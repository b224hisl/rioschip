magic
tech sky130B
magscale 1 2
timestamp 1667228943
<< obsli1 >>
rect 1104 2159 388884 387345
<< obsm1 >>
rect 14 2128 389698 387376
<< metal2 >>
rect 18 389200 74 390000
rect 1306 389200 1362 390000
rect 2594 389200 2650 390000
rect 3882 389200 3938 390000
rect 5170 389200 5226 390000
rect 6458 389200 6514 390000
rect 7746 389200 7802 390000
rect 9034 389200 9090 390000
rect 9678 389200 9734 390000
rect 10966 389200 11022 390000
rect 12254 389200 12310 390000
rect 13542 389200 13598 390000
rect 14830 389200 14886 390000
rect 16118 389200 16174 390000
rect 17406 389200 17462 390000
rect 18694 389200 18750 390000
rect 19982 389200 20038 390000
rect 21270 389200 21326 390000
rect 22558 389200 22614 390000
rect 23846 389200 23902 390000
rect 25134 389200 25190 390000
rect 26422 389200 26478 390000
rect 27710 389200 27766 390000
rect 28998 389200 29054 390000
rect 30286 389200 30342 390000
rect 31574 389200 31630 390000
rect 32862 389200 32918 390000
rect 34150 389200 34206 390000
rect 35438 389200 35494 390000
rect 36726 389200 36782 390000
rect 38014 389200 38070 390000
rect 39302 389200 39358 390000
rect 40590 389200 40646 390000
rect 41878 389200 41934 390000
rect 43166 389200 43222 390000
rect 44454 389200 44510 390000
rect 45742 389200 45798 390000
rect 47030 389200 47086 390000
rect 48318 389200 48374 390000
rect 49606 389200 49662 390000
rect 50894 389200 50950 390000
rect 52182 389200 52238 390000
rect 53470 389200 53526 390000
rect 54758 389200 54814 390000
rect 56046 389200 56102 390000
rect 57334 389200 57390 390000
rect 58622 389200 58678 390000
rect 59910 389200 59966 390000
rect 61198 389200 61254 390000
rect 62486 389200 62542 390000
rect 63774 389200 63830 390000
rect 65062 389200 65118 390000
rect 66350 389200 66406 390000
rect 67638 389200 67694 390000
rect 68926 389200 68982 390000
rect 70214 389200 70270 390000
rect 71502 389200 71558 390000
rect 72790 389200 72846 390000
rect 74078 389200 74134 390000
rect 75366 389200 75422 390000
rect 76654 389200 76710 390000
rect 77942 389200 77998 390000
rect 79230 389200 79286 390000
rect 80518 389200 80574 390000
rect 81806 389200 81862 390000
rect 83094 389200 83150 390000
rect 84382 389200 84438 390000
rect 85670 389200 85726 390000
rect 86958 389200 87014 390000
rect 88246 389200 88302 390000
rect 89534 389200 89590 390000
rect 90822 389200 90878 390000
rect 92110 389200 92166 390000
rect 93398 389200 93454 390000
rect 94686 389200 94742 390000
rect 95974 389200 96030 390000
rect 97262 389200 97318 390000
rect 98550 389200 98606 390000
rect 99838 389200 99894 390000
rect 101126 389200 101182 390000
rect 102414 389200 102470 390000
rect 103702 389200 103758 390000
rect 104990 389200 105046 390000
rect 105634 389200 105690 390000
rect 106922 389200 106978 390000
rect 108210 389200 108266 390000
rect 109498 389200 109554 390000
rect 110786 389200 110842 390000
rect 112074 389200 112130 390000
rect 113362 389200 113418 390000
rect 114650 389200 114706 390000
rect 115938 389200 115994 390000
rect 117226 389200 117282 390000
rect 118514 389200 118570 390000
rect 119802 389200 119858 390000
rect 121090 389200 121146 390000
rect 122378 389200 122434 390000
rect 123666 389200 123722 390000
rect 124954 389200 125010 390000
rect 126242 389200 126298 390000
rect 127530 389200 127586 390000
rect 128818 389200 128874 390000
rect 130106 389200 130162 390000
rect 131394 389200 131450 390000
rect 132682 389200 132738 390000
rect 133970 389200 134026 390000
rect 135258 389200 135314 390000
rect 136546 389200 136602 390000
rect 137834 389200 137890 390000
rect 139122 389200 139178 390000
rect 140410 389200 140466 390000
rect 141698 389200 141754 390000
rect 142986 389200 143042 390000
rect 144274 389200 144330 390000
rect 145562 389200 145618 390000
rect 146850 389200 146906 390000
rect 148138 389200 148194 390000
rect 149426 389200 149482 390000
rect 150714 389200 150770 390000
rect 152002 389200 152058 390000
rect 153290 389200 153346 390000
rect 154578 389200 154634 390000
rect 155866 389200 155922 390000
rect 157154 389200 157210 390000
rect 158442 389200 158498 390000
rect 159730 389200 159786 390000
rect 161018 389200 161074 390000
rect 162306 389200 162362 390000
rect 163594 389200 163650 390000
rect 164882 389200 164938 390000
rect 166170 389200 166226 390000
rect 167458 389200 167514 390000
rect 168746 389200 168802 390000
rect 170034 389200 170090 390000
rect 171322 389200 171378 390000
rect 172610 389200 172666 390000
rect 173898 389200 173954 390000
rect 175186 389200 175242 390000
rect 176474 389200 176530 390000
rect 177762 389200 177818 390000
rect 179050 389200 179106 390000
rect 180338 389200 180394 390000
rect 181626 389200 181682 390000
rect 182914 389200 182970 390000
rect 184202 389200 184258 390000
rect 185490 389200 185546 390000
rect 186778 389200 186834 390000
rect 188066 389200 188122 390000
rect 189354 389200 189410 390000
rect 190642 389200 190698 390000
rect 191930 389200 191986 390000
rect 193218 389200 193274 390000
rect 194506 389200 194562 390000
rect 195794 389200 195850 390000
rect 197082 389200 197138 390000
rect 198370 389200 198426 390000
rect 199658 389200 199714 390000
rect 200302 389200 200358 390000
rect 201590 389200 201646 390000
rect 202878 389200 202934 390000
rect 204166 389200 204222 390000
rect 205454 389200 205510 390000
rect 206742 389200 206798 390000
rect 208030 389200 208086 390000
rect 209318 389200 209374 390000
rect 210606 389200 210662 390000
rect 211894 389200 211950 390000
rect 213182 389200 213238 390000
rect 214470 389200 214526 390000
rect 215758 389200 215814 390000
rect 217046 389200 217102 390000
rect 218334 389200 218390 390000
rect 219622 389200 219678 390000
rect 220910 389200 220966 390000
rect 222198 389200 222254 390000
rect 223486 389200 223542 390000
rect 224774 389200 224830 390000
rect 226062 389200 226118 390000
rect 227350 389200 227406 390000
rect 228638 389200 228694 390000
rect 229926 389200 229982 390000
rect 231214 389200 231270 390000
rect 232502 389200 232558 390000
rect 233790 389200 233846 390000
rect 235078 389200 235134 390000
rect 236366 389200 236422 390000
rect 237654 389200 237710 390000
rect 238942 389200 238998 390000
rect 240230 389200 240286 390000
rect 241518 389200 241574 390000
rect 242806 389200 242862 390000
rect 244094 389200 244150 390000
rect 245382 389200 245438 390000
rect 246670 389200 246726 390000
rect 247958 389200 248014 390000
rect 249246 389200 249302 390000
rect 250534 389200 250590 390000
rect 251822 389200 251878 390000
rect 253110 389200 253166 390000
rect 254398 389200 254454 390000
rect 255686 389200 255742 390000
rect 256974 389200 257030 390000
rect 258262 389200 258318 390000
rect 259550 389200 259606 390000
rect 260838 389200 260894 390000
rect 262126 389200 262182 390000
rect 263414 389200 263470 390000
rect 264702 389200 264758 390000
rect 265990 389200 266046 390000
rect 267278 389200 267334 390000
rect 268566 389200 268622 390000
rect 269854 389200 269910 390000
rect 271142 389200 271198 390000
rect 272430 389200 272486 390000
rect 273718 389200 273774 390000
rect 275006 389200 275062 390000
rect 276294 389200 276350 390000
rect 277582 389200 277638 390000
rect 278870 389200 278926 390000
rect 280158 389200 280214 390000
rect 281446 389200 281502 390000
rect 282734 389200 282790 390000
rect 284022 389200 284078 390000
rect 285310 389200 285366 390000
rect 286598 389200 286654 390000
rect 287886 389200 287942 390000
rect 289174 389200 289230 390000
rect 290462 389200 290518 390000
rect 291750 389200 291806 390000
rect 293038 389200 293094 390000
rect 294326 389200 294382 390000
rect 294970 389200 295026 390000
rect 296258 389200 296314 390000
rect 297546 389200 297602 390000
rect 298834 389200 298890 390000
rect 300122 389200 300178 390000
rect 301410 389200 301466 390000
rect 302698 389200 302754 390000
rect 303986 389200 304042 390000
rect 305274 389200 305330 390000
rect 306562 389200 306618 390000
rect 307850 389200 307906 390000
rect 309138 389200 309194 390000
rect 310426 389200 310482 390000
rect 311714 389200 311770 390000
rect 313002 389200 313058 390000
rect 314290 389200 314346 390000
rect 315578 389200 315634 390000
rect 316866 389200 316922 390000
rect 318154 389200 318210 390000
rect 319442 389200 319498 390000
rect 320730 389200 320786 390000
rect 322018 389200 322074 390000
rect 323306 389200 323362 390000
rect 324594 389200 324650 390000
rect 325882 389200 325938 390000
rect 327170 389200 327226 390000
rect 328458 389200 328514 390000
rect 329746 389200 329802 390000
rect 331034 389200 331090 390000
rect 332322 389200 332378 390000
rect 333610 389200 333666 390000
rect 334898 389200 334954 390000
rect 336186 389200 336242 390000
rect 337474 389200 337530 390000
rect 338762 389200 338818 390000
rect 340050 389200 340106 390000
rect 341338 389200 341394 390000
rect 342626 389200 342682 390000
rect 343914 389200 343970 390000
rect 345202 389200 345258 390000
rect 346490 389200 346546 390000
rect 347778 389200 347834 390000
rect 349066 389200 349122 390000
rect 350354 389200 350410 390000
rect 351642 389200 351698 390000
rect 352930 389200 352986 390000
rect 354218 389200 354274 390000
rect 355506 389200 355562 390000
rect 356794 389200 356850 390000
rect 358082 389200 358138 390000
rect 359370 389200 359426 390000
rect 360658 389200 360714 390000
rect 361946 389200 362002 390000
rect 363234 389200 363290 390000
rect 364522 389200 364578 390000
rect 365810 389200 365866 390000
rect 367098 389200 367154 390000
rect 368386 389200 368442 390000
rect 369674 389200 369730 390000
rect 370962 389200 371018 390000
rect 372250 389200 372306 390000
rect 373538 389200 373594 390000
rect 374826 389200 374882 390000
rect 376114 389200 376170 390000
rect 377402 389200 377458 390000
rect 378690 389200 378746 390000
rect 379978 389200 380034 390000
rect 381266 389200 381322 390000
rect 382554 389200 382610 390000
rect 383842 389200 383898 390000
rect 385130 389200 385186 390000
rect 386418 389200 386474 390000
rect 387706 389200 387762 390000
rect 388994 389200 389050 390000
rect 389638 389200 389694 390000
rect 18 0 74 800
rect 662 0 718 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 30286 0 30342 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36726 0 36782 800
rect 38014 0 38070 800
rect 39302 0 39358 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 43166 0 43222 800
rect 44454 0 44510 800
rect 45742 0 45798 800
rect 47030 0 47086 800
rect 48318 0 48374 800
rect 49606 0 49662 800
rect 50894 0 50950 800
rect 52182 0 52238 800
rect 53470 0 53526 800
rect 54758 0 54814 800
rect 56046 0 56102 800
rect 57334 0 57390 800
rect 58622 0 58678 800
rect 59910 0 59966 800
rect 61198 0 61254 800
rect 62486 0 62542 800
rect 63774 0 63830 800
rect 65062 0 65118 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68926 0 68982 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 77942 0 77998 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 84382 0 84438 800
rect 85670 0 85726 800
rect 86958 0 87014 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 90822 0 90878 800
rect 92110 0 92166 800
rect 93398 0 93454 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 96618 0 96674 800
rect 97906 0 97962 800
rect 99194 0 99250 800
rect 100482 0 100538 800
rect 101770 0 101826 800
rect 103058 0 103114 800
rect 104346 0 104402 800
rect 105634 0 105690 800
rect 106922 0 106978 800
rect 108210 0 108266 800
rect 109498 0 109554 800
rect 110786 0 110842 800
rect 112074 0 112130 800
rect 113362 0 113418 800
rect 114650 0 114706 800
rect 115938 0 115994 800
rect 117226 0 117282 800
rect 118514 0 118570 800
rect 119802 0 119858 800
rect 121090 0 121146 800
rect 122378 0 122434 800
rect 123666 0 123722 800
rect 124954 0 125010 800
rect 126242 0 126298 800
rect 127530 0 127586 800
rect 128818 0 128874 800
rect 130106 0 130162 800
rect 131394 0 131450 800
rect 132682 0 132738 800
rect 133970 0 134026 800
rect 135258 0 135314 800
rect 136546 0 136602 800
rect 137834 0 137890 800
rect 139122 0 139178 800
rect 140410 0 140466 800
rect 141698 0 141754 800
rect 142986 0 143042 800
rect 144274 0 144330 800
rect 145562 0 145618 800
rect 146850 0 146906 800
rect 148138 0 148194 800
rect 149426 0 149482 800
rect 150714 0 150770 800
rect 152002 0 152058 800
rect 153290 0 153346 800
rect 154578 0 154634 800
rect 155866 0 155922 800
rect 157154 0 157210 800
rect 158442 0 158498 800
rect 159730 0 159786 800
rect 161018 0 161074 800
rect 162306 0 162362 800
rect 163594 0 163650 800
rect 164882 0 164938 800
rect 166170 0 166226 800
rect 167458 0 167514 800
rect 168746 0 168802 800
rect 170034 0 170090 800
rect 171322 0 171378 800
rect 172610 0 172666 800
rect 173898 0 173954 800
rect 175186 0 175242 800
rect 176474 0 176530 800
rect 177762 0 177818 800
rect 179050 0 179106 800
rect 180338 0 180394 800
rect 181626 0 181682 800
rect 182914 0 182970 800
rect 184202 0 184258 800
rect 185490 0 185546 800
rect 186778 0 186834 800
rect 188066 0 188122 800
rect 189354 0 189410 800
rect 189998 0 190054 800
rect 191286 0 191342 800
rect 192574 0 192630 800
rect 193862 0 193918 800
rect 195150 0 195206 800
rect 196438 0 196494 800
rect 197726 0 197782 800
rect 199014 0 199070 800
rect 200302 0 200358 800
rect 201590 0 201646 800
rect 202878 0 202934 800
rect 204166 0 204222 800
rect 205454 0 205510 800
rect 206742 0 206798 800
rect 208030 0 208086 800
rect 209318 0 209374 800
rect 210606 0 210662 800
rect 211894 0 211950 800
rect 213182 0 213238 800
rect 214470 0 214526 800
rect 215758 0 215814 800
rect 217046 0 217102 800
rect 218334 0 218390 800
rect 219622 0 219678 800
rect 220910 0 220966 800
rect 222198 0 222254 800
rect 223486 0 223542 800
rect 224774 0 224830 800
rect 226062 0 226118 800
rect 227350 0 227406 800
rect 228638 0 228694 800
rect 229926 0 229982 800
rect 231214 0 231270 800
rect 232502 0 232558 800
rect 233790 0 233846 800
rect 235078 0 235134 800
rect 236366 0 236422 800
rect 237654 0 237710 800
rect 238942 0 238998 800
rect 240230 0 240286 800
rect 241518 0 241574 800
rect 242806 0 242862 800
rect 244094 0 244150 800
rect 245382 0 245438 800
rect 246670 0 246726 800
rect 247958 0 248014 800
rect 249246 0 249302 800
rect 250534 0 250590 800
rect 251822 0 251878 800
rect 253110 0 253166 800
rect 254398 0 254454 800
rect 255686 0 255742 800
rect 256974 0 257030 800
rect 258262 0 258318 800
rect 259550 0 259606 800
rect 260838 0 260894 800
rect 262126 0 262182 800
rect 263414 0 263470 800
rect 264702 0 264758 800
rect 265990 0 266046 800
rect 267278 0 267334 800
rect 268566 0 268622 800
rect 269854 0 269910 800
rect 271142 0 271198 800
rect 272430 0 272486 800
rect 273718 0 273774 800
rect 275006 0 275062 800
rect 276294 0 276350 800
rect 277582 0 277638 800
rect 278870 0 278926 800
rect 280158 0 280214 800
rect 281446 0 281502 800
rect 282734 0 282790 800
rect 284022 0 284078 800
rect 284666 0 284722 800
rect 285954 0 286010 800
rect 287242 0 287298 800
rect 288530 0 288586 800
rect 289818 0 289874 800
rect 291106 0 291162 800
rect 292394 0 292450 800
rect 293682 0 293738 800
rect 294970 0 295026 800
rect 296258 0 296314 800
rect 297546 0 297602 800
rect 298834 0 298890 800
rect 300122 0 300178 800
rect 301410 0 301466 800
rect 302698 0 302754 800
rect 303986 0 304042 800
rect 305274 0 305330 800
rect 306562 0 306618 800
rect 307850 0 307906 800
rect 309138 0 309194 800
rect 310426 0 310482 800
rect 311714 0 311770 800
rect 313002 0 313058 800
rect 314290 0 314346 800
rect 315578 0 315634 800
rect 316866 0 316922 800
rect 318154 0 318210 800
rect 319442 0 319498 800
rect 320730 0 320786 800
rect 322018 0 322074 800
rect 323306 0 323362 800
rect 324594 0 324650 800
rect 325882 0 325938 800
rect 327170 0 327226 800
rect 328458 0 328514 800
rect 329746 0 329802 800
rect 331034 0 331090 800
rect 332322 0 332378 800
rect 333610 0 333666 800
rect 334898 0 334954 800
rect 336186 0 336242 800
rect 337474 0 337530 800
rect 338762 0 338818 800
rect 340050 0 340106 800
rect 341338 0 341394 800
rect 342626 0 342682 800
rect 343914 0 343970 800
rect 345202 0 345258 800
rect 346490 0 346546 800
rect 347778 0 347834 800
rect 349066 0 349122 800
rect 350354 0 350410 800
rect 351642 0 351698 800
rect 352930 0 352986 800
rect 354218 0 354274 800
rect 355506 0 355562 800
rect 356794 0 356850 800
rect 358082 0 358138 800
rect 359370 0 359426 800
rect 360658 0 360714 800
rect 361946 0 362002 800
rect 363234 0 363290 800
rect 364522 0 364578 800
rect 365810 0 365866 800
rect 367098 0 367154 800
rect 368386 0 368442 800
rect 369674 0 369730 800
rect 370962 0 371018 800
rect 372250 0 372306 800
rect 373538 0 373594 800
rect 374826 0 374882 800
rect 376114 0 376170 800
rect 377402 0 377458 800
rect 378690 0 378746 800
rect 379978 0 380034 800
rect 380622 0 380678 800
rect 381910 0 381966 800
rect 383198 0 383254 800
rect 384486 0 384542 800
rect 385774 0 385830 800
rect 387062 0 387118 800
rect 388350 0 388406 800
rect 389638 0 389694 800
<< obsm2 >>
rect 130 389144 1250 389314
rect 1418 389144 2538 389314
rect 2706 389144 3826 389314
rect 3994 389144 5114 389314
rect 5282 389144 6402 389314
rect 6570 389144 7690 389314
rect 7858 389144 8978 389314
rect 9146 389144 9622 389314
rect 9790 389144 10910 389314
rect 11078 389144 12198 389314
rect 12366 389144 13486 389314
rect 13654 389144 14774 389314
rect 14942 389144 16062 389314
rect 16230 389144 17350 389314
rect 17518 389144 18638 389314
rect 18806 389144 19926 389314
rect 20094 389144 21214 389314
rect 21382 389144 22502 389314
rect 22670 389144 23790 389314
rect 23958 389144 25078 389314
rect 25246 389144 26366 389314
rect 26534 389144 27654 389314
rect 27822 389144 28942 389314
rect 29110 389144 30230 389314
rect 30398 389144 31518 389314
rect 31686 389144 32806 389314
rect 32974 389144 34094 389314
rect 34262 389144 35382 389314
rect 35550 389144 36670 389314
rect 36838 389144 37958 389314
rect 38126 389144 39246 389314
rect 39414 389144 40534 389314
rect 40702 389144 41822 389314
rect 41990 389144 43110 389314
rect 43278 389144 44398 389314
rect 44566 389144 45686 389314
rect 45854 389144 46974 389314
rect 47142 389144 48262 389314
rect 48430 389144 49550 389314
rect 49718 389144 50838 389314
rect 51006 389144 52126 389314
rect 52294 389144 53414 389314
rect 53582 389144 54702 389314
rect 54870 389144 55990 389314
rect 56158 389144 57278 389314
rect 57446 389144 58566 389314
rect 58734 389144 59854 389314
rect 60022 389144 61142 389314
rect 61310 389144 62430 389314
rect 62598 389144 63718 389314
rect 63886 389144 65006 389314
rect 65174 389144 66294 389314
rect 66462 389144 67582 389314
rect 67750 389144 68870 389314
rect 69038 389144 70158 389314
rect 70326 389144 71446 389314
rect 71614 389144 72734 389314
rect 72902 389144 74022 389314
rect 74190 389144 75310 389314
rect 75478 389144 76598 389314
rect 76766 389144 77886 389314
rect 78054 389144 79174 389314
rect 79342 389144 80462 389314
rect 80630 389144 81750 389314
rect 81918 389144 83038 389314
rect 83206 389144 84326 389314
rect 84494 389144 85614 389314
rect 85782 389144 86902 389314
rect 87070 389144 88190 389314
rect 88358 389144 89478 389314
rect 89646 389144 90766 389314
rect 90934 389144 92054 389314
rect 92222 389144 93342 389314
rect 93510 389144 94630 389314
rect 94798 389144 95918 389314
rect 96086 389144 97206 389314
rect 97374 389144 98494 389314
rect 98662 389144 99782 389314
rect 99950 389144 101070 389314
rect 101238 389144 102358 389314
rect 102526 389144 103646 389314
rect 103814 389144 104934 389314
rect 105102 389144 105578 389314
rect 105746 389144 106866 389314
rect 107034 389144 108154 389314
rect 108322 389144 109442 389314
rect 109610 389144 110730 389314
rect 110898 389144 112018 389314
rect 112186 389144 113306 389314
rect 113474 389144 114594 389314
rect 114762 389144 115882 389314
rect 116050 389144 117170 389314
rect 117338 389144 118458 389314
rect 118626 389144 119746 389314
rect 119914 389144 121034 389314
rect 121202 389144 122322 389314
rect 122490 389144 123610 389314
rect 123778 389144 124898 389314
rect 125066 389144 126186 389314
rect 126354 389144 127474 389314
rect 127642 389144 128762 389314
rect 128930 389144 130050 389314
rect 130218 389144 131338 389314
rect 131506 389144 132626 389314
rect 132794 389144 133914 389314
rect 134082 389144 135202 389314
rect 135370 389144 136490 389314
rect 136658 389144 137778 389314
rect 137946 389144 139066 389314
rect 139234 389144 140354 389314
rect 140522 389144 141642 389314
rect 141810 389144 142930 389314
rect 143098 389144 144218 389314
rect 144386 389144 145506 389314
rect 145674 389144 146794 389314
rect 146962 389144 148082 389314
rect 148250 389144 149370 389314
rect 149538 389144 150658 389314
rect 150826 389144 151946 389314
rect 152114 389144 153234 389314
rect 153402 389144 154522 389314
rect 154690 389144 155810 389314
rect 155978 389144 157098 389314
rect 157266 389144 158386 389314
rect 158554 389144 159674 389314
rect 159842 389144 160962 389314
rect 161130 389144 162250 389314
rect 162418 389144 163538 389314
rect 163706 389144 164826 389314
rect 164994 389144 166114 389314
rect 166282 389144 167402 389314
rect 167570 389144 168690 389314
rect 168858 389144 169978 389314
rect 170146 389144 171266 389314
rect 171434 389144 172554 389314
rect 172722 389144 173842 389314
rect 174010 389144 175130 389314
rect 175298 389144 176418 389314
rect 176586 389144 177706 389314
rect 177874 389144 178994 389314
rect 179162 389144 180282 389314
rect 180450 389144 181570 389314
rect 181738 389144 182858 389314
rect 183026 389144 184146 389314
rect 184314 389144 185434 389314
rect 185602 389144 186722 389314
rect 186890 389144 188010 389314
rect 188178 389144 189298 389314
rect 189466 389144 190586 389314
rect 190754 389144 191874 389314
rect 192042 389144 193162 389314
rect 193330 389144 194450 389314
rect 194618 389144 195738 389314
rect 195906 389144 197026 389314
rect 197194 389144 198314 389314
rect 198482 389144 199602 389314
rect 199770 389144 200246 389314
rect 200414 389144 201534 389314
rect 201702 389144 202822 389314
rect 202990 389144 204110 389314
rect 204278 389144 205398 389314
rect 205566 389144 206686 389314
rect 206854 389144 207974 389314
rect 208142 389144 209262 389314
rect 209430 389144 210550 389314
rect 210718 389144 211838 389314
rect 212006 389144 213126 389314
rect 213294 389144 214414 389314
rect 214582 389144 215702 389314
rect 215870 389144 216990 389314
rect 217158 389144 218278 389314
rect 218446 389144 219566 389314
rect 219734 389144 220854 389314
rect 221022 389144 222142 389314
rect 222310 389144 223430 389314
rect 223598 389144 224718 389314
rect 224886 389144 226006 389314
rect 226174 389144 227294 389314
rect 227462 389144 228582 389314
rect 228750 389144 229870 389314
rect 230038 389144 231158 389314
rect 231326 389144 232446 389314
rect 232614 389144 233734 389314
rect 233902 389144 235022 389314
rect 235190 389144 236310 389314
rect 236478 389144 237598 389314
rect 237766 389144 238886 389314
rect 239054 389144 240174 389314
rect 240342 389144 241462 389314
rect 241630 389144 242750 389314
rect 242918 389144 244038 389314
rect 244206 389144 245326 389314
rect 245494 389144 246614 389314
rect 246782 389144 247902 389314
rect 248070 389144 249190 389314
rect 249358 389144 250478 389314
rect 250646 389144 251766 389314
rect 251934 389144 253054 389314
rect 253222 389144 254342 389314
rect 254510 389144 255630 389314
rect 255798 389144 256918 389314
rect 257086 389144 258206 389314
rect 258374 389144 259494 389314
rect 259662 389144 260782 389314
rect 260950 389144 262070 389314
rect 262238 389144 263358 389314
rect 263526 389144 264646 389314
rect 264814 389144 265934 389314
rect 266102 389144 267222 389314
rect 267390 389144 268510 389314
rect 268678 389144 269798 389314
rect 269966 389144 271086 389314
rect 271254 389144 272374 389314
rect 272542 389144 273662 389314
rect 273830 389144 274950 389314
rect 275118 389144 276238 389314
rect 276406 389144 277526 389314
rect 277694 389144 278814 389314
rect 278982 389144 280102 389314
rect 280270 389144 281390 389314
rect 281558 389144 282678 389314
rect 282846 389144 283966 389314
rect 284134 389144 285254 389314
rect 285422 389144 286542 389314
rect 286710 389144 287830 389314
rect 287998 389144 289118 389314
rect 289286 389144 290406 389314
rect 290574 389144 291694 389314
rect 291862 389144 292982 389314
rect 293150 389144 294270 389314
rect 294438 389144 294914 389314
rect 295082 389144 296202 389314
rect 296370 389144 297490 389314
rect 297658 389144 298778 389314
rect 298946 389144 300066 389314
rect 300234 389144 301354 389314
rect 301522 389144 302642 389314
rect 302810 389144 303930 389314
rect 304098 389144 305218 389314
rect 305386 389144 306506 389314
rect 306674 389144 307794 389314
rect 307962 389144 309082 389314
rect 309250 389144 310370 389314
rect 310538 389144 311658 389314
rect 311826 389144 312946 389314
rect 313114 389144 314234 389314
rect 314402 389144 315522 389314
rect 315690 389144 316810 389314
rect 316978 389144 318098 389314
rect 318266 389144 319386 389314
rect 319554 389144 320674 389314
rect 320842 389144 321962 389314
rect 322130 389144 323250 389314
rect 323418 389144 324538 389314
rect 324706 389144 325826 389314
rect 325994 389144 327114 389314
rect 327282 389144 328402 389314
rect 328570 389144 329690 389314
rect 329858 389144 330978 389314
rect 331146 389144 332266 389314
rect 332434 389144 333554 389314
rect 333722 389144 334842 389314
rect 335010 389144 336130 389314
rect 336298 389144 337418 389314
rect 337586 389144 338706 389314
rect 338874 389144 339994 389314
rect 340162 389144 341282 389314
rect 341450 389144 342570 389314
rect 342738 389144 343858 389314
rect 344026 389144 345146 389314
rect 345314 389144 346434 389314
rect 346602 389144 347722 389314
rect 347890 389144 349010 389314
rect 349178 389144 350298 389314
rect 350466 389144 351586 389314
rect 351754 389144 352874 389314
rect 353042 389144 354162 389314
rect 354330 389144 355450 389314
rect 355618 389144 356738 389314
rect 356906 389144 358026 389314
rect 358194 389144 359314 389314
rect 359482 389144 360602 389314
rect 360770 389144 361890 389314
rect 362058 389144 363178 389314
rect 363346 389144 364466 389314
rect 364634 389144 365754 389314
rect 365922 389144 367042 389314
rect 367210 389144 368330 389314
rect 368498 389144 369618 389314
rect 369786 389144 370906 389314
rect 371074 389144 372194 389314
rect 372362 389144 373482 389314
rect 373650 389144 374770 389314
rect 374938 389144 376058 389314
rect 376226 389144 377346 389314
rect 377514 389144 378634 389314
rect 378802 389144 379922 389314
rect 380090 389144 381210 389314
rect 381378 389144 382498 389314
rect 382666 389144 383786 389314
rect 383954 389144 385074 389314
rect 385242 389144 386362 389314
rect 386530 389144 387650 389314
rect 387818 389144 388938 389314
rect 389106 389144 389582 389314
rect 20 856 389692 389144
rect 130 734 606 856
rect 774 734 1894 856
rect 2062 734 3182 856
rect 3350 734 4470 856
rect 4638 734 5758 856
rect 5926 734 7046 856
rect 7214 734 8334 856
rect 8502 734 9622 856
rect 9790 734 10910 856
rect 11078 734 12198 856
rect 12366 734 13486 856
rect 13654 734 14774 856
rect 14942 734 16062 856
rect 16230 734 17350 856
rect 17518 734 18638 856
rect 18806 734 19926 856
rect 20094 734 21214 856
rect 21382 734 22502 856
rect 22670 734 23790 856
rect 23958 734 25078 856
rect 25246 734 26366 856
rect 26534 734 27654 856
rect 27822 734 28942 856
rect 29110 734 30230 856
rect 30398 734 31518 856
rect 31686 734 32806 856
rect 32974 734 34094 856
rect 34262 734 35382 856
rect 35550 734 36670 856
rect 36838 734 37958 856
rect 38126 734 39246 856
rect 39414 734 40534 856
rect 40702 734 41822 856
rect 41990 734 43110 856
rect 43278 734 44398 856
rect 44566 734 45686 856
rect 45854 734 46974 856
rect 47142 734 48262 856
rect 48430 734 49550 856
rect 49718 734 50838 856
rect 51006 734 52126 856
rect 52294 734 53414 856
rect 53582 734 54702 856
rect 54870 734 55990 856
rect 56158 734 57278 856
rect 57446 734 58566 856
rect 58734 734 59854 856
rect 60022 734 61142 856
rect 61310 734 62430 856
rect 62598 734 63718 856
rect 63886 734 65006 856
rect 65174 734 66294 856
rect 66462 734 67582 856
rect 67750 734 68870 856
rect 69038 734 70158 856
rect 70326 734 71446 856
rect 71614 734 72734 856
rect 72902 734 74022 856
rect 74190 734 75310 856
rect 75478 734 76598 856
rect 76766 734 77886 856
rect 78054 734 79174 856
rect 79342 734 80462 856
rect 80630 734 81750 856
rect 81918 734 83038 856
rect 83206 734 84326 856
rect 84494 734 85614 856
rect 85782 734 86902 856
rect 87070 734 88190 856
rect 88358 734 89478 856
rect 89646 734 90766 856
rect 90934 734 92054 856
rect 92222 734 93342 856
rect 93510 734 94630 856
rect 94798 734 95274 856
rect 95442 734 96562 856
rect 96730 734 97850 856
rect 98018 734 99138 856
rect 99306 734 100426 856
rect 100594 734 101714 856
rect 101882 734 103002 856
rect 103170 734 104290 856
rect 104458 734 105578 856
rect 105746 734 106866 856
rect 107034 734 108154 856
rect 108322 734 109442 856
rect 109610 734 110730 856
rect 110898 734 112018 856
rect 112186 734 113306 856
rect 113474 734 114594 856
rect 114762 734 115882 856
rect 116050 734 117170 856
rect 117338 734 118458 856
rect 118626 734 119746 856
rect 119914 734 121034 856
rect 121202 734 122322 856
rect 122490 734 123610 856
rect 123778 734 124898 856
rect 125066 734 126186 856
rect 126354 734 127474 856
rect 127642 734 128762 856
rect 128930 734 130050 856
rect 130218 734 131338 856
rect 131506 734 132626 856
rect 132794 734 133914 856
rect 134082 734 135202 856
rect 135370 734 136490 856
rect 136658 734 137778 856
rect 137946 734 139066 856
rect 139234 734 140354 856
rect 140522 734 141642 856
rect 141810 734 142930 856
rect 143098 734 144218 856
rect 144386 734 145506 856
rect 145674 734 146794 856
rect 146962 734 148082 856
rect 148250 734 149370 856
rect 149538 734 150658 856
rect 150826 734 151946 856
rect 152114 734 153234 856
rect 153402 734 154522 856
rect 154690 734 155810 856
rect 155978 734 157098 856
rect 157266 734 158386 856
rect 158554 734 159674 856
rect 159842 734 160962 856
rect 161130 734 162250 856
rect 162418 734 163538 856
rect 163706 734 164826 856
rect 164994 734 166114 856
rect 166282 734 167402 856
rect 167570 734 168690 856
rect 168858 734 169978 856
rect 170146 734 171266 856
rect 171434 734 172554 856
rect 172722 734 173842 856
rect 174010 734 175130 856
rect 175298 734 176418 856
rect 176586 734 177706 856
rect 177874 734 178994 856
rect 179162 734 180282 856
rect 180450 734 181570 856
rect 181738 734 182858 856
rect 183026 734 184146 856
rect 184314 734 185434 856
rect 185602 734 186722 856
rect 186890 734 188010 856
rect 188178 734 189298 856
rect 189466 734 189942 856
rect 190110 734 191230 856
rect 191398 734 192518 856
rect 192686 734 193806 856
rect 193974 734 195094 856
rect 195262 734 196382 856
rect 196550 734 197670 856
rect 197838 734 198958 856
rect 199126 734 200246 856
rect 200414 734 201534 856
rect 201702 734 202822 856
rect 202990 734 204110 856
rect 204278 734 205398 856
rect 205566 734 206686 856
rect 206854 734 207974 856
rect 208142 734 209262 856
rect 209430 734 210550 856
rect 210718 734 211838 856
rect 212006 734 213126 856
rect 213294 734 214414 856
rect 214582 734 215702 856
rect 215870 734 216990 856
rect 217158 734 218278 856
rect 218446 734 219566 856
rect 219734 734 220854 856
rect 221022 734 222142 856
rect 222310 734 223430 856
rect 223598 734 224718 856
rect 224886 734 226006 856
rect 226174 734 227294 856
rect 227462 734 228582 856
rect 228750 734 229870 856
rect 230038 734 231158 856
rect 231326 734 232446 856
rect 232614 734 233734 856
rect 233902 734 235022 856
rect 235190 734 236310 856
rect 236478 734 237598 856
rect 237766 734 238886 856
rect 239054 734 240174 856
rect 240342 734 241462 856
rect 241630 734 242750 856
rect 242918 734 244038 856
rect 244206 734 245326 856
rect 245494 734 246614 856
rect 246782 734 247902 856
rect 248070 734 249190 856
rect 249358 734 250478 856
rect 250646 734 251766 856
rect 251934 734 253054 856
rect 253222 734 254342 856
rect 254510 734 255630 856
rect 255798 734 256918 856
rect 257086 734 258206 856
rect 258374 734 259494 856
rect 259662 734 260782 856
rect 260950 734 262070 856
rect 262238 734 263358 856
rect 263526 734 264646 856
rect 264814 734 265934 856
rect 266102 734 267222 856
rect 267390 734 268510 856
rect 268678 734 269798 856
rect 269966 734 271086 856
rect 271254 734 272374 856
rect 272542 734 273662 856
rect 273830 734 274950 856
rect 275118 734 276238 856
rect 276406 734 277526 856
rect 277694 734 278814 856
rect 278982 734 280102 856
rect 280270 734 281390 856
rect 281558 734 282678 856
rect 282846 734 283966 856
rect 284134 734 284610 856
rect 284778 734 285898 856
rect 286066 734 287186 856
rect 287354 734 288474 856
rect 288642 734 289762 856
rect 289930 734 291050 856
rect 291218 734 292338 856
rect 292506 734 293626 856
rect 293794 734 294914 856
rect 295082 734 296202 856
rect 296370 734 297490 856
rect 297658 734 298778 856
rect 298946 734 300066 856
rect 300234 734 301354 856
rect 301522 734 302642 856
rect 302810 734 303930 856
rect 304098 734 305218 856
rect 305386 734 306506 856
rect 306674 734 307794 856
rect 307962 734 309082 856
rect 309250 734 310370 856
rect 310538 734 311658 856
rect 311826 734 312946 856
rect 313114 734 314234 856
rect 314402 734 315522 856
rect 315690 734 316810 856
rect 316978 734 318098 856
rect 318266 734 319386 856
rect 319554 734 320674 856
rect 320842 734 321962 856
rect 322130 734 323250 856
rect 323418 734 324538 856
rect 324706 734 325826 856
rect 325994 734 327114 856
rect 327282 734 328402 856
rect 328570 734 329690 856
rect 329858 734 330978 856
rect 331146 734 332266 856
rect 332434 734 333554 856
rect 333722 734 334842 856
rect 335010 734 336130 856
rect 336298 734 337418 856
rect 337586 734 338706 856
rect 338874 734 339994 856
rect 340162 734 341282 856
rect 341450 734 342570 856
rect 342738 734 343858 856
rect 344026 734 345146 856
rect 345314 734 346434 856
rect 346602 734 347722 856
rect 347890 734 349010 856
rect 349178 734 350298 856
rect 350466 734 351586 856
rect 351754 734 352874 856
rect 353042 734 354162 856
rect 354330 734 355450 856
rect 355618 734 356738 856
rect 356906 734 358026 856
rect 358194 734 359314 856
rect 359482 734 360602 856
rect 360770 734 361890 856
rect 362058 734 363178 856
rect 363346 734 364466 856
rect 364634 734 365754 856
rect 365922 734 367042 856
rect 367210 734 368330 856
rect 368498 734 369618 856
rect 369786 734 370906 856
rect 371074 734 372194 856
rect 372362 734 373482 856
rect 373650 734 374770 856
rect 374938 734 376058 856
rect 376226 734 377346 856
rect 377514 734 378634 856
rect 378802 734 379922 856
rect 380090 734 380566 856
rect 380734 734 381854 856
rect 382022 734 383142 856
rect 383310 734 384430 856
rect 384598 734 385718 856
rect 385886 734 387006 856
rect 387174 734 388294 856
rect 388462 734 389582 856
<< metal3 >>
rect 0 388968 800 389088
rect 389200 388968 390000 389088
rect 0 387608 800 387728
rect 389200 387608 390000 387728
rect 0 386248 800 386368
rect 389200 386248 390000 386368
rect 0 384888 800 385008
rect 389200 384888 390000 385008
rect 0 383528 800 383648
rect 389200 383528 390000 383648
rect 0 382168 800 382288
rect 389200 382168 390000 382288
rect 0 380808 800 380928
rect 389200 380808 390000 380928
rect 0 379448 800 379568
rect 389200 379448 390000 379568
rect 0 378088 800 378208
rect 389200 378088 390000 378208
rect 0 376728 800 376848
rect 389200 376728 390000 376848
rect 0 375368 800 375488
rect 389200 375368 390000 375488
rect 0 374008 800 374128
rect 389200 374008 390000 374128
rect 0 372648 800 372768
rect 389200 372648 390000 372768
rect 0 371288 800 371408
rect 389200 371288 390000 371408
rect 0 369928 800 370048
rect 389200 369928 390000 370048
rect 0 368568 800 368688
rect 389200 368568 390000 368688
rect 0 367208 800 367328
rect 389200 367208 390000 367328
rect 0 365848 800 365968
rect 389200 365848 390000 365968
rect 0 364488 800 364608
rect 389200 364488 390000 364608
rect 0 363128 800 363248
rect 389200 363128 390000 363248
rect 0 361768 800 361888
rect 389200 361768 390000 361888
rect 0 360408 800 360528
rect 389200 360408 390000 360528
rect 0 359048 800 359168
rect 389200 359048 390000 359168
rect 0 357688 800 357808
rect 389200 357688 390000 357808
rect 0 356328 800 356448
rect 389200 356328 390000 356448
rect 0 354968 800 355088
rect 389200 354968 390000 355088
rect 0 353608 800 353728
rect 389200 353608 390000 353728
rect 0 352248 800 352368
rect 389200 352248 390000 352368
rect 0 350888 800 351008
rect 389200 350888 390000 351008
rect 0 349528 800 349648
rect 389200 349528 390000 349648
rect 0 348168 800 348288
rect 389200 348168 390000 348288
rect 0 346808 800 346928
rect 389200 346808 390000 346928
rect 0 345448 800 345568
rect 389200 345448 390000 345568
rect 0 344088 800 344208
rect 389200 344088 390000 344208
rect 0 342728 800 342848
rect 389200 342728 390000 342848
rect 0 341368 800 341488
rect 389200 341368 390000 341488
rect 0 340008 800 340128
rect 389200 340008 390000 340128
rect 0 338648 800 338768
rect 389200 338648 390000 338768
rect 0 337288 800 337408
rect 389200 337288 390000 337408
rect 0 335928 800 336048
rect 389200 335928 390000 336048
rect 0 334568 800 334688
rect 389200 334568 390000 334688
rect 0 333208 800 333328
rect 389200 333208 390000 333328
rect 0 331848 800 331968
rect 389200 331848 390000 331968
rect 0 330488 800 330608
rect 389200 330488 390000 330608
rect 0 329128 800 329248
rect 389200 329128 390000 329248
rect 0 327768 800 327888
rect 389200 327768 390000 327888
rect 0 326408 800 326528
rect 389200 326408 390000 326528
rect 0 325048 800 325168
rect 389200 325048 390000 325168
rect 0 323688 800 323808
rect 389200 323688 390000 323808
rect 0 322328 800 322448
rect 389200 322328 390000 322448
rect 0 320968 800 321088
rect 389200 320968 390000 321088
rect 0 319608 800 319728
rect 389200 319608 390000 319728
rect 0 318248 800 318368
rect 389200 318248 390000 318368
rect 0 316888 800 317008
rect 389200 316888 390000 317008
rect 0 315528 800 315648
rect 389200 315528 390000 315648
rect 0 314168 800 314288
rect 389200 314168 390000 314288
rect 0 312808 800 312928
rect 389200 312808 390000 312928
rect 0 311448 800 311568
rect 389200 311448 390000 311568
rect 0 310088 800 310208
rect 389200 310088 390000 310208
rect 0 308728 800 308848
rect 389200 308728 390000 308848
rect 0 307368 800 307488
rect 389200 307368 390000 307488
rect 0 306008 800 306128
rect 389200 306008 390000 306128
rect 0 304648 800 304768
rect 389200 304648 390000 304768
rect 0 303288 800 303408
rect 389200 303288 390000 303408
rect 0 301928 800 302048
rect 389200 301928 390000 302048
rect 0 300568 800 300688
rect 389200 300568 390000 300688
rect 0 299888 800 300008
rect 389200 299208 390000 299328
rect 0 298528 800 298648
rect 389200 297848 390000 297968
rect 0 297168 800 297288
rect 389200 296488 390000 296608
rect 0 295808 800 295928
rect 389200 295128 390000 295248
rect 0 294448 800 294568
rect 389200 293768 390000 293888
rect 0 293088 800 293208
rect 389200 292408 390000 292528
rect 0 291728 800 291848
rect 389200 291048 390000 291168
rect 0 290368 800 290488
rect 389200 289688 390000 289808
rect 0 289008 800 289128
rect 389200 289008 390000 289128
rect 0 287648 800 287768
rect 389200 287648 390000 287768
rect 0 286288 800 286408
rect 389200 286288 390000 286408
rect 0 284928 800 285048
rect 389200 284928 390000 285048
rect 0 283568 800 283688
rect 389200 283568 390000 283688
rect 0 282208 800 282328
rect 389200 282208 390000 282328
rect 0 280848 800 280968
rect 389200 280848 390000 280968
rect 0 279488 800 279608
rect 389200 279488 390000 279608
rect 0 278128 800 278248
rect 389200 278128 390000 278248
rect 0 276768 800 276888
rect 389200 276768 390000 276888
rect 0 275408 800 275528
rect 389200 275408 390000 275528
rect 0 274048 800 274168
rect 389200 274048 390000 274168
rect 0 272688 800 272808
rect 389200 272688 390000 272808
rect 0 271328 800 271448
rect 389200 271328 390000 271448
rect 0 269968 800 270088
rect 389200 269968 390000 270088
rect 0 268608 800 268728
rect 389200 268608 390000 268728
rect 0 267248 800 267368
rect 389200 267248 390000 267368
rect 0 265888 800 266008
rect 389200 265888 390000 266008
rect 0 264528 800 264648
rect 389200 264528 390000 264648
rect 0 263168 800 263288
rect 389200 263168 390000 263288
rect 0 261808 800 261928
rect 389200 261808 390000 261928
rect 0 260448 800 260568
rect 389200 260448 390000 260568
rect 0 259088 800 259208
rect 389200 259088 390000 259208
rect 0 257728 800 257848
rect 389200 257728 390000 257848
rect 0 256368 800 256488
rect 389200 256368 390000 256488
rect 0 255008 800 255128
rect 389200 255008 390000 255128
rect 0 253648 800 253768
rect 389200 253648 390000 253768
rect 0 252288 800 252408
rect 389200 252288 390000 252408
rect 0 250928 800 251048
rect 389200 250928 390000 251048
rect 0 249568 800 249688
rect 389200 249568 390000 249688
rect 0 248208 800 248328
rect 389200 248208 390000 248328
rect 0 246848 800 246968
rect 389200 246848 390000 246968
rect 0 245488 800 245608
rect 389200 245488 390000 245608
rect 0 244128 800 244248
rect 389200 244128 390000 244248
rect 0 242768 800 242888
rect 389200 242768 390000 242888
rect 0 241408 800 241528
rect 389200 241408 390000 241528
rect 0 240048 800 240168
rect 389200 240048 390000 240168
rect 0 238688 800 238808
rect 389200 238688 390000 238808
rect 0 237328 800 237448
rect 389200 237328 390000 237448
rect 0 235968 800 236088
rect 389200 235968 390000 236088
rect 0 234608 800 234728
rect 389200 234608 390000 234728
rect 0 233248 800 233368
rect 389200 233248 390000 233368
rect 0 231888 800 232008
rect 389200 231888 390000 232008
rect 0 230528 800 230648
rect 389200 230528 390000 230648
rect 0 229168 800 229288
rect 389200 229168 390000 229288
rect 0 227808 800 227928
rect 389200 227808 390000 227928
rect 0 226448 800 226568
rect 389200 226448 390000 226568
rect 0 225088 800 225208
rect 389200 225088 390000 225208
rect 0 223728 800 223848
rect 389200 223728 390000 223848
rect 0 222368 800 222488
rect 389200 222368 390000 222488
rect 0 221008 800 221128
rect 389200 221008 390000 221128
rect 0 219648 800 219768
rect 389200 219648 390000 219768
rect 0 218288 800 218408
rect 389200 218288 390000 218408
rect 0 216928 800 217048
rect 389200 216928 390000 217048
rect 0 215568 800 215688
rect 389200 215568 390000 215688
rect 0 214208 800 214328
rect 389200 214208 390000 214328
rect 0 212848 800 212968
rect 389200 212848 390000 212968
rect 0 211488 800 211608
rect 389200 211488 390000 211608
rect 0 210128 800 210248
rect 389200 210128 390000 210248
rect 0 208768 800 208888
rect 389200 208768 390000 208888
rect 0 207408 800 207528
rect 389200 207408 390000 207528
rect 0 206048 800 206168
rect 389200 206048 390000 206168
rect 0 204688 800 204808
rect 389200 204688 390000 204808
rect 0 203328 800 203448
rect 389200 203328 390000 203448
rect 0 201968 800 202088
rect 389200 201968 390000 202088
rect 0 200608 800 200728
rect 389200 200608 390000 200728
rect 0 199928 800 200048
rect 389200 199248 390000 199368
rect 0 198568 800 198688
rect 389200 197888 390000 198008
rect 0 197208 800 197328
rect 389200 196528 390000 196648
rect 0 195848 800 195968
rect 389200 195168 390000 195288
rect 0 194488 800 194608
rect 389200 193808 390000 193928
rect 0 193128 800 193248
rect 389200 192448 390000 192568
rect 0 191768 800 191888
rect 389200 191088 390000 191208
rect 0 190408 800 190528
rect 389200 189728 390000 189848
rect 0 189048 800 189168
rect 389200 189048 390000 189168
rect 0 187688 800 187808
rect 389200 187688 390000 187808
rect 0 186328 800 186448
rect 389200 186328 390000 186448
rect 0 184968 800 185088
rect 389200 184968 390000 185088
rect 0 183608 800 183728
rect 389200 183608 390000 183728
rect 0 182248 800 182368
rect 389200 182248 390000 182368
rect 0 180888 800 181008
rect 389200 180888 390000 181008
rect 0 179528 800 179648
rect 389200 179528 390000 179648
rect 0 178168 800 178288
rect 389200 178168 390000 178288
rect 0 176808 800 176928
rect 389200 176808 390000 176928
rect 0 175448 800 175568
rect 389200 175448 390000 175568
rect 0 174088 800 174208
rect 389200 174088 390000 174208
rect 0 172728 800 172848
rect 389200 172728 390000 172848
rect 0 171368 800 171488
rect 389200 171368 390000 171488
rect 0 170008 800 170128
rect 389200 170008 390000 170128
rect 0 168648 800 168768
rect 389200 168648 390000 168768
rect 0 167288 800 167408
rect 389200 167288 390000 167408
rect 0 165928 800 166048
rect 389200 165928 390000 166048
rect 0 164568 800 164688
rect 389200 164568 390000 164688
rect 0 163208 800 163328
rect 389200 163208 390000 163328
rect 0 161848 800 161968
rect 389200 161848 390000 161968
rect 0 160488 800 160608
rect 389200 160488 390000 160608
rect 0 159128 800 159248
rect 389200 159128 390000 159248
rect 0 157768 800 157888
rect 389200 157768 390000 157888
rect 0 156408 800 156528
rect 389200 156408 390000 156528
rect 0 155048 800 155168
rect 389200 155048 390000 155168
rect 0 153688 800 153808
rect 389200 153688 390000 153808
rect 0 152328 800 152448
rect 389200 152328 390000 152448
rect 0 150968 800 151088
rect 389200 150968 390000 151088
rect 0 149608 800 149728
rect 389200 149608 390000 149728
rect 0 148248 800 148368
rect 389200 148248 390000 148368
rect 0 146888 800 147008
rect 389200 146888 390000 147008
rect 0 145528 800 145648
rect 389200 145528 390000 145648
rect 0 144168 800 144288
rect 389200 144168 390000 144288
rect 0 142808 800 142928
rect 389200 142808 390000 142928
rect 0 141448 800 141568
rect 389200 141448 390000 141568
rect 0 140088 800 140208
rect 389200 140088 390000 140208
rect 0 138728 800 138848
rect 389200 138728 390000 138848
rect 0 137368 800 137488
rect 389200 137368 390000 137488
rect 0 136008 800 136128
rect 389200 136008 390000 136128
rect 0 134648 800 134768
rect 389200 134648 390000 134768
rect 0 133288 800 133408
rect 389200 133288 390000 133408
rect 0 131928 800 132048
rect 389200 131928 390000 132048
rect 0 130568 800 130688
rect 389200 130568 390000 130688
rect 0 129208 800 129328
rect 389200 129208 390000 129328
rect 0 127848 800 127968
rect 389200 127848 390000 127968
rect 0 126488 800 126608
rect 389200 126488 390000 126608
rect 0 125128 800 125248
rect 389200 125128 390000 125248
rect 0 123768 800 123888
rect 389200 123768 390000 123888
rect 0 122408 800 122528
rect 389200 122408 390000 122528
rect 0 121048 800 121168
rect 389200 121048 390000 121168
rect 0 119688 800 119808
rect 389200 119688 390000 119808
rect 0 118328 800 118448
rect 389200 118328 390000 118448
rect 0 116968 800 117088
rect 389200 116968 390000 117088
rect 0 115608 800 115728
rect 389200 115608 390000 115728
rect 0 114248 800 114368
rect 389200 114248 390000 114368
rect 0 112888 800 113008
rect 389200 112888 390000 113008
rect 0 111528 800 111648
rect 389200 111528 390000 111648
rect 0 110168 800 110288
rect 389200 110168 390000 110288
rect 0 108808 800 108928
rect 389200 108808 390000 108928
rect 0 107448 800 107568
rect 389200 107448 390000 107568
rect 0 106088 800 106208
rect 389200 106088 390000 106208
rect 0 104728 800 104848
rect 389200 104728 390000 104848
rect 0 103368 800 103488
rect 389200 103368 390000 103488
rect 0 102008 800 102128
rect 389200 102008 390000 102128
rect 0 100648 800 100768
rect 389200 100648 390000 100768
rect 0 99968 800 100088
rect 389200 99288 390000 99408
rect 0 98608 800 98728
rect 389200 97928 390000 98048
rect 0 97248 800 97368
rect 389200 96568 390000 96688
rect 0 95888 800 96008
rect 389200 95208 390000 95328
rect 0 94528 800 94648
rect 389200 93848 390000 93968
rect 0 93168 800 93288
rect 389200 92488 390000 92608
rect 0 91808 800 91928
rect 389200 91128 390000 91248
rect 0 90448 800 90568
rect 389200 89768 390000 89888
rect 0 89088 800 89208
rect 389200 89088 390000 89208
rect 0 87728 800 87848
rect 389200 87728 390000 87848
rect 0 86368 800 86488
rect 389200 86368 390000 86488
rect 0 85008 800 85128
rect 389200 85008 390000 85128
rect 0 83648 800 83768
rect 389200 83648 390000 83768
rect 0 82288 800 82408
rect 389200 82288 390000 82408
rect 0 80928 800 81048
rect 389200 80928 390000 81048
rect 0 79568 800 79688
rect 389200 79568 390000 79688
rect 0 78208 800 78328
rect 389200 78208 390000 78328
rect 0 76848 800 76968
rect 389200 76848 390000 76968
rect 0 75488 800 75608
rect 389200 75488 390000 75608
rect 0 74128 800 74248
rect 389200 74128 390000 74248
rect 0 72768 800 72888
rect 389200 72768 390000 72888
rect 0 71408 800 71528
rect 389200 71408 390000 71528
rect 0 70048 800 70168
rect 389200 70048 390000 70168
rect 0 68688 800 68808
rect 389200 68688 390000 68808
rect 0 67328 800 67448
rect 389200 67328 390000 67448
rect 0 65968 800 66088
rect 389200 65968 390000 66088
rect 0 64608 800 64728
rect 389200 64608 390000 64728
rect 0 63248 800 63368
rect 389200 63248 390000 63368
rect 0 61888 800 62008
rect 389200 61888 390000 62008
rect 0 60528 800 60648
rect 389200 60528 390000 60648
rect 0 59168 800 59288
rect 389200 59168 390000 59288
rect 0 57808 800 57928
rect 389200 57808 390000 57928
rect 0 56448 800 56568
rect 389200 56448 390000 56568
rect 0 55088 800 55208
rect 389200 55088 390000 55208
rect 0 53728 800 53848
rect 389200 53728 390000 53848
rect 0 52368 800 52488
rect 389200 52368 390000 52488
rect 0 51008 800 51128
rect 389200 51008 390000 51128
rect 0 49648 800 49768
rect 389200 49648 390000 49768
rect 0 48288 800 48408
rect 389200 48288 390000 48408
rect 0 46928 800 47048
rect 389200 46928 390000 47048
rect 0 45568 800 45688
rect 389200 45568 390000 45688
rect 0 44208 800 44328
rect 389200 44208 390000 44328
rect 0 42848 800 42968
rect 389200 42848 390000 42968
rect 0 41488 800 41608
rect 389200 41488 390000 41608
rect 0 40128 800 40248
rect 389200 40128 390000 40248
rect 0 38768 800 38888
rect 389200 38768 390000 38888
rect 0 37408 800 37528
rect 389200 37408 390000 37528
rect 0 36048 800 36168
rect 389200 36048 390000 36168
rect 0 34688 800 34808
rect 389200 34688 390000 34808
rect 0 33328 800 33448
rect 389200 33328 390000 33448
rect 0 31968 800 32088
rect 389200 31968 390000 32088
rect 0 30608 800 30728
rect 389200 30608 390000 30728
rect 0 29248 800 29368
rect 389200 29248 390000 29368
rect 0 27888 800 28008
rect 389200 27888 390000 28008
rect 0 26528 800 26648
rect 389200 26528 390000 26648
rect 0 25168 800 25288
rect 389200 25168 390000 25288
rect 0 23808 800 23928
rect 389200 23808 390000 23928
rect 0 22448 800 22568
rect 389200 22448 390000 22568
rect 0 21088 800 21208
rect 389200 21088 390000 21208
rect 0 19728 800 19848
rect 389200 19728 390000 19848
rect 0 18368 800 18488
rect 389200 18368 390000 18488
rect 0 17008 800 17128
rect 389200 17008 390000 17128
rect 0 15648 800 15768
rect 389200 15648 390000 15768
rect 0 14288 800 14408
rect 389200 14288 390000 14408
rect 0 12928 800 13048
rect 389200 12928 390000 13048
rect 0 11568 800 11688
rect 389200 11568 390000 11688
rect 0 10208 800 10328
rect 389200 10208 390000 10328
rect 0 8848 800 8968
rect 389200 8848 390000 8968
rect 0 7488 800 7608
rect 389200 7488 390000 7608
rect 0 6128 800 6248
rect 389200 6128 390000 6248
rect 0 4768 800 4888
rect 389200 4768 390000 4888
rect 0 3408 800 3528
rect 389200 3408 390000 3528
rect 0 2048 800 2168
rect 389200 2048 390000 2168
rect 0 688 800 808
rect 389200 688 390000 808
<< obsm3 >>
rect 880 388888 389120 389061
rect 800 387808 389200 388888
rect 880 387528 389120 387808
rect 800 386448 389200 387528
rect 880 386168 389120 386448
rect 800 385088 389200 386168
rect 880 384808 389120 385088
rect 800 383728 389200 384808
rect 880 383448 389120 383728
rect 800 382368 389200 383448
rect 880 382088 389120 382368
rect 800 381008 389200 382088
rect 880 380728 389120 381008
rect 800 379648 389200 380728
rect 880 379368 389120 379648
rect 800 378288 389200 379368
rect 880 378008 389120 378288
rect 800 376928 389200 378008
rect 880 376648 389120 376928
rect 800 375568 389200 376648
rect 880 375288 389120 375568
rect 800 374208 389200 375288
rect 880 373928 389120 374208
rect 800 372848 389200 373928
rect 880 372568 389120 372848
rect 800 371488 389200 372568
rect 880 371208 389120 371488
rect 800 370128 389200 371208
rect 880 369848 389120 370128
rect 800 368768 389200 369848
rect 880 368488 389120 368768
rect 800 367408 389200 368488
rect 880 367128 389120 367408
rect 800 366048 389200 367128
rect 880 365768 389120 366048
rect 800 364688 389200 365768
rect 880 364408 389120 364688
rect 800 363328 389200 364408
rect 880 363048 389120 363328
rect 800 361968 389200 363048
rect 880 361688 389120 361968
rect 800 360608 389200 361688
rect 880 360328 389120 360608
rect 800 359248 389200 360328
rect 880 358968 389120 359248
rect 800 357888 389200 358968
rect 880 357608 389120 357888
rect 800 356528 389200 357608
rect 880 356248 389120 356528
rect 800 355168 389200 356248
rect 880 354888 389120 355168
rect 800 353808 389200 354888
rect 880 353528 389120 353808
rect 800 352448 389200 353528
rect 880 352168 389120 352448
rect 800 351088 389200 352168
rect 880 350808 389120 351088
rect 800 349728 389200 350808
rect 880 349448 389120 349728
rect 800 348368 389200 349448
rect 880 348088 389120 348368
rect 800 347008 389200 348088
rect 880 346728 389120 347008
rect 800 345648 389200 346728
rect 880 345368 389120 345648
rect 800 344288 389200 345368
rect 880 344008 389120 344288
rect 800 342928 389200 344008
rect 880 342648 389120 342928
rect 800 341568 389200 342648
rect 880 341288 389120 341568
rect 800 340208 389200 341288
rect 880 339928 389120 340208
rect 800 338848 389200 339928
rect 880 338568 389120 338848
rect 800 337488 389200 338568
rect 880 337208 389120 337488
rect 800 336128 389200 337208
rect 880 335848 389120 336128
rect 800 334768 389200 335848
rect 880 334488 389120 334768
rect 800 333408 389200 334488
rect 880 333128 389120 333408
rect 800 332048 389200 333128
rect 880 331768 389120 332048
rect 800 330688 389200 331768
rect 880 330408 389120 330688
rect 800 329328 389200 330408
rect 880 329048 389120 329328
rect 800 327968 389200 329048
rect 880 327688 389120 327968
rect 800 326608 389200 327688
rect 880 326328 389120 326608
rect 800 325248 389200 326328
rect 880 324968 389120 325248
rect 800 323888 389200 324968
rect 880 323608 389120 323888
rect 800 322528 389200 323608
rect 880 322248 389120 322528
rect 800 321168 389200 322248
rect 880 320888 389120 321168
rect 800 319808 389200 320888
rect 880 319528 389120 319808
rect 800 318448 389200 319528
rect 880 318168 389120 318448
rect 800 317088 389200 318168
rect 880 316808 389120 317088
rect 800 315728 389200 316808
rect 880 315448 389120 315728
rect 800 314368 389200 315448
rect 880 314088 389120 314368
rect 800 313008 389200 314088
rect 880 312728 389120 313008
rect 800 311648 389200 312728
rect 880 311368 389120 311648
rect 800 310288 389200 311368
rect 880 310008 389120 310288
rect 800 308928 389200 310008
rect 880 308648 389120 308928
rect 800 307568 389200 308648
rect 880 307288 389120 307568
rect 800 306208 389200 307288
rect 880 305928 389120 306208
rect 800 304848 389200 305928
rect 880 304568 389120 304848
rect 800 303488 389200 304568
rect 880 303208 389120 303488
rect 800 302128 389200 303208
rect 880 301848 389120 302128
rect 800 300768 389200 301848
rect 880 300488 389120 300768
rect 800 300088 389200 300488
rect 880 299808 389200 300088
rect 800 299408 389200 299808
rect 800 299128 389120 299408
rect 800 298728 389200 299128
rect 880 298448 389200 298728
rect 800 298048 389200 298448
rect 800 297768 389120 298048
rect 800 297368 389200 297768
rect 880 297088 389200 297368
rect 800 296688 389200 297088
rect 800 296408 389120 296688
rect 800 296008 389200 296408
rect 880 295728 389200 296008
rect 800 295328 389200 295728
rect 800 295048 389120 295328
rect 800 294648 389200 295048
rect 880 294368 389200 294648
rect 800 293968 389200 294368
rect 800 293688 389120 293968
rect 800 293288 389200 293688
rect 880 293008 389200 293288
rect 800 292608 389200 293008
rect 800 292328 389120 292608
rect 800 291928 389200 292328
rect 880 291648 389200 291928
rect 800 291248 389200 291648
rect 800 290968 389120 291248
rect 800 290568 389200 290968
rect 880 290288 389200 290568
rect 800 289888 389200 290288
rect 800 289608 389120 289888
rect 800 289208 389200 289608
rect 880 288928 389120 289208
rect 800 287848 389200 288928
rect 880 287568 389120 287848
rect 800 286488 389200 287568
rect 880 286208 389120 286488
rect 800 285128 389200 286208
rect 880 284848 389120 285128
rect 800 283768 389200 284848
rect 880 283488 389120 283768
rect 800 282408 389200 283488
rect 880 282128 389120 282408
rect 800 281048 389200 282128
rect 880 280768 389120 281048
rect 800 279688 389200 280768
rect 880 279408 389120 279688
rect 800 278328 389200 279408
rect 880 278048 389120 278328
rect 800 276968 389200 278048
rect 880 276688 389120 276968
rect 800 275608 389200 276688
rect 880 275328 389120 275608
rect 800 274248 389200 275328
rect 880 273968 389120 274248
rect 800 272888 389200 273968
rect 880 272608 389120 272888
rect 800 271528 389200 272608
rect 880 271248 389120 271528
rect 800 270168 389200 271248
rect 880 269888 389120 270168
rect 800 268808 389200 269888
rect 880 268528 389120 268808
rect 800 267448 389200 268528
rect 880 267168 389120 267448
rect 800 266088 389200 267168
rect 880 265808 389120 266088
rect 800 264728 389200 265808
rect 880 264448 389120 264728
rect 800 263368 389200 264448
rect 880 263088 389120 263368
rect 800 262008 389200 263088
rect 880 261728 389120 262008
rect 800 260648 389200 261728
rect 880 260368 389120 260648
rect 800 259288 389200 260368
rect 880 259008 389120 259288
rect 800 257928 389200 259008
rect 880 257648 389120 257928
rect 800 256568 389200 257648
rect 880 256288 389120 256568
rect 800 255208 389200 256288
rect 880 254928 389120 255208
rect 800 253848 389200 254928
rect 880 253568 389120 253848
rect 800 252488 389200 253568
rect 880 252208 389120 252488
rect 800 251128 389200 252208
rect 880 250848 389120 251128
rect 800 249768 389200 250848
rect 880 249488 389120 249768
rect 800 248408 389200 249488
rect 880 248128 389120 248408
rect 800 247048 389200 248128
rect 880 246768 389120 247048
rect 800 245688 389200 246768
rect 880 245408 389120 245688
rect 800 244328 389200 245408
rect 880 244048 389120 244328
rect 800 242968 389200 244048
rect 880 242688 389120 242968
rect 800 241608 389200 242688
rect 880 241328 389120 241608
rect 800 240248 389200 241328
rect 880 239968 389120 240248
rect 800 238888 389200 239968
rect 880 238608 389120 238888
rect 800 237528 389200 238608
rect 880 237248 389120 237528
rect 800 236168 389200 237248
rect 880 235888 389120 236168
rect 800 234808 389200 235888
rect 880 234528 389120 234808
rect 800 233448 389200 234528
rect 880 233168 389120 233448
rect 800 232088 389200 233168
rect 880 231808 389120 232088
rect 800 230728 389200 231808
rect 880 230448 389120 230728
rect 800 229368 389200 230448
rect 880 229088 389120 229368
rect 800 228008 389200 229088
rect 880 227728 389120 228008
rect 800 226648 389200 227728
rect 880 226368 389120 226648
rect 800 225288 389200 226368
rect 880 225008 389120 225288
rect 800 223928 389200 225008
rect 880 223648 389120 223928
rect 800 222568 389200 223648
rect 880 222288 389120 222568
rect 800 221208 389200 222288
rect 880 220928 389120 221208
rect 800 219848 389200 220928
rect 880 219568 389120 219848
rect 800 218488 389200 219568
rect 880 218208 389120 218488
rect 800 217128 389200 218208
rect 880 216848 389120 217128
rect 800 215768 389200 216848
rect 880 215488 389120 215768
rect 800 214408 389200 215488
rect 880 214128 389120 214408
rect 800 213048 389200 214128
rect 880 212768 389120 213048
rect 800 211688 389200 212768
rect 880 211408 389120 211688
rect 800 210328 389200 211408
rect 880 210048 389120 210328
rect 800 208968 389200 210048
rect 880 208688 389120 208968
rect 800 207608 389200 208688
rect 880 207328 389120 207608
rect 800 206248 389200 207328
rect 880 205968 389120 206248
rect 800 204888 389200 205968
rect 880 204608 389120 204888
rect 800 203528 389200 204608
rect 880 203248 389120 203528
rect 800 202168 389200 203248
rect 880 201888 389120 202168
rect 800 200808 389200 201888
rect 880 200528 389120 200808
rect 800 200128 389200 200528
rect 880 199848 389200 200128
rect 800 199448 389200 199848
rect 800 199168 389120 199448
rect 800 198768 389200 199168
rect 880 198488 389200 198768
rect 800 198088 389200 198488
rect 800 197808 389120 198088
rect 800 197408 389200 197808
rect 880 197128 389200 197408
rect 800 196728 389200 197128
rect 800 196448 389120 196728
rect 800 196048 389200 196448
rect 880 195768 389200 196048
rect 800 195368 389200 195768
rect 800 195088 389120 195368
rect 800 194688 389200 195088
rect 880 194408 389200 194688
rect 800 194008 389200 194408
rect 800 193728 389120 194008
rect 800 193328 389200 193728
rect 880 193048 389200 193328
rect 800 192648 389200 193048
rect 800 192368 389120 192648
rect 800 191968 389200 192368
rect 880 191688 389200 191968
rect 800 191288 389200 191688
rect 800 191008 389120 191288
rect 800 190608 389200 191008
rect 880 190328 389200 190608
rect 800 189928 389200 190328
rect 800 189648 389120 189928
rect 800 189248 389200 189648
rect 880 188968 389120 189248
rect 800 187888 389200 188968
rect 880 187608 389120 187888
rect 800 186528 389200 187608
rect 880 186248 389120 186528
rect 800 185168 389200 186248
rect 880 184888 389120 185168
rect 800 183808 389200 184888
rect 880 183528 389120 183808
rect 800 182448 389200 183528
rect 880 182168 389120 182448
rect 800 181088 389200 182168
rect 880 180808 389120 181088
rect 800 179728 389200 180808
rect 880 179448 389120 179728
rect 800 178368 389200 179448
rect 880 178088 389120 178368
rect 800 177008 389200 178088
rect 880 176728 389120 177008
rect 800 175648 389200 176728
rect 880 175368 389120 175648
rect 800 174288 389200 175368
rect 880 174008 389120 174288
rect 800 172928 389200 174008
rect 880 172648 389120 172928
rect 800 171568 389200 172648
rect 880 171288 389120 171568
rect 800 170208 389200 171288
rect 880 169928 389120 170208
rect 800 168848 389200 169928
rect 880 168568 389120 168848
rect 800 167488 389200 168568
rect 880 167208 389120 167488
rect 800 166128 389200 167208
rect 880 165848 389120 166128
rect 800 164768 389200 165848
rect 880 164488 389120 164768
rect 800 163408 389200 164488
rect 880 163128 389120 163408
rect 800 162048 389200 163128
rect 880 161768 389120 162048
rect 800 160688 389200 161768
rect 880 160408 389120 160688
rect 800 159328 389200 160408
rect 880 159048 389120 159328
rect 800 157968 389200 159048
rect 880 157688 389120 157968
rect 800 156608 389200 157688
rect 880 156328 389120 156608
rect 800 155248 389200 156328
rect 880 154968 389120 155248
rect 800 153888 389200 154968
rect 880 153608 389120 153888
rect 800 152528 389200 153608
rect 880 152248 389120 152528
rect 800 151168 389200 152248
rect 880 150888 389120 151168
rect 800 149808 389200 150888
rect 880 149528 389120 149808
rect 800 148448 389200 149528
rect 880 148168 389120 148448
rect 800 147088 389200 148168
rect 880 146808 389120 147088
rect 800 145728 389200 146808
rect 880 145448 389120 145728
rect 800 144368 389200 145448
rect 880 144088 389120 144368
rect 800 143008 389200 144088
rect 880 142728 389120 143008
rect 800 141648 389200 142728
rect 880 141368 389120 141648
rect 800 140288 389200 141368
rect 880 140008 389120 140288
rect 800 138928 389200 140008
rect 880 138648 389120 138928
rect 800 137568 389200 138648
rect 880 137288 389120 137568
rect 800 136208 389200 137288
rect 880 135928 389120 136208
rect 800 134848 389200 135928
rect 880 134568 389120 134848
rect 800 133488 389200 134568
rect 880 133208 389120 133488
rect 800 132128 389200 133208
rect 880 131848 389120 132128
rect 800 130768 389200 131848
rect 880 130488 389120 130768
rect 800 129408 389200 130488
rect 880 129128 389120 129408
rect 800 128048 389200 129128
rect 880 127768 389120 128048
rect 800 126688 389200 127768
rect 880 126408 389120 126688
rect 800 125328 389200 126408
rect 880 125048 389120 125328
rect 800 123968 389200 125048
rect 880 123688 389120 123968
rect 800 122608 389200 123688
rect 880 122328 389120 122608
rect 800 121248 389200 122328
rect 880 120968 389120 121248
rect 800 119888 389200 120968
rect 880 119608 389120 119888
rect 800 118528 389200 119608
rect 880 118248 389120 118528
rect 800 117168 389200 118248
rect 880 116888 389120 117168
rect 800 115808 389200 116888
rect 880 115528 389120 115808
rect 800 114448 389200 115528
rect 880 114168 389120 114448
rect 800 113088 389200 114168
rect 880 112808 389120 113088
rect 800 111728 389200 112808
rect 880 111448 389120 111728
rect 800 110368 389200 111448
rect 880 110088 389120 110368
rect 800 109008 389200 110088
rect 880 108728 389120 109008
rect 800 107648 389200 108728
rect 880 107368 389120 107648
rect 800 106288 389200 107368
rect 880 106008 389120 106288
rect 800 104928 389200 106008
rect 880 104648 389120 104928
rect 800 103568 389200 104648
rect 880 103288 389120 103568
rect 800 102208 389200 103288
rect 880 101928 389120 102208
rect 800 100848 389200 101928
rect 880 100568 389120 100848
rect 800 100168 389200 100568
rect 880 99888 389200 100168
rect 800 99488 389200 99888
rect 800 99208 389120 99488
rect 800 98808 389200 99208
rect 880 98528 389200 98808
rect 800 98128 389200 98528
rect 800 97848 389120 98128
rect 800 97448 389200 97848
rect 880 97168 389200 97448
rect 800 96768 389200 97168
rect 800 96488 389120 96768
rect 800 96088 389200 96488
rect 880 95808 389200 96088
rect 800 95408 389200 95808
rect 800 95128 389120 95408
rect 800 94728 389200 95128
rect 880 94448 389200 94728
rect 800 94048 389200 94448
rect 800 93768 389120 94048
rect 800 93368 389200 93768
rect 880 93088 389200 93368
rect 800 92688 389200 93088
rect 800 92408 389120 92688
rect 800 92008 389200 92408
rect 880 91728 389200 92008
rect 800 91328 389200 91728
rect 800 91048 389120 91328
rect 800 90648 389200 91048
rect 880 90368 389200 90648
rect 800 89968 389200 90368
rect 800 89688 389120 89968
rect 800 89288 389200 89688
rect 880 89008 389120 89288
rect 800 87928 389200 89008
rect 880 87648 389120 87928
rect 800 86568 389200 87648
rect 880 86288 389120 86568
rect 800 85208 389200 86288
rect 880 84928 389120 85208
rect 800 83848 389200 84928
rect 880 83568 389120 83848
rect 800 82488 389200 83568
rect 880 82208 389120 82488
rect 800 81128 389200 82208
rect 880 80848 389120 81128
rect 800 79768 389200 80848
rect 880 79488 389120 79768
rect 800 78408 389200 79488
rect 880 78128 389120 78408
rect 800 77048 389200 78128
rect 880 76768 389120 77048
rect 800 75688 389200 76768
rect 880 75408 389120 75688
rect 800 74328 389200 75408
rect 880 74048 389120 74328
rect 800 72968 389200 74048
rect 880 72688 389120 72968
rect 800 71608 389200 72688
rect 880 71328 389120 71608
rect 800 70248 389200 71328
rect 880 69968 389120 70248
rect 800 68888 389200 69968
rect 880 68608 389120 68888
rect 800 67528 389200 68608
rect 880 67248 389120 67528
rect 800 66168 389200 67248
rect 880 65888 389120 66168
rect 800 64808 389200 65888
rect 880 64528 389120 64808
rect 800 63448 389200 64528
rect 880 63168 389120 63448
rect 800 62088 389200 63168
rect 880 61808 389120 62088
rect 800 60728 389200 61808
rect 880 60448 389120 60728
rect 800 59368 389200 60448
rect 880 59088 389120 59368
rect 800 58008 389200 59088
rect 880 57728 389120 58008
rect 800 56648 389200 57728
rect 880 56368 389120 56648
rect 800 55288 389200 56368
rect 880 55008 389120 55288
rect 800 53928 389200 55008
rect 880 53648 389120 53928
rect 800 52568 389200 53648
rect 880 52288 389120 52568
rect 800 51208 389200 52288
rect 880 50928 389120 51208
rect 800 49848 389200 50928
rect 880 49568 389120 49848
rect 800 48488 389200 49568
rect 880 48208 389120 48488
rect 800 47128 389200 48208
rect 880 46848 389120 47128
rect 800 45768 389200 46848
rect 880 45488 389120 45768
rect 800 44408 389200 45488
rect 880 44128 389120 44408
rect 800 43048 389200 44128
rect 880 42768 389120 43048
rect 800 41688 389200 42768
rect 880 41408 389120 41688
rect 800 40328 389200 41408
rect 880 40048 389120 40328
rect 800 38968 389200 40048
rect 880 38688 389120 38968
rect 800 37608 389200 38688
rect 880 37328 389120 37608
rect 800 36248 389200 37328
rect 880 35968 389120 36248
rect 800 34888 389200 35968
rect 880 34608 389120 34888
rect 800 33528 389200 34608
rect 880 33248 389120 33528
rect 800 32168 389200 33248
rect 880 31888 389120 32168
rect 800 30808 389200 31888
rect 880 30528 389120 30808
rect 800 29448 389200 30528
rect 880 29168 389120 29448
rect 800 28088 389200 29168
rect 880 27808 389120 28088
rect 800 26728 389200 27808
rect 880 26448 389120 26728
rect 800 25368 389200 26448
rect 880 25088 389120 25368
rect 800 24008 389200 25088
rect 880 23728 389120 24008
rect 800 22648 389200 23728
rect 880 22368 389120 22648
rect 800 21288 389200 22368
rect 880 21008 389120 21288
rect 800 19928 389200 21008
rect 880 19648 389120 19928
rect 800 18568 389200 19648
rect 880 18288 389120 18568
rect 800 17208 389200 18288
rect 880 16928 389120 17208
rect 800 15848 389200 16928
rect 880 15568 389120 15848
rect 800 14488 389200 15568
rect 880 14208 389120 14488
rect 800 13128 389200 14208
rect 880 12848 389120 13128
rect 800 11768 389200 12848
rect 880 11488 389120 11768
rect 800 10408 389200 11488
rect 880 10128 389120 10408
rect 800 9048 389200 10128
rect 880 8768 389120 9048
rect 800 7688 389200 8768
rect 880 7408 389120 7688
rect 800 6328 389200 7408
rect 880 6048 389120 6328
rect 800 4968 389200 6048
rect 880 4688 389120 4968
rect 800 3608 389200 4688
rect 880 3328 389120 3608
rect 800 2248 389200 3328
rect 880 2075 389120 2248
<< metal4 >>
rect 4208 2128 4528 387376
rect 19568 2128 19888 387376
rect 34928 2128 35248 387376
rect 50288 2128 50608 387376
rect 65648 2128 65968 387376
rect 81008 2128 81328 387376
rect 96368 2128 96688 387376
rect 111728 2128 112048 387376
rect 127088 2128 127408 387376
rect 142448 2128 142768 387376
rect 157808 2128 158128 387376
rect 173168 2128 173488 387376
rect 188528 2128 188848 387376
rect 203888 2128 204208 387376
rect 219248 2128 219568 387376
rect 234608 2128 234928 387376
rect 249968 2128 250288 387376
rect 265328 2128 265648 387376
rect 280688 2128 281008 387376
rect 296048 2128 296368 387376
rect 311408 2128 311728 387376
rect 326768 2128 327088 387376
rect 342128 2128 342448 387376
rect 357488 2128 357808 387376
rect 372848 2128 373168 387376
rect 388208 2128 388528 387376
<< obsm4 >>
rect 12203 2347 19488 387021
rect 19968 2347 34848 387021
rect 35328 2347 50208 387021
rect 50688 2347 65568 387021
rect 66048 2347 80928 387021
rect 81408 2347 96288 387021
rect 96768 2347 111648 387021
rect 112128 2347 127008 387021
rect 127488 2347 142368 387021
rect 142848 2347 157728 387021
rect 158208 2347 173088 387021
rect 173568 2347 188448 387021
rect 188928 2347 203808 387021
rect 204288 2347 219168 387021
rect 219648 2347 234528 387021
rect 235008 2347 249888 387021
rect 250368 2347 265248 387021
rect 265728 2347 280608 387021
rect 281088 2347 295968 387021
rect 296448 2347 311328 387021
rect 311808 2347 326688 387021
rect 327168 2347 342048 387021
rect 342528 2347 356165 387021
<< labels >>
rlabel metal3 s 389200 201968 390000 202088 6 clk
port 1 nsew signal input
rlabel metal3 s 389200 121048 390000 121168 6 dcache_data_chip_en_1
port 2 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 dcache_data_chip_en_2
port 3 nsew signal input
rlabel metal3 s 0 376728 800 376848 6 dcache_data_in_1[0]
port 4 nsew signal input
rlabel metal3 s 389200 222368 390000 222488 6 dcache_data_in_1[10]
port 5 nsew signal input
rlabel metal2 s 144274 389200 144330 390000 6 dcache_data_in_1[11]
port 6 nsew signal input
rlabel metal3 s 0 255008 800 255128 6 dcache_data_in_1[12]
port 7 nsew signal input
rlabel metal2 s 123666 389200 123722 390000 6 dcache_data_in_1[13]
port 8 nsew signal input
rlabel metal2 s 222198 389200 222254 390000 6 dcache_data_in_1[14]
port 9 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 dcache_data_in_1[15]
port 10 nsew signal input
rlabel metal2 s 267278 0 267334 800 6 dcache_data_in_1[16]
port 11 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 dcache_data_in_1[17]
port 12 nsew signal input
rlabel metal2 s 47030 389200 47086 390000 6 dcache_data_in_1[18]
port 13 nsew signal input
rlabel metal2 s 194506 389200 194562 390000 6 dcache_data_in_1[19]
port 14 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 dcache_data_in_1[1]
port 15 nsew signal input
rlabel metal2 s 378690 389200 378746 390000 6 dcache_data_in_1[20]
port 16 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 dcache_data_in_1[21]
port 17 nsew signal input
rlabel metal2 s 189354 389200 189410 390000 6 dcache_data_in_1[22]
port 18 nsew signal input
rlabel metal2 s 97262 389200 97318 390000 6 dcache_data_in_1[23]
port 19 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 dcache_data_in_1[24]
port 20 nsew signal input
rlabel metal3 s 0 356328 800 356448 6 dcache_data_in_1[25]
port 21 nsew signal input
rlabel metal2 s 214470 389200 214526 390000 6 dcache_data_in_1[26]
port 22 nsew signal input
rlabel metal2 s 220910 0 220966 800 6 dcache_data_in_1[27]
port 23 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 dcache_data_in_1[28]
port 24 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 dcache_data_in_1[29]
port 25 nsew signal input
rlabel metal3 s 389200 199248 390000 199368 6 dcache_data_in_1[2]
port 26 nsew signal input
rlabel metal2 s 387062 0 387118 800 6 dcache_data_in_1[30]
port 27 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 dcache_data_in_1[31]
port 28 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 dcache_data_in_1[3]
port 29 nsew signal input
rlabel metal3 s 0 315528 800 315648 6 dcache_data_in_1[4]
port 30 nsew signal input
rlabel metal2 s 294970 0 295026 800 6 dcache_data_in_1[5]
port 31 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 dcache_data_in_1[6]
port 32 nsew signal input
rlabel metal3 s 389200 278128 390000 278248 6 dcache_data_in_1[7]
port 33 nsew signal input
rlabel metal2 s 253110 0 253166 800 6 dcache_data_in_1[8]
port 34 nsew signal input
rlabel metal2 s 110786 389200 110842 390000 6 dcache_data_in_1[9]
port 35 nsew signal input
rlabel metal3 s 389200 244128 390000 244248 6 dcache_data_in_2[0]
port 36 nsew signal input
rlabel metal3 s 0 268608 800 268728 6 dcache_data_in_2[10]
port 37 nsew signal input
rlabel metal3 s 389200 130568 390000 130688 6 dcache_data_in_2[11]
port 38 nsew signal input
rlabel metal2 s 363234 389200 363290 390000 6 dcache_data_in_2[12]
port 39 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 dcache_data_in_2[13]
port 40 nsew signal input
rlabel metal3 s 0 289008 800 289128 6 dcache_data_in_2[14]
port 41 nsew signal input
rlabel metal2 s 152002 389200 152058 390000 6 dcache_data_in_2[15]
port 42 nsew signal input
rlabel metal2 s 272430 389200 272486 390000 6 dcache_data_in_2[16]
port 43 nsew signal input
rlabel metal3 s 389200 103368 390000 103488 6 dcache_data_in_2[17]
port 44 nsew signal input
rlabel metal3 s 0 352248 800 352368 6 dcache_data_in_2[18]
port 45 nsew signal input
rlabel metal3 s 389200 30608 390000 30728 6 dcache_data_in_2[19]
port 46 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 dcache_data_in_2[1]
port 47 nsew signal input
rlabel metal3 s 389200 323688 390000 323808 6 dcache_data_in_2[20]
port 48 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 dcache_data_in_2[21]
port 49 nsew signal input
rlabel metal2 s 88246 389200 88302 390000 6 dcache_data_in_2[22]
port 50 nsew signal input
rlabel metal3 s 389200 95208 390000 95328 6 dcache_data_in_2[23]
port 51 nsew signal input
rlabel metal3 s 389200 314168 390000 314288 6 dcache_data_in_2[24]
port 52 nsew signal input
rlabel metal2 s 136546 389200 136602 390000 6 dcache_data_in_2[25]
port 53 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 dcache_data_in_2[26]
port 54 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 dcache_data_in_2[27]
port 55 nsew signal input
rlabel metal3 s 389200 65968 390000 66088 6 dcache_data_in_2[28]
port 56 nsew signal input
rlabel metal3 s 389200 60528 390000 60648 6 dcache_data_in_2[29]
port 57 nsew signal input
rlabel metal2 s 140410 389200 140466 390000 6 dcache_data_in_2[2]
port 58 nsew signal input
rlabel metal3 s 0 223728 800 223848 6 dcache_data_in_2[30]
port 59 nsew signal input
rlabel metal2 s 262126 389200 262182 390000 6 dcache_data_in_2[31]
port 60 nsew signal input
rlabel metal2 s 228638 389200 228694 390000 6 dcache_data_in_2[3]
port 61 nsew signal input
rlabel metal3 s 0 340008 800 340128 6 dcache_data_in_2[4]
port 62 nsew signal input
rlabel metal2 s 290462 389200 290518 390000 6 dcache_data_in_2[5]
port 63 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 dcache_data_in_2[6]
port 64 nsew signal input
rlabel metal3 s 0 300568 800 300688 6 dcache_data_in_2[7]
port 65 nsew signal input
rlabel metal2 s 206742 389200 206798 390000 6 dcache_data_in_2[8]
port 66 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 dcache_data_in_2[9]
port 67 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 dcache_data_index_1[0]
port 68 nsew signal input
rlabel metal3 s 389200 350888 390000 351008 6 dcache_data_index_1[1]
port 69 nsew signal input
rlabel metal2 s 373538 0 373594 800 6 dcache_data_index_1[2]
port 70 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 dcache_data_index_1[3]
port 71 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 dcache_data_index_1[4]
port 72 nsew signal input
rlabel metal3 s 389200 380808 390000 380928 6 dcache_data_index_1[5]
port 73 nsew signal input
rlabel metal2 s 161018 389200 161074 390000 6 dcache_data_index_1[6]
port 74 nsew signal input
rlabel metal2 s 48318 389200 48374 390000 6 dcache_data_index_1[7]
port 75 nsew signal input
rlabel metal2 s 149426 389200 149482 390000 6 dcache_data_index_2[0]
port 76 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 dcache_data_index_2[1]
port 77 nsew signal input
rlabel metal3 s 389200 116968 390000 117088 6 dcache_data_index_2[2]
port 78 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 dcache_data_index_2[3]
port 79 nsew signal input
rlabel metal2 s 309138 389200 309194 390000 6 dcache_data_index_2[4]
port 80 nsew signal input
rlabel metal2 s 241518 0 241574 800 6 dcache_data_index_2[5]
port 81 nsew signal input
rlabel metal2 s 71502 389200 71558 390000 6 dcache_data_index_2[6]
port 82 nsew signal input
rlabel metal3 s 389200 284928 390000 285048 6 dcache_data_index_2[7]
port 83 nsew signal input
rlabel metal2 s 132682 389200 132738 390000 6 dcache_data_out_1[0]
port 84 nsew signal output
rlabel metal2 s 197082 389200 197138 390000 6 dcache_data_out_1[10]
port 85 nsew signal output
rlabel metal3 s 0 311448 800 311568 6 dcache_data_out_1[11]
port 86 nsew signal output
rlabel metal2 s 328458 0 328514 800 6 dcache_data_out_1[12]
port 87 nsew signal output
rlabel metal3 s 0 335928 800 336048 6 dcache_data_out_1[13]
port 88 nsew signal output
rlabel metal2 s 218334 0 218390 800 6 dcache_data_out_1[14]
port 89 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 dcache_data_out_1[15]
port 90 nsew signal output
rlabel metal3 s 389200 311448 390000 311568 6 dcache_data_out_1[16]
port 91 nsew signal output
rlabel metal3 s 0 260448 800 260568 6 dcache_data_out_1[17]
port 92 nsew signal output
rlabel metal3 s 0 219648 800 219768 6 dcache_data_out_1[18]
port 93 nsew signal output
rlabel metal2 s 39302 389200 39358 390000 6 dcache_data_out_1[19]
port 94 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 dcache_data_out_1[1]
port 95 nsew signal output
rlabel metal3 s 389200 319608 390000 319728 6 dcache_data_out_1[20]
port 96 nsew signal output
rlabel metal3 s 389200 153688 390000 153808 6 dcache_data_out_1[21]
port 97 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 dcache_data_out_1[22]
port 98 nsew signal output
rlabel metal2 s 287242 0 287298 800 6 dcache_data_out_1[23]
port 99 nsew signal output
rlabel metal2 s 332322 0 332378 800 6 dcache_data_out_1[24]
port 100 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 dcache_data_out_1[25]
port 101 nsew signal output
rlabel metal3 s 389200 165928 390000 166048 6 dcache_data_out_1[26]
port 102 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 dcache_data_out_1[27]
port 103 nsew signal output
rlabel metal2 s 311714 389200 311770 390000 6 dcache_data_out_1[28]
port 104 nsew signal output
rlabel metal2 s 220910 389200 220966 390000 6 dcache_data_out_1[29]
port 105 nsew signal output
rlabel metal3 s 389200 329128 390000 329248 6 dcache_data_out_1[2]
port 106 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 dcache_data_out_1[30]
port 107 nsew signal output
rlabel metal3 s 389200 134648 390000 134768 6 dcache_data_out_1[31]
port 108 nsew signal output
rlabel metal2 s 18 389200 74 390000 6 dcache_data_out_1[3]
port 109 nsew signal output
rlabel metal3 s 389200 348168 390000 348288 6 dcache_data_out_1[4]
port 110 nsew signal output
rlabel metal2 s 189998 0 190054 800 6 dcache_data_out_1[5]
port 111 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 dcache_data_out_1[6]
port 112 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 dcache_data_out_1[7]
port 113 nsew signal output
rlabel metal2 s 388350 0 388406 800 6 dcache_data_out_1[8]
port 114 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 dcache_data_out_1[9]
port 115 nsew signal output
rlabel metal3 s 0 210128 800 210248 6 dcache_data_out_2[0]
port 116 nsew signal output
rlabel metal3 s 389200 76848 390000 76968 6 dcache_data_out_2[10]
port 117 nsew signal output
rlabel metal3 s 0 331848 800 331968 6 dcache_data_out_2[11]
port 118 nsew signal output
rlabel metal3 s 389200 331848 390000 331968 6 dcache_data_out_2[12]
port 119 nsew signal output
rlabel metal3 s 389200 263168 390000 263288 6 dcache_data_out_2[13]
port 120 nsew signal output
rlabel metal2 s 65062 389200 65118 390000 6 dcache_data_out_2[14]
port 121 nsew signal output
rlabel metal2 s 80518 389200 80574 390000 6 dcache_data_out_2[15]
port 122 nsew signal output
rlabel metal3 s 389200 107448 390000 107568 6 dcache_data_out_2[16]
port 123 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 dcache_data_out_2[17]
port 124 nsew signal output
rlabel metal3 s 389200 233248 390000 233368 6 dcache_data_out_2[18]
port 125 nsew signal output
rlabel metal2 s 242806 389200 242862 390000 6 dcache_data_out_2[19]
port 126 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 dcache_data_out_2[1]
port 127 nsew signal output
rlabel metal2 s 99838 389200 99894 390000 6 dcache_data_out_2[20]
port 128 nsew signal output
rlabel metal2 s 369674 389200 369730 390000 6 dcache_data_out_2[21]
port 129 nsew signal output
rlabel metal2 s 217046 389200 217102 390000 6 dcache_data_out_2[22]
port 130 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 dcache_data_out_2[23]
port 131 nsew signal output
rlabel metal2 s 367098 389200 367154 390000 6 dcache_data_out_2[24]
port 132 nsew signal output
rlabel metal2 s 662 0 718 800 6 dcache_data_out_2[25]
port 133 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 dcache_data_out_2[26]
port 134 nsew signal output
rlabel metal3 s 389200 89088 390000 89208 6 dcache_data_out_2[27]
port 135 nsew signal output
rlabel metal2 s 184202 0 184258 800 6 dcache_data_out_2[28]
port 136 nsew signal output
rlabel metal3 s 0 195848 800 195968 6 dcache_data_out_2[29]
port 137 nsew signal output
rlabel metal3 s 389200 25168 390000 25288 6 dcache_data_out_2[2]
port 138 nsew signal output
rlabel metal2 s 98550 389200 98606 390000 6 dcache_data_out_2[30]
port 139 nsew signal output
rlabel metal2 s 9034 389200 9090 390000 6 dcache_data_out_2[31]
port 140 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 dcache_data_out_2[3]
port 141 nsew signal output
rlabel metal3 s 0 159128 800 159248 6 dcache_data_out_2[4]
port 142 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 dcache_data_out_2[5]
port 143 nsew signal output
rlabel metal2 s 75366 389200 75422 390000 6 dcache_data_out_2[6]
port 144 nsew signal output
rlabel metal3 s 389200 345448 390000 345568 6 dcache_data_out_2[7]
port 145 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 dcache_data_out_2[8]
port 146 nsew signal output
rlabel metal3 s 0 357688 800 357808 6 dcache_data_out_2[9]
port 147 nsew signal output
rlabel metal3 s 389200 267248 390000 267368 6 dcache_data_write_en_1
port 148 nsew signal input
rlabel metal2 s 72790 389200 72846 390000 6 dcache_data_write_en_2
port 149 nsew signal input
rlabel metal2 s 342626 0 342682 800 6 dcache_tag_chip_en
port 150 nsew signal input
rlabel metal3 s 389200 46928 390000 47048 6 dcache_tag_data_in[0]
port 151 nsew signal input
rlabel metal2 s 26422 389200 26478 390000 6 dcache_tag_data_in[10]
port 152 nsew signal input
rlabel metal2 s 359370 0 359426 800 6 dcache_tag_data_in[11]
port 153 nsew signal input
rlabel metal3 s 389200 123768 390000 123888 6 dcache_tag_data_in[12]
port 154 nsew signal input
rlabel metal2 s 292394 0 292450 800 6 dcache_tag_data_in[13]
port 155 nsew signal input
rlabel metal2 s 150714 389200 150770 390000 6 dcache_tag_data_in[14]
port 156 nsew signal input
rlabel metal3 s 0 225088 800 225208 6 dcache_tag_data_in[15]
port 157 nsew signal input
rlabel metal3 s 0 203328 800 203448 6 dcache_tag_data_in[16]
port 158 nsew signal input
rlabel metal3 s 389200 231888 390000 232008 6 dcache_tag_data_in[17]
port 159 nsew signal input
rlabel metal3 s 389200 249568 390000 249688 6 dcache_tag_data_in[18]
port 160 nsew signal input
rlabel metal2 s 109498 389200 109554 390000 6 dcache_tag_data_in[19]
port 161 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 dcache_tag_data_in[1]
port 162 nsew signal input
rlabel metal2 s 105634 389200 105690 390000 6 dcache_tag_data_in[20]
port 163 nsew signal input
rlabel metal2 s 385774 0 385830 800 6 dcache_tag_data_in[21]
port 164 nsew signal input
rlabel metal3 s 389200 306008 390000 306128 6 dcache_tag_data_in[22]
port 165 nsew signal input
rlabel metal2 s 320730 389200 320786 390000 6 dcache_tag_data_in[23]
port 166 nsew signal input
rlabel metal3 s 0 348168 800 348288 6 dcache_tag_data_in[24]
port 167 nsew signal input
rlabel metal3 s 389200 10208 390000 10328 6 dcache_tag_data_in[25]
port 168 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 dcache_tag_data_in[26]
port 169 nsew signal input
rlabel metal2 s 334898 0 334954 800 6 dcache_tag_data_in[27]
port 170 nsew signal input
rlabel metal3 s 389200 248208 390000 248328 6 dcache_tag_data_in[28]
port 171 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 dcache_tag_data_in[29]
port 172 nsew signal input
rlabel metal3 s 0 338648 800 338768 6 dcache_tag_data_in[2]
port 173 nsew signal input
rlabel metal3 s 389200 320968 390000 321088 6 dcache_tag_data_in[30]
port 174 nsew signal input
rlabel metal2 s 175186 389200 175242 390000 6 dcache_tag_data_in[31]
port 175 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 dcache_tag_data_in[3]
port 176 nsew signal input
rlabel metal3 s 0 249568 800 249688 6 dcache_tag_data_in[4]
port 177 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 dcache_tag_data_in[5]
port 178 nsew signal input
rlabel metal3 s 0 246848 800 246968 6 dcache_tag_data_in[6]
port 179 nsew signal input
rlabel metal3 s 0 241408 800 241528 6 dcache_tag_data_in[7]
port 180 nsew signal input
rlabel metal2 s 253110 389200 253166 390000 6 dcache_tag_data_in[8]
port 181 nsew signal input
rlabel metal3 s 0 344088 800 344208 6 dcache_tag_data_in[9]
port 182 nsew signal input
rlabel metal2 s 117226 389200 117282 390000 6 dcache_tag_index[0]
port 183 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 dcache_tag_index[1]
port 184 nsew signal input
rlabel metal3 s 389200 338648 390000 338768 6 dcache_tag_index[2]
port 185 nsew signal input
rlabel metal3 s 389200 322328 390000 322448 6 dcache_tag_index[3]
port 186 nsew signal input
rlabel metal3 s 0 346808 800 346928 6 dcache_tag_index[4]
port 187 nsew signal input
rlabel metal3 s 0 341368 800 341488 6 dcache_tag_index[5]
port 188 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 dcache_tag_index[6]
port 189 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 dcache_tag_index[7]
port 190 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 dcache_tag_out[0]
port 191 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 dcache_tag_out[10]
port 192 nsew signal output
rlabel metal2 s 135258 389200 135314 390000 6 dcache_tag_out[11]
port 193 nsew signal output
rlabel metal3 s 389200 78208 390000 78328 6 dcache_tag_out[12]
port 194 nsew signal output
rlabel metal2 s 276294 389200 276350 390000 6 dcache_tag_out[13]
port 195 nsew signal output
rlabel metal2 s 329746 389200 329802 390000 6 dcache_tag_out[14]
port 196 nsew signal output
rlabel metal3 s 389200 6128 390000 6248 6 dcache_tag_out[15]
port 197 nsew signal output
rlabel metal2 s 199658 389200 199714 390000 6 dcache_tag_out[16]
port 198 nsew signal output
rlabel metal2 s 50894 389200 50950 390000 6 dcache_tag_out[17]
port 199 nsew signal output
rlabel metal3 s 0 298528 800 298648 6 dcache_tag_out[18]
port 200 nsew signal output
rlabel metal3 s 0 267248 800 267368 6 dcache_tag_out[19]
port 201 nsew signal output
rlabel metal3 s 0 382168 800 382288 6 dcache_tag_out[1]
port 202 nsew signal output
rlabel metal2 s 61198 389200 61254 390000 6 dcache_tag_out[20]
port 203 nsew signal output
rlabel metal2 s 320730 0 320786 800 6 dcache_tag_out[21]
port 204 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 dcache_tag_out[22]
port 205 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 dcache_tag_out[23]
port 206 nsew signal output
rlabel metal3 s 389200 102008 390000 102128 6 dcache_tag_out[24]
port 207 nsew signal output
rlabel metal2 s 23846 389200 23902 390000 6 dcache_tag_out[25]
port 208 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 dcache_tag_out[26]
port 209 nsew signal output
rlabel metal2 s 67638 389200 67694 390000 6 dcache_tag_out[27]
port 210 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 dcache_tag_out[28]
port 211 nsew signal output
rlabel metal2 s 235078 389200 235134 390000 6 dcache_tag_out[29]
port 212 nsew signal output
rlabel metal2 s 260838 0 260894 800 6 dcache_tag_out[2]
port 213 nsew signal output
rlabel metal3 s 389200 291048 390000 291168 6 dcache_tag_out[30]
port 214 nsew signal output
rlabel metal2 s 302698 0 302754 800 6 dcache_tag_out[31]
port 215 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 dcache_tag_out[3]
port 216 nsew signal output
rlabel metal2 s 364522 0 364578 800 6 dcache_tag_out[4]
port 217 nsew signal output
rlabel metal3 s 389200 59168 390000 59288 6 dcache_tag_out[5]
port 218 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 dcache_tag_out[6]
port 219 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 dcache_tag_out[7]
port 220 nsew signal output
rlabel metal2 s 287886 389200 287942 390000 6 dcache_tag_out[8]
port 221 nsew signal output
rlabel metal2 s 211894 389200 211950 390000 6 dcache_tag_out[9]
port 222 nsew signal output
rlabel metal3 s 389200 365848 390000 365968 6 dcache_tag_write_en
port 223 nsew signal input
rlabel metal3 s 0 310088 800 310208 6 dcache_write_data_mask_1[0]
port 224 nsew signal input
rlabel metal2 s 145562 389200 145618 390000 6 dcache_write_data_mask_1[1]
port 225 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 dcache_write_data_mask_1[2]
port 226 nsew signal input
rlabel metal3 s 389200 275408 390000 275528 6 dcache_write_data_mask_1[3]
port 227 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 dcache_write_data_mask_2[0]
port 228 nsew signal input
rlabel metal3 s 0 342728 800 342848 6 dcache_write_data_mask_2[1]
port 229 nsew signal input
rlabel metal2 s 361946 0 362002 800 6 dcache_write_data_mask_2[2]
port 230 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 dcache_write_data_mask_2[3]
port 231 nsew signal input
rlabel metal3 s 389200 307368 390000 307488 6 dcache_write_tag_mask[0]
port 232 nsew signal input
rlabel metal2 s 206742 0 206798 800 6 dcache_write_tag_mask[1]
port 233 nsew signal input
rlabel metal2 s 54758 389200 54814 390000 6 dcache_write_tag_mask[2]
port 234 nsew signal input
rlabel metal3 s 389200 214208 390000 214328 6 dcache_write_tag_mask[3]
port 235 nsew signal input
rlabel metal3 s 0 189048 800 189168 6 dram_addr0[0]
port 236 nsew signal input
rlabel metal2 s 345202 389200 345258 390000 6 dram_addr0[1]
port 237 nsew signal input
rlabel metal3 s 389200 82288 390000 82408 6 dram_addr0[2]
port 238 nsew signal input
rlabel metal2 s 282734 389200 282790 390000 6 dram_addr0[3]
port 239 nsew signal input
rlabel metal2 s 148138 389200 148194 390000 6 dram_addr0[4]
port 240 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 dram_addr0[5]
port 241 nsew signal input
rlabel metal2 s 275006 0 275062 800 6 dram_addr0[6]
port 242 nsew signal input
rlabel metal3 s 389200 237328 390000 237448 6 dram_addr0[7]
port 243 nsew signal input
rlabel metal2 s 314290 389200 314346 390000 6 dram_clk0
port 244 nsew signal input
rlabel metal3 s 0 216928 800 217048 6 dram_csb0
port 245 nsew signal input
rlabel metal2 s 300122 389200 300178 390000 6 dram_din0[0]
port 246 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 dram_din0[10]
port 247 nsew signal input
rlabel metal3 s 389200 80928 390000 81048 6 dram_din0[11]
port 248 nsew signal input
rlabel metal3 s 0 279488 800 279608 6 dram_din0[12]
port 249 nsew signal input
rlabel metal3 s 389200 376728 390000 376848 6 dram_din0[13]
port 250 nsew signal input
rlabel metal3 s 389200 163208 390000 163328 6 dram_din0[14]
port 251 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 dram_din0[15]
port 252 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 dram_din0[16]
port 253 nsew signal input
rlabel metal3 s 389200 378088 390000 378208 6 dram_din0[17]
port 254 nsew signal input
rlabel metal3 s 389200 286288 390000 286408 6 dram_din0[18]
port 255 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 dram_din0[19]
port 256 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 dram_din0[1]
port 257 nsew signal input
rlabel metal3 s 389200 192448 390000 192568 6 dram_din0[20]
port 258 nsew signal input
rlabel metal2 s 186778 389200 186834 390000 6 dram_din0[21]
port 259 nsew signal input
rlabel metal3 s 0 383528 800 383648 6 dram_din0[22]
port 260 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 dram_din0[23]
port 261 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 dram_din0[24]
port 262 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 dram_din0[25]
port 263 nsew signal input
rlabel metal3 s 0 201968 800 202088 6 dram_din0[26]
port 264 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 dram_din0[27]
port 265 nsew signal input
rlabel metal2 s 95974 389200 96030 390000 6 dram_din0[28]
port 266 nsew signal input
rlabel metal2 s 280158 0 280214 800 6 dram_din0[29]
port 267 nsew signal input
rlabel metal3 s 389200 129208 390000 129328 6 dram_din0[2]
port 268 nsew signal input
rlabel metal2 s 370962 0 371018 800 6 dram_din0[30]
port 269 nsew signal input
rlabel metal3 s 389200 21088 390000 21208 6 dram_din0[31]
port 270 nsew signal input
rlabel metal3 s 0 345448 800 345568 6 dram_din0[3]
port 271 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 dram_din0[4]
port 272 nsew signal input
rlabel metal2 s 199014 0 199070 800 6 dram_din0[5]
port 273 nsew signal input
rlabel metal3 s 0 257728 800 257848 6 dram_din0[6]
port 274 nsew signal input
rlabel metal2 s 389638 0 389694 800 6 dram_din0[7]
port 275 nsew signal input
rlabel metal2 s 333610 389200 333666 390000 6 dram_din0[8]
port 276 nsew signal input
rlabel metal3 s 389200 136008 390000 136128 6 dram_din0[9]
port 277 nsew signal input
rlabel metal2 s 191930 389200 191986 390000 6 dram_dout0[0]
port 278 nsew signal output
rlabel metal3 s 389200 99288 390000 99408 6 dram_dout0[10]
port 279 nsew signal output
rlabel metal2 s 303986 389200 304042 390000 6 dram_dout0[11]
port 280 nsew signal output
rlabel metal3 s 389200 274048 390000 274168 6 dram_dout0[12]
port 281 nsew signal output
rlabel metal3 s 0 256368 800 256488 6 dram_dout0[13]
port 282 nsew signal output
rlabel metal2 s 260838 389200 260894 390000 6 dram_dout0[14]
port 283 nsew signal output
rlabel metal3 s 0 244128 800 244248 6 dram_dout0[15]
port 284 nsew signal output
rlabel metal3 s 389200 23808 390000 23928 6 dram_dout0[16]
port 285 nsew signal output
rlabel metal3 s 0 248208 800 248328 6 dram_dout0[17]
port 286 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 dram_dout0[18]
port 287 nsew signal output
rlabel metal3 s 389200 157768 390000 157888 6 dram_dout0[19]
port 288 nsew signal output
rlabel metal3 s 389200 178168 390000 178288 6 dram_dout0[1]
port 289 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 dram_dout0[20]
port 290 nsew signal output
rlabel metal3 s 0 199928 800 200048 6 dram_dout0[21]
port 291 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 dram_dout0[22]
port 292 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 dram_dout0[23]
port 293 nsew signal output
rlabel metal2 s 282734 0 282790 800 6 dram_dout0[24]
port 294 nsew signal output
rlabel metal2 s 38014 389200 38070 390000 6 dram_dout0[25]
port 295 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 dram_dout0[26]
port 296 nsew signal output
rlabel metal3 s 389200 19728 390000 19848 6 dram_dout0[27]
port 297 nsew signal output
rlabel metal2 s 92110 389200 92166 390000 6 dram_dout0[28]
port 298 nsew signal output
rlabel metal2 s 159730 389200 159786 390000 6 dram_dout0[29]
port 299 nsew signal output
rlabel metal3 s 389200 330488 390000 330608 6 dram_dout0[2]
port 300 nsew signal output
rlabel metal2 s 52182 389200 52238 390000 6 dram_dout0[30]
port 301 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 dram_dout0[31]
port 302 nsew signal output
rlabel metal3 s 389200 241408 390000 241528 6 dram_dout0[3]
port 303 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 dram_dout0[4]
port 304 nsew signal output
rlabel metal2 s 370962 389200 371018 390000 6 dram_dout0[5]
port 305 nsew signal output
rlabel metal2 s 193218 389200 193274 390000 6 dram_dout0[6]
port 306 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 dram_dout0[7]
port 307 nsew signal output
rlabel metal3 s 389200 49648 390000 49768 6 dram_dout0[8]
port 308 nsew signal output
rlabel metal2 s 201590 0 201646 800 6 dram_dout0[9]
port 309 nsew signal output
rlabel metal3 s 389200 303288 390000 303408 6 dram_web0
port 310 nsew signal input
rlabel metal2 s 265990 389200 266046 390000 6 dram_wmask0[0]
port 311 nsew signal input
rlabel metal2 s 281446 0 281502 800 6 dram_wmask0[1]
port 312 nsew signal input
rlabel metal2 s 70214 389200 70270 390000 6 dram_wmask0[2]
port 313 nsew signal input
rlabel metal2 s 329746 0 329802 800 6 dram_wmask0[3]
port 314 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 icache_data_chip_en
port 315 nsew signal input
rlabel metal3 s 389200 253648 390000 253768 6 icache_data_in[0]
port 316 nsew signal input
rlabel metal2 s 6458 389200 6514 390000 6 icache_data_in[10]
port 317 nsew signal input
rlabel metal2 s 128818 389200 128874 390000 6 icache_data_in[11]
port 318 nsew signal input
rlabel metal2 s 185490 389200 185546 390000 6 icache_data_in[12]
port 319 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 icache_data_in[13]
port 320 nsew signal input
rlabel metal2 s 343914 0 343970 800 6 icache_data_in[14]
port 321 nsew signal input
rlabel metal2 s 213182 389200 213238 390000 6 icache_data_in[15]
port 322 nsew signal input
rlabel metal2 s 356794 0 356850 800 6 icache_data_in[16]
port 323 nsew signal input
rlabel metal3 s 0 367208 800 367328 6 icache_data_in[17]
port 324 nsew signal input
rlabel metal2 s 356794 389200 356850 390000 6 icache_data_in[18]
port 325 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 icache_data_in[19]
port 326 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 icache_data_in[1]
port 327 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 icache_data_in[20]
port 328 nsew signal input
rlabel metal2 s 226062 389200 226118 390000 6 icache_data_in[21]
port 329 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 icache_data_in[22]
port 330 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 icache_data_in[23]
port 331 nsew signal input
rlabel metal3 s 389200 64608 390000 64728 6 icache_data_in[24]
port 332 nsew signal input
rlabel metal2 s 223486 389200 223542 390000 6 icache_data_in[25]
port 333 nsew signal input
rlabel metal3 s 389200 161848 390000 161968 6 icache_data_in[26]
port 334 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 icache_data_in[27]
port 335 nsew signal input
rlabel metal3 s 389200 100648 390000 100768 6 icache_data_in[28]
port 336 nsew signal input
rlabel metal2 s 373538 389200 373594 390000 6 icache_data_in[29]
port 337 nsew signal input
rlabel metal3 s 389200 361768 390000 361888 6 icache_data_in[2]
port 338 nsew signal input
rlabel metal3 s 389200 42848 390000 42968 6 icache_data_in[30]
port 339 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 icache_data_in[31]
port 340 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 icache_data_in[3]
port 341 nsew signal input
rlabel metal3 s 0 371288 800 371408 6 icache_data_in[4]
port 342 nsew signal input
rlabel metal2 s 334898 389200 334954 390000 6 icache_data_in[5]
port 343 nsew signal input
rlabel metal3 s 389200 180888 390000 181008 6 icache_data_in[6]
port 344 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 icache_data_in[7]
port 345 nsew signal input
rlabel metal3 s 389200 184968 390000 185088 6 icache_data_in[8]
port 346 nsew signal input
rlabel metal3 s 0 235968 800 236088 6 icache_data_in[9]
port 347 nsew signal input
rlabel metal2 s 162306 389200 162362 390000 6 icache_data_index[0]
port 348 nsew signal input
rlabel metal3 s 389200 333208 390000 333328 6 icache_data_index[1]
port 349 nsew signal input
rlabel metal2 s 336186 0 336242 800 6 icache_data_index[2]
port 350 nsew signal input
rlabel metal3 s 0 295808 800 295928 6 icache_data_index[3]
port 351 nsew signal input
rlabel metal3 s 0 253648 800 253768 6 icache_data_index[4]
port 352 nsew signal input
rlabel metal2 s 385130 389200 385186 390000 6 icache_data_index[5]
port 353 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 icache_data_index[6]
port 354 nsew signal input
rlabel metal2 s 272430 0 272486 800 6 icache_data_index[7]
port 355 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 icache_data_out[0]
port 356 nsew signal output
rlabel metal3 s 389200 335928 390000 336048 6 icache_data_out[10]
port 357 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 icache_data_out[11]
port 358 nsew signal output
rlabel metal2 s 10966 389200 11022 390000 6 icache_data_out[12]
port 359 nsew signal output
rlabel metal3 s 389200 146888 390000 147008 6 icache_data_out[13]
port 360 nsew signal output
rlabel metal3 s 0 316888 800 317008 6 icache_data_out[14]
port 361 nsew signal output
rlabel metal2 s 35438 389200 35494 390000 6 icache_data_out[15]
port 362 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 icache_data_out[16]
port 363 nsew signal output
rlabel metal3 s 389200 55088 390000 55208 6 icache_data_out[17]
port 364 nsew signal output
rlabel metal3 s 0 282208 800 282328 6 icache_data_out[18]
port 365 nsew signal output
rlabel metal3 s 389200 56448 390000 56568 6 icache_data_out[19]
port 366 nsew signal output
rlabel metal2 s 85670 389200 85726 390000 6 icache_data_out[1]
port 367 nsew signal output
rlabel metal2 s 359370 389200 359426 390000 6 icache_data_out[20]
port 368 nsew signal output
rlabel metal2 s 275006 389200 275062 390000 6 icache_data_out[21]
port 369 nsew signal output
rlabel metal3 s 389200 234608 390000 234728 6 icache_data_out[22]
port 370 nsew signal output
rlabel metal3 s 389200 11568 390000 11688 6 icache_data_out[23]
port 371 nsew signal output
rlabel metal3 s 0 329128 800 329248 6 icache_data_out[24]
port 372 nsew signal output
rlabel metal3 s 0 290368 800 290488 6 icache_data_out[25]
port 373 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 icache_data_out[26]
port 374 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 icache_data_out[27]
port 375 nsew signal output
rlabel metal3 s 0 242768 800 242888 6 icache_data_out[28]
port 376 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 icache_data_out[29]
port 377 nsew signal output
rlabel metal3 s 0 222368 800 222488 6 icache_data_out[2]
port 378 nsew signal output
rlabel metal2 s 112074 389200 112130 390000 6 icache_data_out[30]
port 379 nsew signal output
rlabel metal3 s 389200 167288 390000 167408 6 icache_data_out[31]
port 380 nsew signal output
rlabel metal3 s 0 149608 800 149728 6 icache_data_out[3]
port 381 nsew signal output
rlabel metal2 s 268566 389200 268622 390000 6 icache_data_out[4]
port 382 nsew signal output
rlabel metal2 s 319442 389200 319498 390000 6 icache_data_out[5]
port 383 nsew signal output
rlabel metal2 s 247958 0 248014 800 6 icache_data_out[6]
port 384 nsew signal output
rlabel metal3 s 0 354968 800 355088 6 icache_data_out[7]
port 385 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 icache_data_out[8]
port 386 nsew signal output
rlabel metal2 s 79230 389200 79286 390000 6 icache_data_out[9]
port 387 nsew signal output
rlabel metal3 s 0 259088 800 259208 6 icache_data_write_en
port 388 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 icache_tag_chip_en
port 389 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 icache_tag_data_in[0]
port 390 nsew signal input
rlabel metal2 s 157154 389200 157210 390000 6 icache_tag_data_in[10]
port 391 nsew signal input
rlabel metal2 s 376114 0 376170 800 6 icache_tag_data_in[11]
port 392 nsew signal input
rlabel metal3 s 389200 216928 390000 217048 6 icache_tag_data_in[12]
port 393 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 icache_tag_data_in[13]
port 394 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 icache_tag_data_in[14]
port 395 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 icache_tag_data_in[15]
port 396 nsew signal input
rlabel metal3 s 389200 304648 390000 304768 6 icache_tag_data_in[16]
port 397 nsew signal input
rlabel metal3 s 389200 352248 390000 352368 6 icache_tag_data_in[17]
port 398 nsew signal input
rlabel metal3 s 389200 316888 390000 317008 6 icache_tag_data_in[18]
port 399 nsew signal input
rlabel metal3 s 0 245488 800 245608 6 icache_tag_data_in[19]
port 400 nsew signal input
rlabel metal2 s 296258 0 296314 800 6 icache_tag_data_in[1]
port 401 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 icache_tag_data_in[20]
port 402 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 icache_tag_data_in[21]
port 403 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 icache_tag_data_in[22]
port 404 nsew signal input
rlabel metal2 s 5170 389200 5226 390000 6 icache_tag_data_in[23]
port 405 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 icache_tag_data_in[24]
port 406 nsew signal input
rlabel metal3 s 389200 310088 390000 310208 6 icache_tag_data_in[25]
port 407 nsew signal input
rlabel metal2 s 198370 389200 198426 390000 6 icache_tag_data_in[26]
port 408 nsew signal input
rlabel metal2 s 300122 0 300178 800 6 icache_tag_data_in[27]
port 409 nsew signal input
rlabel metal3 s 389200 238688 390000 238808 6 icache_tag_data_in[28]
port 410 nsew signal input
rlabel metal3 s 0 319608 800 319728 6 icache_tag_data_in[29]
port 411 nsew signal input
rlabel metal3 s 0 276768 800 276888 6 icache_tag_data_in[2]
port 412 nsew signal input
rlabel metal3 s 389200 282208 390000 282328 6 icache_tag_data_in[30]
port 413 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 icache_tag_data_in[31]
port 414 nsew signal input
rlabel metal2 s 349066 389200 349122 390000 6 icache_tag_data_in[3]
port 415 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 icache_tag_data_in[4]
port 416 nsew signal input
rlabel metal3 s 389200 131928 390000 132048 6 icache_tag_data_in[5]
port 417 nsew signal input
rlabel metal3 s 389200 40128 390000 40248 6 icache_tag_data_in[6]
port 418 nsew signal input
rlabel metal2 s 368386 389200 368442 390000 6 icache_tag_data_in[7]
port 419 nsew signal input
rlabel metal3 s 389200 3408 390000 3528 6 icache_tag_data_in[8]
port 420 nsew signal input
rlabel metal3 s 0 186328 800 186448 6 icache_tag_data_in[9]
port 421 nsew signal input
rlabel metal3 s 389200 372648 390000 372768 6 icache_tag_index[0]
port 422 nsew signal input
rlabel metal3 s 389200 312808 390000 312928 6 icache_tag_index[1]
port 423 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 icache_tag_index[2]
port 424 nsew signal input
rlabel metal3 s 389200 182248 390000 182368 6 icache_tag_index[3]
port 425 nsew signal input
rlabel metal2 s 208030 389200 208086 390000 6 icache_tag_index[4]
port 426 nsew signal input
rlabel metal2 s 377402 0 377458 800 6 icache_tag_index[5]
port 427 nsew signal input
rlabel metal3 s 389200 383528 390000 383648 6 icache_tag_index[6]
port 428 nsew signal input
rlabel metal3 s 389200 212848 390000 212968 6 icache_tag_index[7]
port 429 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 icache_tag_out[0]
port 430 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 icache_tag_out[10]
port 431 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 icache_tag_out[11]
port 432 nsew signal output
rlabel metal2 s 188066 0 188122 800 6 icache_tag_out[12]
port 433 nsew signal output
rlabel metal2 s 255686 389200 255742 390000 6 icache_tag_out[13]
port 434 nsew signal output
rlabel metal2 s 101126 389200 101182 390000 6 icache_tag_out[14]
port 435 nsew signal output
rlabel metal3 s 389200 386248 390000 386368 6 icache_tag_out[15]
port 436 nsew signal output
rlabel metal3 s 389200 189728 390000 189848 6 icache_tag_out[16]
port 437 nsew signal output
rlabel metal2 s 294970 389200 295026 390000 6 icache_tag_out[17]
port 438 nsew signal output
rlabel metal2 s 388994 389200 389050 390000 6 icache_tag_out[18]
port 439 nsew signal output
rlabel metal2 s 121090 389200 121146 390000 6 icache_tag_out[19]
port 440 nsew signal output
rlabel metal3 s 0 179528 800 179648 6 icache_tag_out[1]
port 441 nsew signal output
rlabel metal3 s 389200 225088 390000 225208 6 icache_tag_out[20]
port 442 nsew signal output
rlabel metal2 s 349066 0 349122 800 6 icache_tag_out[21]
port 443 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 icache_tag_out[22]
port 444 nsew signal output
rlabel metal2 s 351642 389200 351698 390000 6 icache_tag_out[23]
port 445 nsew signal output
rlabel metal3 s 0 369928 800 370048 6 icache_tag_out[24]
port 446 nsew signal output
rlabel metal2 s 44454 389200 44510 390000 6 icache_tag_out[25]
port 447 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 icache_tag_out[26]
port 448 nsew signal output
rlabel metal3 s 0 278128 800 278248 6 icache_tag_out[27]
port 449 nsew signal output
rlabel metal2 s 346490 389200 346546 390000 6 icache_tag_out[28]
port 450 nsew signal output
rlabel metal2 s 338762 389200 338818 390000 6 icache_tag_out[29]
port 451 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 icache_tag_out[2]
port 452 nsew signal output
rlabel metal2 s 301410 389200 301466 390000 6 icache_tag_out[30]
port 453 nsew signal output
rlabel metal3 s 0 349528 800 349648 6 icache_tag_out[31]
port 454 nsew signal output
rlabel metal3 s 389200 235968 390000 236088 6 icache_tag_out[3]
port 455 nsew signal output
rlabel metal2 s 387706 389200 387762 390000 6 icache_tag_out[4]
port 456 nsew signal output
rlabel metal3 s 389200 92488 390000 92608 6 icache_tag_out[5]
port 457 nsew signal output
rlabel metal2 s 224774 0 224830 800 6 icache_tag_out[6]
port 458 nsew signal output
rlabel metal2 s 367098 0 367154 800 6 icache_tag_out[7]
port 459 nsew signal output
rlabel metal3 s 389200 172728 390000 172848 6 icache_tag_out[8]
port 460 nsew signal output
rlabel metal2 s 200302 389200 200358 390000 6 icache_tag_out[9]
port 461 nsew signal output
rlabel metal2 s 322018 0 322074 800 6 icache_tag_write_en
port 462 nsew signal input
rlabel metal3 s 389200 93848 390000 93968 6 icache_write_data_mask[0]
port 463 nsew signal input
rlabel metal2 s 307850 389200 307906 390000 6 icache_write_data_mask[1]
port 464 nsew signal input
rlabel metal3 s 0 375368 800 375488 6 icache_write_data_mask[2]
port 465 nsew signal input
rlabel metal3 s 389200 300568 390000 300688 6 icache_write_data_mask[3]
port 466 nsew signal input
rlabel metal2 s 285310 389200 285366 390000 6 icache_write_tag_mask[0]
port 467 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 icache_write_tag_mask[1]
port 468 nsew signal input
rlabel metal3 s 0 227808 800 227928 6 icache_write_tag_mask[2]
port 469 nsew signal input
rlabel metal3 s 0 286288 800 286408 6 icache_write_tag_mask[3]
port 470 nsew signal input
rlabel metal2 s 267278 389200 267334 390000 6 io_in[0]
port 471 nsew signal input
rlabel metal2 s 342626 389200 342682 390000 6 io_in[10]
port 472 nsew signal input
rlabel metal2 s 384486 0 384542 800 6 io_in[11]
port 473 nsew signal input
rlabel metal2 s 354218 0 354274 800 6 io_in[12]
port 474 nsew signal input
rlabel metal3 s 389200 142808 390000 142928 6 io_in[13]
port 475 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 io_in[14]
port 476 nsew signal input
rlabel metal3 s 389200 195168 390000 195288 6 io_in[15]
port 477 nsew signal input
rlabel metal3 s 0 323688 800 323808 6 io_in[16]
port 478 nsew signal input
rlabel metal2 s 154578 389200 154634 390000 6 io_in[17]
port 479 nsew signal input
rlabel metal3 s 0 238688 800 238808 6 io_in[18]
port 480 nsew signal input
rlabel metal3 s 0 365848 800 365968 6 io_in[19]
port 481 nsew signal input
rlabel metal2 s 158442 389200 158498 390000 6 io_in[1]
port 482 nsew signal input
rlabel metal2 s 280158 389200 280214 390000 6 io_in[20]
port 483 nsew signal input
rlabel metal3 s 389200 17008 390000 17128 6 io_in[21]
port 484 nsew signal input
rlabel metal2 s 333610 0 333666 800 6 io_in[22]
port 485 nsew signal input
rlabel metal3 s 389200 149608 390000 149728 6 io_in[23]
port 486 nsew signal input
rlabel metal2 s 311714 0 311770 800 6 io_in[24]
port 487 nsew signal input
rlabel metal2 s 313002 0 313058 800 6 io_in[25]
port 488 nsew signal input
rlabel metal3 s 389200 203328 390000 203448 6 io_in[26]
port 489 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 io_in[27]
port 490 nsew signal input
rlabel metal2 s 93398 389200 93454 390000 6 io_in[28]
port 491 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 io_in[29]
port 492 nsew signal input
rlabel metal2 s 59910 389200 59966 390000 6 io_in[2]
port 493 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 io_in[30]
port 494 nsew signal input
rlabel metal3 s 389200 179528 390000 179648 6 io_in[31]
port 495 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 io_in[32]
port 496 nsew signal input
rlabel metal2 s 202878 389200 202934 390000 6 io_in[33]
port 497 nsew signal input
rlabel metal2 s 13542 389200 13598 390000 6 io_in[34]
port 498 nsew signal input
rlabel metal2 s 28998 389200 29054 390000 6 io_in[35]
port 499 nsew signal input
rlabel metal3 s 0 269968 800 270088 6 io_in[36]
port 500 nsew signal input
rlabel metal3 s 389200 26528 390000 26648 6 io_in[37]
port 501 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 io_in[3]
port 502 nsew signal input
rlabel metal3 s 389200 308728 390000 308848 6 io_in[4]
port 503 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 io_in[5]
port 504 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 io_in[6]
port 505 nsew signal input
rlabel metal3 s 0 274048 800 274168 6 io_in[7]
port 506 nsew signal input
rlabel metal3 s 389200 140088 390000 140208 6 io_in[8]
port 507 nsew signal input
rlabel metal3 s 0 240048 800 240168 6 io_in[9]
port 508 nsew signal input
rlabel metal2 s 310426 389200 310482 390000 6 io_oeb[0]
port 509 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 io_oeb[10]
port 510 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_oeb[11]
port 511 nsew signal output
rlabel metal2 s 309138 0 309194 800 6 io_oeb[12]
port 512 nsew signal output
rlabel metal2 s 313002 389200 313058 390000 6 io_oeb[13]
port 513 nsew signal output
rlabel metal3 s 389200 75488 390000 75608 6 io_oeb[14]
port 514 nsew signal output
rlabel metal3 s 389200 268608 390000 268728 6 io_oeb[15]
port 515 nsew signal output
rlabel metal3 s 389200 183608 390000 183728 6 io_oeb[16]
port 516 nsew signal output
rlabel metal2 s 389638 389200 389694 390000 6 io_oeb[17]
port 517 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 io_oeb[18]
port 518 nsew signal output
rlabel metal3 s 0 157768 800 157888 6 io_oeb[19]
port 519 nsew signal output
rlabel metal3 s 389200 387608 390000 387728 6 io_oeb[1]
port 520 nsew signal output
rlabel metal2 s 263414 389200 263470 390000 6 io_oeb[20]
port 521 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 io_oeb[21]
port 522 nsew signal output
rlabel metal2 s 227350 0 227406 800 6 io_oeb[22]
port 523 nsew signal output
rlabel metal3 s 0 306008 800 306128 6 io_oeb[23]
port 524 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 io_oeb[24]
port 525 nsew signal output
rlabel metal3 s 389200 125128 390000 125248 6 io_oeb[25]
port 526 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 io_oeb[26]
port 527 nsew signal output
rlabel metal2 s 103702 389200 103758 390000 6 io_oeb[27]
port 528 nsew signal output
rlabel metal2 s 381910 0 381966 800 6 io_oeb[28]
port 529 nsew signal output
rlabel metal3 s 389200 327768 390000 327888 6 io_oeb[29]
port 530 nsew signal output
rlabel metal3 s 0 265888 800 266008 6 io_oeb[2]
port 531 nsew signal output
rlabel metal3 s 0 380808 800 380928 6 io_oeb[30]
port 532 nsew signal output
rlabel metal3 s 389200 112888 390000 113008 6 io_oeb[31]
port 533 nsew signal output
rlabel metal3 s 389200 27888 390000 28008 6 io_oeb[32]
port 534 nsew signal output
rlabel metal2 s 297546 0 297602 800 6 io_oeb[33]
port 535 nsew signal output
rlabel metal3 s 389200 364488 390000 364608 6 io_oeb[34]
port 536 nsew signal output
rlabel metal3 s 389200 63248 390000 63368 6 io_oeb[35]
port 537 nsew signal output
rlabel metal2 s 264702 389200 264758 390000 6 io_oeb[36]
port 538 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 io_oeb[37]
port 539 nsew signal output
rlabel metal3 s 389200 283568 390000 283688 6 io_oeb[3]
port 540 nsew signal output
rlabel metal3 s 389200 53728 390000 53848 6 io_oeb[4]
port 541 nsew signal output
rlabel metal2 s 374826 389200 374882 390000 6 io_oeb[5]
port 542 nsew signal output
rlabel metal2 s 337474 389200 337530 390000 6 io_oeb[6]
port 543 nsew signal output
rlabel metal2 s 318154 389200 318210 390000 6 io_oeb[7]
port 544 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 io_oeb[8]
port 545 nsew signal output
rlabel metal3 s 389200 114248 390000 114368 6 io_oeb[9]
port 546 nsew signal output
rlabel metal2 s 269854 389200 269910 390000 6 io_out[0]
port 547 nsew signal output
rlabel metal3 s 0 330488 800 330608 6 io_out[10]
port 548 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 io_out[11]
port 549 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 io_out[12]
port 550 nsew signal output
rlabel metal3 s 0 284928 800 285048 6 io_out[13]
port 551 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 io_out[14]
port 552 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 io_out[15]
port 553 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 io_out[16]
port 554 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 io_out[17]
port 555 nsew signal output
rlabel metal3 s 389200 357688 390000 357808 6 io_out[18]
port 556 nsew signal output
rlabel metal3 s 0 299888 800 300008 6 io_out[19]
port 557 nsew signal output
rlabel metal3 s 389200 111528 390000 111648 6 io_out[1]
port 558 nsew signal output
rlabel metal2 s 1306 389200 1362 390000 6 io_out[20]
port 559 nsew signal output
rlabel metal2 s 21270 389200 21326 390000 6 io_out[21]
port 560 nsew signal output
rlabel metal2 s 9678 389200 9734 390000 6 io_out[22]
port 561 nsew signal output
rlabel metal2 s 179050 389200 179106 390000 6 io_out[23]
port 562 nsew signal output
rlabel metal3 s 0 215568 800 215688 6 io_out[24]
port 563 nsew signal output
rlabel metal3 s 0 182248 800 182368 6 io_out[25]
port 564 nsew signal output
rlabel metal2 s 180338 0 180394 800 6 io_out[26]
port 565 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 io_out[27]
port 566 nsew signal output
rlabel metal3 s 0 261808 800 261928 6 io_out[28]
port 567 nsew signal output
rlabel metal2 s 318154 0 318210 800 6 io_out[29]
port 568 nsew signal output
rlabel metal2 s 184202 389200 184258 390000 6 io_out[2]
port 569 nsew signal output
rlabel metal3 s 0 364488 800 364608 6 io_out[30]
port 570 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 io_out[31]
port 571 nsew signal output
rlabel metal3 s 389200 200608 390000 200728 6 io_out[32]
port 572 nsew signal output
rlabel metal2 s 377402 389200 377458 390000 6 io_out[33]
port 573 nsew signal output
rlabel metal2 s 205454 389200 205510 390000 6 io_out[34]
port 574 nsew signal output
rlabel metal2 s 296258 389200 296314 390000 6 io_out[35]
port 575 nsew signal output
rlabel metal3 s 0 174088 800 174208 6 io_out[36]
port 576 nsew signal output
rlabel metal3 s 389200 342728 390000 342848 6 io_out[37]
port 577 nsew signal output
rlabel metal3 s 389200 349528 390000 349648 6 io_out[3]
port 578 nsew signal output
rlabel metal2 s 383842 389200 383898 390000 6 io_out[4]
port 579 nsew signal output
rlabel metal2 s 168746 389200 168802 390000 6 io_out[5]
port 580 nsew signal output
rlabel metal2 s 77942 389200 77998 390000 6 io_out[6]
port 581 nsew signal output
rlabel metal3 s 389200 87728 390000 87848 6 io_out[7]
port 582 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 io_out[8]
port 583 nsew signal output
rlabel metal3 s 389200 12928 390000 13048 6 io_out[9]
port 584 nsew signal output
rlabel metal2 s 306562 0 306618 800 6 iram_addr0[0]
port 585 nsew signal input
rlabel metal3 s 0 360408 800 360528 6 iram_addr0[1]
port 586 nsew signal input
rlabel metal2 s 89534 389200 89590 390000 6 iram_addr0[2]
port 587 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 iram_addr0[3]
port 588 nsew signal input
rlabel metal3 s 389200 256368 390000 256488 6 iram_addr0[4]
port 589 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 iram_addr0[5]
port 590 nsew signal input
rlabel metal2 s 345202 0 345258 800 6 iram_addr0[6]
port 591 nsew signal input
rlabel metal3 s 0 372648 800 372768 6 iram_addr0[7]
port 592 nsew signal input
rlabel metal3 s 389200 360408 390000 360528 6 iram_clk0
port 593 nsew signal input
rlabel metal2 s 19982 389200 20038 390000 6 iram_csb0_A
port 594 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 iram_csb0_B
port 595 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 iram_din0[0]
port 596 nsew signal input
rlabel metal3 s 389200 255008 390000 255128 6 iram_din0[10]
port 597 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 iram_din0[11]
port 598 nsew signal input
rlabel metal2 s 305274 389200 305330 390000 6 iram_din0[12]
port 599 nsew signal input
rlabel metal3 s 0 208768 800 208888 6 iram_din0[13]
port 600 nsew signal input
rlabel metal2 s 84382 389200 84438 390000 6 iram_din0[14]
port 601 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 iram_din0[15]
port 602 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 iram_din0[16]
port 603 nsew signal input
rlabel metal3 s 0 350888 800 351008 6 iram_din0[17]
port 604 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 iram_din0[18]
port 605 nsew signal input
rlabel metal2 s 360658 389200 360714 390000 6 iram_din0[19]
port 606 nsew signal input
rlabel metal2 s 108210 389200 108266 390000 6 iram_din0[1]
port 607 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 iram_din0[20]
port 608 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 iram_din0[21]
port 609 nsew signal input
rlabel metal2 s 354218 389200 354274 390000 6 iram_din0[22]
port 610 nsew signal input
rlabel metal3 s 0 322328 800 322448 6 iram_din0[23]
port 611 nsew signal input
rlabel metal2 s 223486 0 223542 800 6 iram_din0[24]
port 612 nsew signal input
rlabel metal3 s 0 304648 800 304768 6 iram_din0[25]
port 613 nsew signal input
rlabel metal3 s 389200 37408 390000 37528 6 iram_din0[26]
port 614 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 iram_din0[27]
port 615 nsew signal input
rlabel metal2 s 365810 0 365866 800 6 iram_din0[28]
port 616 nsew signal input
rlabel metal2 s 271142 389200 271198 390000 6 iram_din0[29]
port 617 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 iram_din0[2]
port 618 nsew signal input
rlabel metal3 s 0 163208 800 163328 6 iram_din0[30]
port 619 nsew signal input
rlabel metal3 s 389200 71408 390000 71528 6 iram_din0[31]
port 620 nsew signal input
rlabel metal3 s 0 233248 800 233368 6 iram_din0[3]
port 621 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 iram_din0[4]
port 622 nsew signal input
rlabel metal3 s 389200 74128 390000 74248 6 iram_din0[5]
port 623 nsew signal input
rlabel metal2 s 316866 389200 316922 390000 6 iram_din0[6]
port 624 nsew signal input
rlabel metal2 s 237654 389200 237710 390000 6 iram_din0[7]
port 625 nsew signal input
rlabel metal2 s 113362 389200 113418 390000 6 iram_din0[8]
port 626 nsew signal input
rlabel metal3 s 389200 337288 390000 337408 6 iram_din0[9]
port 627 nsew signal input
rlabel metal3 s 0 161848 800 161968 6 iram_dout0_A[0]
port 628 nsew signal output
rlabel metal2 s 241518 389200 241574 390000 6 iram_dout0_A[10]
port 629 nsew signal output
rlabel metal3 s 389200 264528 390000 264648 6 iram_dout0_A[11]
port 630 nsew signal output
rlabel metal2 s 319442 0 319498 800 6 iram_dout0_A[12]
port 631 nsew signal output
rlabel metal3 s 389200 186328 390000 186448 6 iram_dout0_A[13]
port 632 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 iram_dout0_A[14]
port 633 nsew signal output
rlabel metal3 s 389200 144168 390000 144288 6 iram_dout0_A[15]
port 634 nsew signal output
rlabel metal2 s 166170 389200 166226 390000 6 iram_dout0_A[16]
port 635 nsew signal output
rlabel metal2 s 124954 389200 125010 390000 6 iram_dout0_A[17]
port 636 nsew signal output
rlabel metal3 s 389200 126488 390000 126608 6 iram_dout0_A[18]
port 637 nsew signal output
rlabel metal2 s 139122 389200 139178 390000 6 iram_dout0_A[19]
port 638 nsew signal output
rlabel metal2 s 163594 389200 163650 390000 6 iram_dout0_A[1]
port 639 nsew signal output
rlabel metal3 s 389200 29248 390000 29368 6 iram_dout0_A[20]
port 640 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 iram_dout0_A[21]
port 641 nsew signal output
rlabel metal3 s 389200 379448 390000 379568 6 iram_dout0_A[22]
port 642 nsew signal output
rlabel metal3 s 389200 118328 390000 118448 6 iram_dout0_A[23]
port 643 nsew signal output
rlabel metal2 s 190642 389200 190698 390000 6 iram_dout0_A[24]
port 644 nsew signal output
rlabel metal2 s 231214 389200 231270 390000 6 iram_dout0_A[25]
port 645 nsew signal output
rlabel metal3 s 389200 293768 390000 293888 6 iram_dout0_A[26]
port 646 nsew signal output
rlabel metal3 s 0 206048 800 206168 6 iram_dout0_A[27]
port 647 nsew signal output
rlabel metal2 s 141698 389200 141754 390000 6 iram_dout0_A[28]
port 648 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 iram_dout0_A[29]
port 649 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 iram_dout0_A[2]
port 650 nsew signal output
rlabel metal3 s 389200 72768 390000 72888 6 iram_dout0_A[30]
port 651 nsew signal output
rlabel metal3 s 0 314168 800 314288 6 iram_dout0_A[31]
port 652 nsew signal output
rlabel metal3 s 389200 211488 390000 211608 6 iram_dout0_A[3]
port 653 nsew signal output
rlabel metal2 s 240230 389200 240286 390000 6 iram_dout0_A[4]
port 654 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 iram_dout0_A[5]
port 655 nsew signal output
rlabel metal3 s 389200 204688 390000 204808 6 iram_dout0_A[6]
port 656 nsew signal output
rlabel metal3 s 389200 340008 390000 340128 6 iram_dout0_A[7]
port 657 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 iram_dout0_A[8]
port 658 nsew signal output
rlabel metal2 s 27710 389200 27766 390000 6 iram_dout0_A[9]
port 659 nsew signal output
rlabel metal3 s 389200 369928 390000 370048 6 iram_dout0_B[0]
port 660 nsew signal output
rlabel metal3 s 0 190408 800 190528 6 iram_dout0_B[10]
port 661 nsew signal output
rlabel metal2 s 172610 389200 172666 390000 6 iram_dout0_B[11]
port 662 nsew signal output
rlabel metal2 s 214470 0 214526 800 6 iram_dout0_B[12]
port 663 nsew signal output
rlabel metal2 s 94686 389200 94742 390000 6 iram_dout0_B[13]
port 664 nsew signal output
rlabel metal2 s 303986 0 304042 800 6 iram_dout0_B[14]
port 665 nsew signal output
rlabel metal2 s 306562 389200 306618 390000 6 iram_dout0_B[15]
port 666 nsew signal output
rlabel metal3 s 389200 191088 390000 191208 6 iram_dout0_B[16]
port 667 nsew signal output
rlabel metal3 s 389200 141448 390000 141568 6 iram_dout0_B[17]
port 668 nsew signal output
rlabel metal2 s 177762 0 177818 800 6 iram_dout0_B[18]
port 669 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 iram_dout0_B[19]
port 670 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 iram_dout0_B[1]
port 671 nsew signal output
rlabel metal3 s 389200 104728 390000 104848 6 iram_dout0_B[20]
port 672 nsew signal output
rlabel metal2 s 350354 389200 350410 390000 6 iram_dout0_B[21]
port 673 nsew signal output
rlabel metal3 s 389200 221008 390000 221128 6 iram_dout0_B[22]
port 674 nsew signal output
rlabel metal3 s 389200 356328 390000 356448 6 iram_dout0_B[23]
port 675 nsew signal output
rlabel metal2 s 341338 389200 341394 390000 6 iram_dout0_B[24]
port 676 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 iram_dout0_B[25]
port 677 nsew signal output
rlabel metal3 s 389200 96568 390000 96688 6 iram_dout0_B[26]
port 678 nsew signal output
rlabel metal2 s 323306 0 323362 800 6 iram_dout0_B[27]
port 679 nsew signal output
rlabel metal3 s 0 326408 800 326528 6 iram_dout0_B[28]
port 680 nsew signal output
rlabel metal3 s 389200 33328 390000 33448 6 iram_dout0_B[29]
port 681 nsew signal output
rlabel metal2 s 276294 0 276350 800 6 iram_dout0_B[2]
port 682 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 iram_dout0_B[30]
port 683 nsew signal output
rlabel metal3 s 389200 374008 390000 374128 6 iram_dout0_B[31]
port 684 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 iram_dout0_B[3]
port 685 nsew signal output
rlabel metal2 s 337474 0 337530 800 6 iram_dout0_B[4]
port 686 nsew signal output
rlabel metal2 s 36726 389200 36782 390000 6 iram_dout0_B[5]
port 687 nsew signal output
rlabel metal2 s 258262 0 258318 800 6 iram_dout0_B[6]
port 688 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 iram_dout0_B[7]
port 689 nsew signal output
rlabel metal2 s 30286 389200 30342 390000 6 iram_dout0_B[8]
port 690 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 iram_dout0_B[9]
port 691 nsew signal output
rlabel metal2 s 256974 389200 257030 390000 6 iram_web0
port 692 nsew signal input
rlabel metal3 s 0 318248 800 318368 6 iram_wmask0[0]
port 693 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 iram_wmask0[1]
port 694 nsew signal input
rlabel metal3 s 389200 106088 390000 106208 6 iram_wmask0[2]
port 695 nsew signal input
rlabel metal2 s 380622 0 380678 800 6 iram_wmask0[3]
port 696 nsew signal input
rlabel metal2 s 195794 389200 195850 390000 6 la_data_in[0]
port 697 nsew signal input
rlabel metal2 s 322018 389200 322074 390000 6 la_data_in[100]
port 698 nsew signal input
rlabel metal2 s 106922 389200 106978 390000 6 la_data_in[101]
port 699 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_data_in[102]
port 700 nsew signal input
rlabel metal3 s 389200 295128 390000 295248 6 la_data_in[103]
port 701 nsew signal input
rlabel metal2 s 331034 0 331090 800 6 la_data_in[104]
port 702 nsew signal input
rlabel metal2 s 355506 389200 355562 390000 6 la_data_in[105]
port 703 nsew signal input
rlabel metal2 s 325882 389200 325938 390000 6 la_data_in[106]
port 704 nsew signal input
rlabel metal3 s 0 291728 800 291848 6 la_data_in[107]
port 705 nsew signal input
rlabel metal2 s 133970 389200 134026 390000 6 la_data_in[108]
port 706 nsew signal input
rlabel metal3 s 389200 36048 390000 36168 6 la_data_in[109]
port 707 nsew signal input
rlabel metal3 s 0 379448 800 379568 6 la_data_in[10]
port 708 nsew signal input
rlabel metal2 s 247958 389200 248014 390000 6 la_data_in[110]
port 709 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[111]
port 710 nsew signal input
rlabel metal3 s 0 271328 800 271448 6 la_data_in[112]
port 711 nsew signal input
rlabel metal3 s 389200 207408 390000 207528 6 la_data_in[113]
port 712 nsew signal input
rlabel metal2 s 45742 389200 45798 390000 6 la_data_in[114]
port 713 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 la_data_in[115]
port 714 nsew signal input
rlabel metal3 s 389200 138728 390000 138848 6 la_data_in[116]
port 715 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 la_data_in[117]
port 716 nsew signal input
rlabel metal3 s 389200 70048 390000 70168 6 la_data_in[118]
port 717 nsew signal input
rlabel metal3 s 389200 287648 390000 287768 6 la_data_in[119]
port 718 nsew signal input
rlabel metal2 s 210606 0 210662 800 6 la_data_in[11]
port 719 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[120]
port 720 nsew signal input
rlabel metal3 s 0 170008 800 170128 6 la_data_in[121]
port 721 nsew signal input
rlabel metal3 s 389200 67328 390000 67448 6 la_data_in[122]
port 722 nsew signal input
rlabel metal3 s 389200 240048 390000 240168 6 la_data_in[123]
port 723 nsew signal input
rlabel metal3 s 389200 150968 390000 151088 6 la_data_in[124]
port 724 nsew signal input
rlabel metal3 s 389200 218288 390000 218408 6 la_data_in[125]
port 725 nsew signal input
rlabel metal3 s 389200 79568 390000 79688 6 la_data_in[126]
port 726 nsew signal input
rlabel metal2 s 324594 0 324650 800 6 la_data_in[127]
port 727 nsew signal input
rlabel metal3 s 389200 368568 390000 368688 6 la_data_in[12]
port 728 nsew signal input
rlabel metal3 s 389200 14288 390000 14408 6 la_data_in[13]
port 729 nsew signal input
rlabel metal3 s 0 172728 800 172848 6 la_data_in[14]
port 730 nsew signal input
rlabel metal2 s 302698 389200 302754 390000 6 la_data_in[15]
port 731 nsew signal input
rlabel metal2 s 315578 389200 315634 390000 6 la_data_in[16]
port 732 nsew signal input
rlabel metal3 s 389200 68688 390000 68808 6 la_data_in[17]
port 733 nsew signal input
rlabel metal2 s 368386 0 368442 800 6 la_data_in[18]
port 734 nsew signal input
rlabel metal2 s 229926 389200 229982 390000 6 la_data_in[19]
port 735 nsew signal input
rlabel metal2 s 53470 389200 53526 390000 6 la_data_in[1]
port 736 nsew signal input
rlabel metal2 s 57334 389200 57390 390000 6 la_data_in[20]
port 737 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_data_in[21]
port 738 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_data_in[22]
port 739 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_data_in[23]
port 740 nsew signal input
rlabel metal3 s 389200 223728 390000 223848 6 la_data_in[24]
port 741 nsew signal input
rlabel metal2 s 347778 0 347834 800 6 la_data_in[25]
port 742 nsew signal input
rlabel metal3 s 0 226448 800 226568 6 la_data_in[26]
port 743 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[27]
port 744 nsew signal input
rlabel metal3 s 389200 133288 390000 133408 6 la_data_in[28]
port 745 nsew signal input
rlabel metal3 s 389200 159128 390000 159248 6 la_data_in[29]
port 746 nsew signal input
rlabel metal3 s 0 378088 800 378208 6 la_data_in[2]
port 747 nsew signal input
rlabel metal3 s 389200 250928 390000 251048 6 la_data_in[30]
port 748 nsew signal input
rlabel metal2 s 104990 389200 105046 390000 6 la_data_in[31]
port 749 nsew signal input
rlabel metal2 s 336186 389200 336242 390000 6 la_data_in[32]
port 750 nsew signal input
rlabel metal2 s 131394 389200 131450 390000 6 la_data_in[33]
port 751 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 la_data_in[34]
port 752 nsew signal input
rlabel metal2 s 351642 0 351698 800 6 la_data_in[35]
port 753 nsew signal input
rlabel metal2 s 16118 389200 16174 390000 6 la_data_in[36]
port 754 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 la_data_in[37]
port 755 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 la_data_in[38]
port 756 nsew signal input
rlabel metal3 s 389200 91128 390000 91248 6 la_data_in[39]
port 757 nsew signal input
rlabel metal2 s 228638 0 228694 800 6 la_data_in[3]
port 758 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_data_in[40]
port 759 nsew signal input
rlabel metal3 s 0 320968 800 321088 6 la_data_in[41]
port 760 nsew signal input
rlabel metal3 s 0 388968 800 389088 6 la_data_in[42]
port 761 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_data_in[43]
port 762 nsew signal input
rlabel metal2 s 180338 389200 180394 390000 6 la_data_in[44]
port 763 nsew signal input
rlabel metal3 s 389200 260448 390000 260568 6 la_data_in[45]
port 764 nsew signal input
rlabel metal3 s 389200 51008 390000 51128 6 la_data_in[46]
port 765 nsew signal input
rlabel metal3 s 389200 301928 390000 302048 6 la_data_in[47]
port 766 nsew signal input
rlabel metal3 s 389200 89768 390000 89888 6 la_data_in[48]
port 767 nsew signal input
rlabel metal3 s 389200 156408 390000 156528 6 la_data_in[49]
port 768 nsew signal input
rlabel metal2 s 298834 0 298890 800 6 la_data_in[4]
port 769 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_data_in[50]
port 770 nsew signal input
rlabel metal2 s 278870 0 278926 800 6 la_data_in[51]
port 771 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[52]
port 772 nsew signal input
rlabel metal2 s 188066 389200 188122 390000 6 la_data_in[53]
port 773 nsew signal input
rlabel metal3 s 389200 280848 390000 280968 6 la_data_in[54]
port 774 nsew signal input
rlabel metal2 s 218334 389200 218390 390000 6 la_data_in[55]
port 775 nsew signal input
rlabel metal3 s 0 184968 800 185088 6 la_data_in[56]
port 776 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 la_data_in[57]
port 777 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 la_data_in[58]
port 778 nsew signal input
rlabel metal3 s 389200 197888 390000 198008 6 la_data_in[59]
port 779 nsew signal input
rlabel metal3 s 389200 226448 390000 226568 6 la_data_in[5]
port 780 nsew signal input
rlabel metal3 s 389200 292408 390000 292528 6 la_data_in[60]
port 781 nsew signal input
rlabel metal2 s 137834 389200 137890 390000 6 la_data_in[61]
port 782 nsew signal input
rlabel metal2 s 364522 389200 364578 390000 6 la_data_in[62]
port 783 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[63]
port 784 nsew signal input
rlabel metal2 s 210606 389200 210662 390000 6 la_data_in[64]
port 785 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[65]
port 786 nsew signal input
rlabel metal2 s 294326 389200 294382 390000 6 la_data_in[66]
port 787 nsew signal input
rlabel metal3 s 389200 269968 390000 270088 6 la_data_in[67]
port 788 nsew signal input
rlabel metal2 s 254398 389200 254454 390000 6 la_data_in[68]
port 789 nsew signal input
rlabel metal2 s 361946 389200 362002 390000 6 la_data_in[69]
port 790 nsew signal input
rlabel metal2 s 25134 389200 25190 390000 6 la_data_in[6]
port 791 nsew signal input
rlabel metal2 s 49606 389200 49662 390000 6 la_data_in[70]
port 792 nsew signal input
rlabel metal2 s 281446 389200 281502 390000 6 la_data_in[71]
port 793 nsew signal input
rlabel metal2 s 238942 389200 238998 390000 6 la_data_in[72]
port 794 nsew signal input
rlabel metal2 s 289174 389200 289230 390000 6 la_data_in[73]
port 795 nsew signal input
rlabel metal2 s 81806 389200 81862 390000 6 la_data_in[74]
port 796 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 la_data_in[75]
port 797 nsew signal input
rlabel metal3 s 0 237328 800 237448 6 la_data_in[76]
port 798 nsew signal input
rlabel metal3 s 0 293088 800 293208 6 la_data_in[77]
port 799 nsew signal input
rlabel metal3 s 0 387608 800 387728 6 la_data_in[78]
port 800 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_data_in[79]
port 801 nsew signal input
rlabel metal3 s 389200 272688 390000 272808 6 la_data_in[7]
port 802 nsew signal input
rlabel metal2 s 244094 389200 244150 390000 6 la_data_in[80]
port 803 nsew signal input
rlabel metal2 s 115938 389200 115994 390000 6 la_data_in[81]
port 804 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 la_data_in[82]
port 805 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 la_data_in[83]
port 806 nsew signal input
rlabel metal2 s 86958 389200 87014 390000 6 la_data_in[84]
port 807 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[85]
port 808 nsew signal input
rlabel metal2 s 119802 389200 119858 390000 6 la_data_in[86]
port 809 nsew signal input
rlabel metal2 s 249246 0 249302 800 6 la_data_in[87]
port 810 nsew signal input
rlabel metal3 s 0 187688 800 187808 6 la_data_in[88]
port 811 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 la_data_in[89]
port 812 nsew signal input
rlabel metal3 s 389200 155048 390000 155168 6 la_data_in[8]
port 813 nsew signal input
rlabel metal3 s 389200 196528 390000 196648 6 la_data_in[90]
port 814 nsew signal input
rlabel metal2 s 126242 389200 126298 390000 6 la_data_in[91]
port 815 nsew signal input
rlabel metal2 s 297546 389200 297602 390000 6 la_data_in[92]
port 816 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 la_data_in[93]
port 817 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 la_data_in[94]
port 818 nsew signal input
rlabel metal2 s 238942 0 238998 800 6 la_data_in[95]
port 819 nsew signal input
rlabel metal2 s 269854 0 269910 800 6 la_data_in[96]
port 820 nsew signal input
rlabel metal3 s 389200 359048 390000 359168 6 la_data_in[97]
port 821 nsew signal input
rlabel metal2 s 227350 389200 227406 390000 6 la_data_in[98]
port 822 nsew signal input
rlabel metal3 s 389200 189048 390000 189168 6 la_data_in[99]
port 823 nsew signal input
rlabel metal2 s 176474 389200 176530 390000 6 la_data_in[9]
port 824 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 la_data_out[0]
port 825 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[100]
port 826 nsew signal output
rlabel metal3 s 0 337288 800 337408 6 la_data_out[101]
port 827 nsew signal output
rlabel metal2 s 360658 0 360714 800 6 la_data_out[102]
port 828 nsew signal output
rlabel metal3 s 389200 344088 390000 344208 6 la_data_out[103]
port 829 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 la_data_out[104]
port 830 nsew signal output
rlabel metal2 s 259550 389200 259606 390000 6 la_data_out[105]
port 831 nsew signal output
rlabel metal2 s 153290 389200 153346 390000 6 la_data_out[106]
port 832 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 la_data_out[107]
port 833 nsew signal output
rlabel metal3 s 0 218288 800 218408 6 la_data_out[108]
port 834 nsew signal output
rlabel metal3 s 0 374008 800 374128 6 la_data_out[109]
port 835 nsew signal output
rlabel metal3 s 389200 367208 390000 367328 6 la_data_out[10]
port 836 nsew signal output
rlabel metal2 s 142986 389200 143042 390000 6 la_data_out[110]
port 837 nsew signal output
rlabel metal2 s 186778 0 186834 800 6 la_data_out[111]
port 838 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[112]
port 839 nsew signal output
rlabel metal3 s 389200 318248 390000 318368 6 la_data_out[113]
port 840 nsew signal output
rlabel metal2 s 374826 0 374882 800 6 la_data_out[114]
port 841 nsew signal output
rlabel metal2 s 242806 0 242862 800 6 la_data_out[115]
port 842 nsew signal output
rlabel metal3 s 0 280848 800 280968 6 la_data_out[116]
port 843 nsew signal output
rlabel metal3 s 389200 171368 390000 171488 6 la_data_out[117]
port 844 nsew signal output
rlabel metal3 s 0 234608 800 234728 6 la_data_out[118]
port 845 nsew signal output
rlabel metal3 s 0 197208 800 197328 6 la_data_out[119]
port 846 nsew signal output
rlabel metal2 s 237654 0 237710 800 6 la_data_out[11]
port 847 nsew signal output
rlabel metal3 s 0 176808 800 176928 6 la_data_out[120]
port 848 nsew signal output
rlabel metal2 s 352930 0 352986 800 6 la_data_out[121]
port 849 nsew signal output
rlabel metal3 s 389200 265888 390000 266008 6 la_data_out[122]
port 850 nsew signal output
rlabel metal2 s 215758 389200 215814 390000 6 la_data_out[123]
port 851 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 la_data_out[124]
port 852 nsew signal output
rlabel metal3 s 389200 388968 390000 389088 6 la_data_out[125]
port 853 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 la_data_out[126]
port 854 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 la_data_out[127]
port 855 nsew signal output
rlabel metal2 s 350354 0 350410 800 6 la_data_out[12]
port 856 nsew signal output
rlabel metal2 s 164882 0 164938 800 6 la_data_out[13]
port 857 nsew signal output
rlabel metal2 s 233790 389200 233846 390000 6 la_data_out[14]
port 858 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 la_data_out[15]
port 859 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[16]
port 860 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 la_data_out[17]
port 861 nsew signal output
rlabel metal3 s 389200 210128 390000 210248 6 la_data_out[18]
port 862 nsew signal output
rlabel metal3 s 389200 52368 390000 52488 6 la_data_out[19]
port 863 nsew signal output
rlabel metal2 s 43166 389200 43222 390000 6 la_data_out[1]
port 864 nsew signal output
rlabel metal2 s 62486 389200 62542 390000 6 la_data_out[20]
port 865 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 la_data_out[21]
port 866 nsew signal output
rlabel metal3 s 389200 137368 390000 137488 6 la_data_out[22]
port 867 nsew signal output
rlabel metal3 s 389200 18368 390000 18488 6 la_data_out[23]
port 868 nsew signal output
rlabel metal2 s 258262 389200 258318 390000 6 la_data_out[24]
port 869 nsew signal output
rlabel metal2 s 340050 389200 340106 390000 6 la_data_out[25]
port 870 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 la_data_out[26]
port 871 nsew signal output
rlabel metal3 s 0 193128 800 193248 6 la_data_out[27]
port 872 nsew signal output
rlabel metal3 s 389200 22448 390000 22568 6 la_data_out[28]
port 873 nsew signal output
rlabel metal2 s 298834 389200 298890 390000 6 la_data_out[29]
port 874 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[2]
port 875 nsew signal output
rlabel metal3 s 389200 382168 390000 382288 6 la_data_out[30]
port 876 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 la_data_out[31]
port 877 nsew signal output
rlabel metal2 s 17406 389200 17462 390000 6 la_data_out[32]
port 878 nsew signal output
rlabel metal3 s 389200 242768 390000 242888 6 la_data_out[33]
port 879 nsew signal output
rlabel metal3 s 0 363128 800 363248 6 la_data_out[34]
port 880 nsew signal output
rlabel metal3 s 389200 119688 390000 119808 6 la_data_out[35]
port 881 nsew signal output
rlabel metal3 s 389200 170008 390000 170128 6 la_data_out[36]
port 882 nsew signal output
rlabel metal3 s 0 275408 800 275528 6 la_data_out[37]
port 883 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 la_data_out[38]
port 884 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 la_data_out[39]
port 885 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 la_data_out[3]
port 886 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 la_data_out[40]
port 887 nsew signal output
rlabel metal2 s 118514 389200 118570 390000 6 la_data_out[41]
port 888 nsew signal output
rlabel metal3 s 0 194488 800 194608 6 la_data_out[42]
port 889 nsew signal output
rlabel metal2 s 315578 0 315634 800 6 la_data_out[43]
port 890 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 la_data_out[44]
port 891 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[45]
port 892 nsew signal output
rlabel metal3 s 389200 83648 390000 83768 6 la_data_out[46]
port 893 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 la_data_out[47]
port 894 nsew signal output
rlabel metal2 s 31574 389200 31630 390000 6 la_data_out[48]
port 895 nsew signal output
rlabel metal3 s 389200 325048 390000 325168 6 la_data_out[49]
port 896 nsew signal output
rlabel metal2 s 305274 0 305330 800 6 la_data_out[4]
port 897 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[50]
port 898 nsew signal output
rlabel metal3 s 0 303288 800 303408 6 la_data_out[51]
port 899 nsew signal output
rlabel metal3 s 0 334568 800 334688 6 la_data_out[52]
port 900 nsew signal output
rlabel metal2 s 170034 0 170090 800 6 la_data_out[53]
port 901 nsew signal output
rlabel metal2 s 346490 0 346546 800 6 la_data_out[54]
port 902 nsew signal output
rlabel metal2 s 327170 389200 327226 390000 6 la_data_out[55]
port 903 nsew signal output
rlabel metal3 s 0 353608 800 353728 6 la_data_out[56]
port 904 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 la_data_out[57]
port 905 nsew signal output
rlabel metal2 s 291106 0 291162 800 6 la_data_out[58]
port 906 nsew signal output
rlabel metal2 s 284666 0 284722 800 6 la_data_out[59]
port 907 nsew signal output
rlabel metal2 s 32862 389200 32918 390000 6 la_data_out[5]
port 908 nsew signal output
rlabel metal2 s 293682 0 293738 800 6 la_data_out[60]
port 909 nsew signal output
rlabel metal3 s 0 272688 800 272808 6 la_data_out[61]
port 910 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 la_data_out[62]
port 911 nsew signal output
rlabel metal3 s 0 230528 800 230648 6 la_data_out[63]
port 912 nsew signal output
rlabel metal3 s 389200 85008 390000 85128 6 la_data_out[64]
port 913 nsew signal output
rlabel metal3 s 0 175448 800 175568 6 la_data_out[65]
port 914 nsew signal output
rlabel metal3 s 389200 276768 390000 276888 6 la_data_out[66]
port 915 nsew signal output
rlabel metal3 s 389200 229168 390000 229288 6 la_data_out[67]
port 916 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 la_data_out[68]
port 917 nsew signal output
rlabel metal2 s 378690 0 378746 800 6 la_data_out[69]
port 918 nsew signal output
rlabel metal2 s 196438 0 196494 800 6 la_data_out[6]
port 919 nsew signal output
rlabel metal2 s 40590 389200 40646 390000 6 la_data_out[70]
port 920 nsew signal output
rlabel metal2 s 285954 0 286010 800 6 la_data_out[71]
port 921 nsew signal output
rlabel metal3 s 389200 7488 390000 7608 6 la_data_out[72]
port 922 nsew signal output
rlabel metal2 s 316866 0 316922 800 6 la_data_out[73]
port 923 nsew signal output
rlabel metal3 s 0 264528 800 264648 6 la_data_out[74]
port 924 nsew signal output
rlabel metal2 s 331034 389200 331090 390000 6 la_data_out[75]
port 925 nsew signal output
rlabel metal2 s 262126 0 262182 800 6 la_data_out[76]
port 926 nsew signal output
rlabel metal3 s 389200 193808 390000 193928 6 la_data_out[77]
port 927 nsew signal output
rlabel metal3 s 389200 110168 390000 110288 6 la_data_out[78]
port 928 nsew signal output
rlabel metal3 s 389200 257728 390000 257848 6 la_data_out[79]
port 929 nsew signal output
rlabel metal3 s 389200 227808 390000 227928 6 la_data_out[7]
port 930 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 la_data_out[80]
port 931 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 la_data_out[81]
port 932 nsew signal output
rlabel metal3 s 0 307368 800 307488 6 la_data_out[82]
port 933 nsew signal output
rlabel metal2 s 122378 389200 122434 390000 6 la_data_out[83]
port 934 nsew signal output
rlabel metal3 s 389200 31968 390000 32088 6 la_data_out[84]
port 935 nsew signal output
rlabel metal3 s 0 325048 800 325168 6 la_data_out[85]
port 936 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 la_data_out[86]
port 937 nsew signal output
rlabel metal3 s 0 287648 800 287768 6 la_data_out[87]
port 938 nsew signal output
rlabel metal3 s 0 308728 800 308848 6 la_data_out[88]
port 939 nsew signal output
rlabel metal2 s 273718 0 273774 800 6 la_data_out[89]
port 940 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 la_data_out[8]
port 941 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 la_data_out[90]
port 942 nsew signal output
rlabel metal2 s 56046 389200 56102 390000 6 la_data_out[91]
port 943 nsew signal output
rlabel metal2 s 383198 0 383254 800 6 la_data_out[92]
port 944 nsew signal output
rlabel metal3 s 389200 41488 390000 41608 6 la_data_out[93]
port 945 nsew signal output
rlabel metal2 s 66350 389200 66406 390000 6 la_data_out[94]
port 946 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[95]
port 947 nsew signal output
rlabel metal2 s 171322 389200 171378 390000 6 la_data_out[96]
port 948 nsew signal output
rlabel metal3 s 389200 2048 390000 2168 6 la_data_out[97]
port 949 nsew signal output
rlabel metal3 s 389200 279488 390000 279608 6 la_data_out[98]
port 950 nsew signal output
rlabel metal2 s 76654 389200 76710 390000 6 la_data_out[99]
port 951 nsew signal output
rlabel metal3 s 0 301928 800 302048 6 la_data_out[9]
port 952 nsew signal output
rlabel metal3 s 389200 122408 390000 122528 6 la_oenb[0]
port 953 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 la_oenb[100]
port 954 nsew signal input
rlabel metal2 s 265990 0 266046 800 6 la_oenb[101]
port 955 nsew signal input
rlabel metal2 s 167458 389200 167514 390000 6 la_oenb[102]
port 956 nsew signal input
rlabel metal3 s 389200 176808 390000 176928 6 la_oenb[103]
port 957 nsew signal input
rlabel metal2 s 83094 389200 83150 390000 6 la_oenb[104]
port 958 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_oenb[105]
port 959 nsew signal input
rlabel metal2 s 372250 389200 372306 390000 6 la_oenb[106]
port 960 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 la_oenb[107]
port 961 nsew signal input
rlabel metal2 s 155866 389200 155922 390000 6 la_oenb[108]
port 962 nsew signal input
rlabel metal2 s 381266 389200 381322 390000 6 la_oenb[109]
port 963 nsew signal input
rlabel metal2 s 3882 389200 3938 390000 6 la_oenb[10]
port 964 nsew signal input
rlabel metal3 s 0 198568 800 198688 6 la_oenb[110]
port 965 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_oenb[111]
port 966 nsew signal input
rlabel metal3 s 0 212848 800 212968 6 la_oenb[112]
port 967 nsew signal input
rlabel metal2 s 358082 0 358138 800 6 la_oenb[113]
port 968 nsew signal input
rlabel metal3 s 389200 371288 390000 371408 6 la_oenb[114]
port 969 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[115]
port 970 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 la_oenb[116]
port 971 nsew signal input
rlabel metal2 s 284022 0 284078 800 6 la_oenb[117]
port 972 nsew signal input
rlabel metal2 s 251822 0 251878 800 6 la_oenb[118]
port 973 nsew signal input
rlabel metal3 s 0 200608 800 200728 6 la_oenb[119]
port 974 nsew signal input
rlabel metal3 s 389200 297848 390000 297968 6 la_oenb[11]
port 975 nsew signal input
rlabel metal3 s 389200 127848 390000 127968 6 la_oenb[120]
port 976 nsew signal input
rlabel metal3 s 389200 384888 390000 385008 6 la_oenb[121]
port 977 nsew signal input
rlabel metal2 s 310426 0 310482 800 6 la_oenb[122]
port 978 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_oenb[123]
port 979 nsew signal input
rlabel metal2 s 12254 389200 12310 390000 6 la_oenb[124]
port 980 nsew signal input
rlabel metal2 s 277582 389200 277638 390000 6 la_oenb[125]
port 981 nsew signal input
rlabel metal3 s 389200 261808 390000 261928 6 la_oenb[126]
port 982 nsew signal input
rlabel metal3 s 389200 334568 390000 334688 6 la_oenb[127]
port 983 nsew signal input
rlabel metal3 s 389200 4768 390000 4888 6 la_oenb[12]
port 984 nsew signal input
rlabel metal3 s 389200 219648 390000 219768 6 la_oenb[13]
port 985 nsew signal input
rlabel metal3 s 0 207408 800 207528 6 la_oenb[14]
port 986 nsew signal input
rlabel metal2 s 18694 389200 18750 390000 6 la_oenb[15]
port 987 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_oenb[16]
port 988 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_oenb[17]
port 989 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[18]
port 990 nsew signal input
rlabel metal3 s 389200 175448 390000 175568 6 la_oenb[19]
port 991 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_oenb[1]
port 992 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[20]
port 993 nsew signal input
rlabel metal3 s 389200 160488 390000 160608 6 la_oenb[21]
port 994 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_oenb[22]
port 995 nsew signal input
rlabel metal3 s 389200 289688 390000 289808 6 la_oenb[23]
port 996 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[24]
port 997 nsew signal input
rlabel metal3 s 389200 252288 390000 252408 6 la_oenb[25]
port 998 nsew signal input
rlabel metal2 s 325882 0 325938 800 6 la_oenb[26]
port 999 nsew signal input
rlabel metal2 s 164882 389200 164938 390000 6 la_oenb[27]
port 1000 nsew signal input
rlabel metal2 s 301410 0 301466 800 6 la_oenb[28]
port 1001 nsew signal input
rlabel metal3 s 389200 346808 390000 346928 6 la_oenb[29]
port 1002 nsew signal input
rlabel metal2 s 224774 389200 224830 390000 6 la_oenb[2]
port 1003 nsew signal input
rlabel metal2 s 173898 389200 173954 390000 6 la_oenb[30]
port 1004 nsew signal input
rlabel metal2 s 58622 389200 58678 390000 6 la_oenb[31]
port 1005 nsew signal input
rlabel metal2 s 232502 389200 232558 390000 6 la_oenb[32]
port 1006 nsew signal input
rlabel metal3 s 0 283568 800 283688 6 la_oenb[33]
port 1007 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oenb[34]
port 1008 nsew signal input
rlabel metal3 s 389200 108808 390000 108928 6 la_oenb[35]
port 1009 nsew signal input
rlabel metal3 s 389200 230528 390000 230648 6 la_oenb[36]
port 1010 nsew signal input
rlabel metal3 s 389200 353608 390000 353728 6 la_oenb[37]
port 1011 nsew signal input
rlabel metal2 s 2594 389200 2650 390000 6 la_oenb[38]
port 1012 nsew signal input
rlabel metal2 s 355506 0 355562 800 6 la_oenb[39]
port 1013 nsew signal input
rlabel metal2 s 323306 389200 323362 390000 6 la_oenb[3]
port 1014 nsew signal input
rlabel metal2 s 382554 389200 382610 390000 6 la_oenb[40]
port 1015 nsew signal input
rlabel metal2 s 201590 389200 201646 390000 6 la_oenb[41]
port 1016 nsew signal input
rlabel metal2 s 284022 389200 284078 390000 6 la_oenb[42]
port 1017 nsew signal input
rlabel metal3 s 389200 34688 390000 34808 6 la_oenb[43]
port 1018 nsew signal input
rlabel metal2 s 278870 389200 278926 390000 6 la_oenb[44]
port 1019 nsew signal input
rlabel metal3 s 389200 15648 390000 15768 6 la_oenb[45]
port 1020 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 la_oenb[46]
port 1021 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[47]
port 1022 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_oenb[48]
port 1023 nsew signal input
rlabel metal3 s 389200 44208 390000 44328 6 la_oenb[49]
port 1024 nsew signal input
rlabel metal3 s 389200 208768 390000 208888 6 la_oenb[4]
port 1025 nsew signal input
rlabel metal2 s 332322 389200 332378 390000 6 la_oenb[50]
port 1026 nsew signal input
rlabel metal2 s 34150 389200 34206 390000 6 la_oenb[51]
port 1027 nsew signal input
rlabel metal2 s 14830 389200 14886 390000 6 la_oenb[52]
port 1028 nsew signal input
rlabel metal3 s 0 333208 800 333328 6 la_oenb[53]
port 1029 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_oenb[54]
port 1030 nsew signal input
rlabel metal2 s 291750 389200 291806 390000 6 la_oenb[55]
port 1031 nsew signal input
rlabel metal3 s 389200 86368 390000 86488 6 la_oenb[56]
port 1032 nsew signal input
rlabel metal3 s 0 312808 800 312928 6 la_oenb[57]
port 1033 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[58]
port 1034 nsew signal input
rlabel metal2 s 347778 389200 347834 390000 6 la_oenb[59]
port 1035 nsew signal input
rlabel metal2 s 127530 389200 127586 390000 6 la_oenb[5]
port 1036 nsew signal input
rlabel metal2 s 102414 389200 102470 390000 6 la_oenb[60]
port 1037 nsew signal input
rlabel metal2 s 182914 389200 182970 390000 6 la_oenb[61]
port 1038 nsew signal input
rlabel metal2 s 204166 389200 204222 390000 6 la_oenb[62]
port 1039 nsew signal input
rlabel metal2 s 209318 389200 209374 390000 6 la_oenb[63]
port 1040 nsew signal input
rlabel metal2 s 263414 0 263470 800 6 la_oenb[64]
port 1041 nsew signal input
rlabel metal2 s 63774 389200 63830 390000 6 la_oenb[65]
port 1042 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 la_oenb[66]
port 1043 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 la_oenb[67]
port 1044 nsew signal input
rlabel metal3 s 389200 688 390000 808 6 la_oenb[68]
port 1045 nsew signal input
rlabel metal2 s 264702 0 264758 800 6 la_oenb[69]
port 1046 nsew signal input
rlabel metal3 s 389200 145528 390000 145648 6 la_oenb[6]
port 1047 nsew signal input
rlabel metal2 s 114650 389200 114706 390000 6 la_oenb[70]
port 1048 nsew signal input
rlabel metal3 s 0 688 800 808 6 la_oenb[71]
port 1049 nsew signal input
rlabel metal3 s 0 204688 800 204808 6 la_oenb[72]
port 1050 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_oenb[73]
port 1051 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[74]
port 1052 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_oenb[75]
port 1053 nsew signal input
rlabel metal2 s 68926 389200 68982 390000 6 la_oenb[76]
port 1054 nsew signal input
rlabel metal3 s 389200 8848 390000 8968 6 la_oenb[77]
port 1055 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_oenb[78]
port 1056 nsew signal input
rlabel metal2 s 372250 0 372306 800 6 la_oenb[79]
port 1057 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 la_oenb[7]
port 1058 nsew signal input
rlabel metal2 s 328458 389200 328514 390000 6 la_oenb[80]
port 1059 nsew signal input
rlabel metal2 s 379978 0 380034 800 6 la_oenb[81]
port 1060 nsew signal input
rlabel metal3 s 0 221008 800 221128 6 la_oenb[82]
port 1061 nsew signal input
rlabel metal3 s 389200 97928 390000 98048 6 la_oenb[83]
port 1062 nsew signal input
rlabel metal2 s 352930 389200 352986 390000 6 la_oenb[84]
port 1063 nsew signal input
rlabel metal2 s 22558 389200 22614 390000 6 la_oenb[85]
port 1064 nsew signal input
rlabel metal3 s 389200 363128 390000 363248 6 la_oenb[86]
port 1065 nsew signal input
rlabel metal2 s 369674 0 369730 800 6 la_oenb[87]
port 1066 nsew signal input
rlabel metal2 s 130106 389200 130162 390000 6 la_oenb[88]
port 1067 nsew signal input
rlabel metal3 s 389200 148248 390000 148368 6 la_oenb[89]
port 1068 nsew signal input
rlabel metal3 s 0 386248 800 386368 6 la_oenb[8]
port 1069 nsew signal input
rlabel metal3 s 389200 57808 390000 57928 6 la_oenb[90]
port 1070 nsew signal input
rlabel metal3 s 0 214208 800 214328 6 la_oenb[91]
port 1071 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[92]
port 1072 nsew signal input
rlabel metal3 s 389200 341368 390000 341488 6 la_oenb[93]
port 1073 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 la_oenb[94]
port 1074 nsew signal input
rlabel metal2 s 365810 389200 365866 390000 6 la_oenb[95]
port 1075 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oenb[96]
port 1076 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 la_oenb[97]
port 1077 nsew signal input
rlabel metal3 s 0 263168 800 263288 6 la_oenb[98]
port 1078 nsew signal input
rlabel metal2 s 146850 389200 146906 390000 6 la_oenb[99]
port 1079 nsew signal input
rlabel metal2 s 324594 389200 324650 390000 6 la_oenb[9]
port 1080 nsew signal input
rlabel metal3 s 0 252288 800 252408 6 user_irq[0]
port 1081 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 user_irq[1]
port 1082 nsew signal output
rlabel metal3 s 389200 164568 390000 164688 6 user_irq[2]
port 1083 nsew signal output
rlabel metal4 s 4208 2128 4528 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 387376 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 387376 6 vssd1
port 1085 nsew ground bidirectional
rlabel metal3 s 0 229168 800 229288 6 wb_rst_i
port 1086 nsew signal input
rlabel metal3 s 389200 245488 390000 245608 6 wbs_ack_o
port 1087 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 wbs_adr_i[0]
port 1088 nsew signal input
rlabel metal3 s 0 368568 800 368688 6 wbs_adr_i[10]
port 1089 nsew signal input
rlabel metal3 s 0 180888 800 181008 6 wbs_adr_i[11]
port 1090 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_adr_i[12]
port 1091 nsew signal input
rlabel metal2 s 256974 0 257030 800 6 wbs_adr_i[13]
port 1092 nsew signal input
rlabel metal2 s 358082 389200 358138 390000 6 wbs_adr_i[14]
port 1093 nsew signal input
rlabel metal2 s 386418 389200 386474 390000 6 wbs_adr_i[15]
port 1094 nsew signal input
rlabel metal2 s 289818 0 289874 800 6 wbs_adr_i[16]
port 1095 nsew signal input
rlabel metal3 s 389200 354968 390000 355088 6 wbs_adr_i[17]
port 1096 nsew signal input
rlabel metal3 s 389200 215568 390000 215688 6 wbs_adr_i[18]
port 1097 nsew signal input
rlabel metal3 s 389200 48288 390000 48408 6 wbs_adr_i[19]
port 1098 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wbs_adr_i[1]
port 1099 nsew signal input
rlabel metal2 s 219622 389200 219678 390000 6 wbs_adr_i[20]
port 1100 nsew signal input
rlabel metal2 s 255686 0 255742 800 6 wbs_adr_i[21]
port 1101 nsew signal input
rlabel metal2 s 363234 0 363290 800 6 wbs_adr_i[22]
port 1102 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 wbs_adr_i[23]
port 1103 nsew signal input
rlabel metal3 s 0 250928 800 251048 6 wbs_adr_i[24]
port 1104 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 wbs_adr_i[25]
port 1105 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_adr_i[26]
port 1106 nsew signal input
rlabel metal3 s 0 361768 800 361888 6 wbs_adr_i[27]
port 1107 nsew signal input
rlabel metal3 s 389200 326408 390000 326528 6 wbs_adr_i[28]
port 1108 nsew signal input
rlabel metal2 s 286598 389200 286654 390000 6 wbs_adr_i[29]
port 1109 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 wbs_adr_i[2]
port 1110 nsew signal input
rlabel metal2 s 181626 389200 181682 390000 6 wbs_adr_i[30]
port 1111 nsew signal input
rlabel metal3 s 389200 246848 390000 246968 6 wbs_adr_i[31]
port 1112 nsew signal input
rlabel metal2 s 341338 0 341394 800 6 wbs_adr_i[3]
port 1113 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wbs_adr_i[4]
port 1114 nsew signal input
rlabel metal2 s 327170 0 327226 800 6 wbs_adr_i[5]
port 1115 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 wbs_adr_i[6]
port 1116 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[7]
port 1117 nsew signal input
rlabel metal3 s 389200 45568 390000 45688 6 wbs_adr_i[8]
port 1118 nsew signal input
rlabel metal3 s 389200 168648 390000 168768 6 wbs_adr_i[9]
port 1119 nsew signal input
rlabel metal3 s 0 384888 800 385008 6 wbs_cyc_i
port 1120 nsew signal input
rlabel metal2 s 343914 389200 343970 390000 6 wbs_dat_i[0]
port 1121 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 wbs_dat_i[10]
port 1122 nsew signal input
rlabel metal3 s 0 178168 800 178288 6 wbs_dat_i[11]
port 1123 nsew signal input
rlabel metal3 s 0 167288 800 167408 6 wbs_dat_i[12]
port 1124 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[13]
port 1125 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 wbs_dat_i[14]
port 1126 nsew signal input
rlabel metal3 s 389200 271328 390000 271448 6 wbs_dat_i[15]
port 1127 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 wbs_dat_i[16]
port 1128 nsew signal input
rlabel metal2 s 170034 389200 170090 390000 6 wbs_dat_i[17]
port 1129 nsew signal input
rlabel metal2 s 273718 389200 273774 390000 6 wbs_dat_i[18]
port 1130 nsew signal input
rlabel metal3 s 0 294448 800 294568 6 wbs_dat_i[19]
port 1131 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 wbs_dat_i[1]
port 1132 nsew signal input
rlabel metal3 s 389200 299208 390000 299328 6 wbs_dat_i[20]
port 1133 nsew signal input
rlabel metal2 s 293038 389200 293094 390000 6 wbs_dat_i[21]
port 1134 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 wbs_dat_i[22]
port 1135 nsew signal input
rlabel metal3 s 389200 375368 390000 375488 6 wbs_dat_i[23]
port 1136 nsew signal input
rlabel metal3 s 389200 174088 390000 174208 6 wbs_dat_i[24]
port 1137 nsew signal input
rlabel metal2 s 288530 0 288586 800 6 wbs_dat_i[25]
port 1138 nsew signal input
rlabel metal2 s 250534 389200 250590 390000 6 wbs_dat_i[26]
port 1139 nsew signal input
rlabel metal2 s 7746 389200 7802 390000 6 wbs_dat_i[27]
port 1140 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 wbs_dat_i[28]
port 1141 nsew signal input
rlabel metal3 s 389200 289008 390000 289128 6 wbs_dat_i[29]
port 1142 nsew signal input
rlabel metal2 s 338762 0 338818 800 6 wbs_dat_i[2]
port 1143 nsew signal input
rlabel metal3 s 389200 152328 390000 152448 6 wbs_dat_i[30]
port 1144 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 wbs_dat_i[31]
port 1145 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 wbs_dat_i[3]
port 1146 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_i[4]
port 1147 nsew signal input
rlabel metal2 s 202878 0 202934 800 6 wbs_dat_i[5]
port 1148 nsew signal input
rlabel metal3 s 389200 206048 390000 206168 6 wbs_dat_i[6]
port 1149 nsew signal input
rlabel metal2 s 251822 389200 251878 390000 6 wbs_dat_i[7]
port 1150 nsew signal input
rlabel metal2 s 379978 389200 380034 390000 6 wbs_dat_i[8]
port 1151 nsew signal input
rlabel metal3 s 389200 38768 390000 38888 6 wbs_dat_i[9]
port 1152 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[0]
port 1153 nsew signal output
rlabel metal3 s 389200 259088 390000 259208 6 wbs_dat_o[10]
port 1154 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[11]
port 1155 nsew signal output
rlabel metal2 s 376114 389200 376170 390000 6 wbs_dat_o[12]
port 1156 nsew signal output
rlabel metal2 s 246670 389200 246726 390000 6 wbs_dat_o[13]
port 1157 nsew signal output
rlabel metal3 s 389200 61888 390000 62008 6 wbs_dat_o[14]
port 1158 nsew signal output
rlabel metal2 s 236366 389200 236422 390000 6 wbs_dat_o[15]
port 1159 nsew signal output
rlabel metal2 s 271142 0 271198 800 6 wbs_dat_o[16]
port 1160 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 wbs_dat_o[17]
port 1161 nsew signal output
rlabel metal2 s 268566 0 268622 800 6 wbs_dat_o[18]
port 1162 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 1163 nsew signal output
rlabel metal2 s 314290 0 314346 800 6 wbs_dat_o[1]
port 1164 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 wbs_dat_o[20]
port 1165 nsew signal output
rlabel metal3 s 0 297168 800 297288 6 wbs_dat_o[21]
port 1166 nsew signal output
rlabel metal2 s 74078 389200 74134 390000 6 wbs_dat_o[22]
port 1167 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 wbs_dat_o[23]
port 1168 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 wbs_dat_o[24]
port 1169 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[25]
port 1170 nsew signal output
rlabel metal2 s 177762 389200 177818 390000 6 wbs_dat_o[26]
port 1171 nsew signal output
rlabel metal2 s 90822 389200 90878 390000 6 wbs_dat_o[27]
port 1172 nsew signal output
rlabel metal2 s 213182 0 213238 800 6 wbs_dat_o[28]
port 1173 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 wbs_dat_o[29]
port 1174 nsew signal output
rlabel metal3 s 389200 115608 390000 115728 6 wbs_dat_o[2]
port 1175 nsew signal output
rlabel metal3 s 0 231888 800 232008 6 wbs_dat_o[30]
port 1176 nsew signal output
rlabel metal3 s 389200 315528 390000 315648 6 wbs_dat_o[31]
port 1177 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 wbs_dat_o[3]
port 1178 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 wbs_dat_o[4]
port 1179 nsew signal output
rlabel metal2 s 233790 0 233846 800 6 wbs_dat_o[5]
port 1180 nsew signal output
rlabel metal3 s 389200 296488 390000 296608 6 wbs_dat_o[6]
port 1181 nsew signal output
rlabel metal2 s 235078 0 235134 800 6 wbs_dat_o[7]
port 1182 nsew signal output
rlabel metal2 s 249246 389200 249302 390000 6 wbs_dat_o[8]
port 1183 nsew signal output
rlabel metal2 s 245382 389200 245438 390000 6 wbs_dat_o[9]
port 1184 nsew signal output
rlabel metal3 s 0 359048 800 359168 6 wbs_sel_i[0]
port 1185 nsew signal input
rlabel metal2 s 41878 389200 41934 390000 6 wbs_sel_i[1]
port 1186 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 wbs_sel_i[2]
port 1187 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 wbs_sel_i[3]
port 1188 nsew signal input
rlabel metal3 s 0 327768 800 327888 6 wbs_stb_i
port 1189 nsew signal input
rlabel metal3 s 389200 187688 390000 187808 6 wbs_we_i
port 1190 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 390000 390000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 186833032
string GDS_FILE /work/stu/yzhu/ai-chip/rioschip/openlane/top/runs/22_10_31_22_03/results/signoff/top.magic.gds
string GDS_START 1586186
<< end >>

