magic
tech sky130B
magscale 1 2
timestamp 1662987572
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 1104 2128 28888 27792
<< metal2 >>
rect 18 29200 74 30000
rect 1306 29200 1362 30000
rect 1950 29200 2006 30000
rect 2594 29200 2650 30000
rect 3882 29200 3938 30000
rect 4526 29200 4582 30000
rect 5814 29200 5870 30000
rect 6458 29200 6514 30000
rect 7746 29200 7802 30000
rect 8390 29200 8446 30000
rect 9034 29200 9090 30000
rect 10322 29200 10378 30000
rect 10966 29200 11022 30000
rect 12254 29200 12310 30000
rect 12898 29200 12954 30000
rect 13542 29200 13598 30000
rect 14830 29200 14886 30000
rect 15474 29200 15530 30000
rect 16118 29200 16174 30000
rect 17406 29200 17462 30000
rect 18050 29200 18106 30000
rect 19338 29200 19394 30000
rect 19982 29200 20038 30000
rect 20626 29200 20682 30000
rect 21914 29200 21970 30000
rect 22558 29200 22614 30000
rect 23846 29200 23902 30000
rect 24490 29200 24546 30000
rect 25134 29200 25190 30000
rect 26422 29200 26478 30000
rect 27066 29200 27122 30000
rect 28354 29200 28410 30000
rect 28998 29200 29054 30000
rect 29642 29200 29698 30000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 29642 0 29698 800
<< obsm2 >>
rect 4424 856 28226 27781
rect 4424 800 4470 856
rect 4638 800 5114 856
rect 5282 800 5758 856
rect 5926 800 7046 856
rect 7214 800 7690 856
rect 7858 800 8978 856
rect 9146 800 9622 856
rect 9790 800 10266 856
rect 10434 800 11554 856
rect 11722 800 12198 856
rect 12366 800 13486 856
rect 13654 800 14130 856
rect 14298 800 14774 856
rect 14942 800 16062 856
rect 16230 800 16706 856
rect 16874 800 17994 856
rect 18162 800 18638 856
rect 18806 800 19282 856
rect 19450 800 20570 856
rect 20738 800 21214 856
rect 21382 800 22502 856
rect 22670 800 23146 856
rect 23314 800 23790 856
rect 23958 800 25078 856
rect 25246 800 25722 856
rect 25890 800 27010 856
rect 27178 800 27654 856
rect 27822 800 28226 856
<< metal3 >>
rect 0 29248 800 29368
rect 29200 28568 30000 28688
rect 0 27888 800 28008
rect 29200 27888 30000 28008
rect 0 27208 800 27328
rect 0 26528 800 26648
rect 29200 26528 30000 26648
rect 29200 25848 30000 25968
rect 0 25168 800 25288
rect 29200 25168 30000 25288
rect 0 24488 800 24608
rect 29200 23808 30000 23928
rect 0 23128 800 23248
rect 29200 23128 30000 23248
rect 0 22448 800 22568
rect 0 21768 800 21888
rect 29200 21768 30000 21888
rect 29200 21088 30000 21208
rect 0 20408 800 20528
rect 29200 20408 30000 20528
rect 0 19728 800 19848
rect 29200 19048 30000 19168
rect 0 18368 800 18488
rect 29200 18368 30000 18488
rect 0 17688 800 17808
rect 0 17008 800 17128
rect 29200 17008 30000 17128
rect 29200 16328 30000 16448
rect 0 15648 800 15768
rect 29200 15648 30000 15768
rect 0 14968 800 15088
rect 29200 14288 30000 14408
rect 0 13608 800 13728
rect 29200 13608 30000 13728
rect 0 12928 800 13048
rect 0 12248 800 12368
rect 29200 12248 30000 12368
rect 29200 11568 30000 11688
rect 0 10888 800 11008
rect 0 10208 800 10328
rect 29200 10208 30000 10328
rect 29200 9528 30000 9648
rect 0 8848 800 8968
rect 29200 8848 30000 8968
rect 0 8168 800 8288
rect 0 7488 800 7608
rect 29200 7488 30000 7608
rect 29200 6808 30000 6928
rect 0 6128 800 6248
rect 29200 6128 30000 6248
rect 0 5448 800 5568
rect 29200 4768 30000 4888
rect 0 4088 800 4208
rect 29200 4088 30000 4208
rect 0 3408 800 3528
rect 0 2728 800 2848
rect 29200 2728 30000 2848
rect 29200 2048 30000 2168
rect 0 1368 800 1488
rect 29200 1368 30000 1488
rect 0 688 800 808
rect 29200 8 30000 128
<< obsm3 >>
rect 4420 26728 29200 27777
rect 4420 26448 29120 26728
rect 4420 26048 29200 26448
rect 4420 25768 29120 26048
rect 4420 25368 29200 25768
rect 4420 25088 29120 25368
rect 4420 24008 29200 25088
rect 4420 23728 29120 24008
rect 4420 23328 29200 23728
rect 4420 23048 29120 23328
rect 4420 21968 29200 23048
rect 4420 21688 29120 21968
rect 4420 21288 29200 21688
rect 4420 21008 29120 21288
rect 4420 20608 29200 21008
rect 4420 20328 29120 20608
rect 4420 19248 29200 20328
rect 4420 18968 29120 19248
rect 4420 18568 29200 18968
rect 4420 18288 29120 18568
rect 4420 17208 29200 18288
rect 4420 16928 29120 17208
rect 4420 16528 29200 16928
rect 4420 16248 29120 16528
rect 4420 15848 29200 16248
rect 4420 15568 29120 15848
rect 4420 14488 29200 15568
rect 4420 14208 29120 14488
rect 4420 13808 29200 14208
rect 4420 13528 29120 13808
rect 4420 12448 29200 13528
rect 4420 12168 29120 12448
rect 4420 11768 29200 12168
rect 4420 11488 29120 11768
rect 4420 10408 29200 11488
rect 4420 10128 29120 10408
rect 4420 9728 29200 10128
rect 4420 9448 29120 9728
rect 4420 9048 29200 9448
rect 4420 8768 29120 9048
rect 4420 7688 29200 8768
rect 4420 7408 29120 7688
rect 4420 7008 29200 7408
rect 4420 6728 29120 7008
rect 4420 6328 29200 6728
rect 4420 6048 29120 6328
rect 4420 4968 29200 6048
rect 4420 4688 29120 4968
rect 4420 4288 29200 4688
rect 4420 4008 29120 4288
rect 4420 2928 29200 4008
rect 4420 2648 29120 2928
rect 4420 2248 29200 2648
rect 4420 2143 29120 2248
<< metal4 >>
rect 4418 2128 4738 27792
rect 7892 2128 8212 27792
rect 11366 2128 11686 27792
rect 14840 2128 15160 27792
rect 18314 2128 18634 27792
rect 21788 2128 22108 27792
rect 25262 2128 25582 27792
<< labels >>
rlabel metal2 s 7102 0 7158 800 6 hehe_rstn
port 1 nsew signal output
rlabel metal3 s 29200 16328 30000 16448 6 la_data_in[0]
port 2 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[100]
port 3 nsew signal input
rlabel metal3 s 29200 21768 30000 21888 6 la_data_in[101]
port 4 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_data_in[102]
port 5 nsew signal input
rlabel metal2 s 29642 29200 29698 30000 6 la_data_in[103]
port 6 nsew signal input
rlabel metal3 s 29200 6808 30000 6928 6 la_data_in[104]
port 7 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 la_data_in[105]
port 8 nsew signal input
rlabel metal2 s 12898 29200 12954 30000 6 la_data_in[106]
port 9 nsew signal input
rlabel metal2 s 15474 29200 15530 30000 6 la_data_in[107]
port 10 nsew signal input
rlabel metal2 s 26422 29200 26478 30000 6 la_data_in[108]
port 11 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 la_data_in[109]
port 12 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_data_in[10]
port 13 nsew signal input
rlabel metal2 s 28998 29200 29054 30000 6 la_data_in[110]
port 14 nsew signal input
rlabel metal2 s 2594 29200 2650 30000 6 la_data_in[111]
port 15 nsew signal input
rlabel metal2 s 24490 29200 24546 30000 6 la_data_in[112]
port 16 nsew signal input
rlabel metal2 s 12254 29200 12310 30000 6 la_data_in[113]
port 17 nsew signal input
rlabel metal3 s 29200 10208 30000 10328 6 la_data_in[114]
port 18 nsew signal input
rlabel metal3 s 29200 14288 30000 14408 6 la_data_in[115]
port 19 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[116]
port 20 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la_data_in[117]
port 21 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 la_data_in[118]
port 22 nsew signal input
rlabel metal2 s 7746 29200 7802 30000 6 la_data_in[119]
port 23 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_data_in[11]
port 24 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 la_data_in[120]
port 25 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_data_in[121]
port 26 nsew signal input
rlabel metal3 s 29200 17008 30000 17128 6 la_data_in[122]
port 27 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_data_in[123]
port 28 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_data_in[124]
port 29 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 la_data_in[125]
port 30 nsew signal input
rlabel metal3 s 29200 21088 30000 21208 6 la_data_in[126]
port 31 nsew signal input
rlabel metal2 s 8390 29200 8446 30000 6 la_data_in[127]
port 32 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_data_in[12]
port 33 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 la_data_in[13]
port 34 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 la_data_in[14]
port 35 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 la_data_in[15]
port 36 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 la_data_in[16]
port 37 nsew signal input
rlabel metal2 s 28354 29200 28410 30000 6 la_data_in[17]
port 38 nsew signal input
rlabel metal2 s 25134 29200 25190 30000 6 la_data_in[18]
port 39 nsew signal input
rlabel metal2 s 6458 29200 6514 30000 6 la_data_in[19]
port 40 nsew signal input
rlabel metal3 s 29200 9528 30000 9648 6 la_data_in[1]
port 41 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 la_data_in[20]
port 42 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 la_data_in[21]
port 43 nsew signal input
rlabel metal2 s 4526 29200 4582 30000 6 la_data_in[22]
port 44 nsew signal input
rlabel metal2 s 16118 29200 16174 30000 6 la_data_in[23]
port 45 nsew signal input
rlabel metal2 s 662 0 718 800 6 la_data_in[24]
port 46 nsew signal input
rlabel metal2 s 20626 29200 20682 30000 6 la_data_in[25]
port 47 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 la_data_in[26]
port 48 nsew signal input
rlabel metal2 s 19982 29200 20038 30000 6 la_data_in[27]
port 49 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_data_in[28]
port 50 nsew signal input
rlabel metal3 s 29200 27888 30000 28008 6 la_data_in[29]
port 51 nsew signal input
rlabel metal3 s 29200 23128 30000 23248 6 la_data_in[2]
port 52 nsew signal input
rlabel metal3 s 29200 19048 30000 19168 6 la_data_in[30]
port 53 nsew signal input
rlabel metal3 s 29200 2048 30000 2168 6 la_data_in[31]
port 54 nsew signal input
rlabel metal2 s 10322 29200 10378 30000 6 la_data_in[32]
port 55 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 la_data_in[33]
port 56 nsew signal input
rlabel metal3 s 29200 28568 30000 28688 6 la_data_in[34]
port 57 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 la_data_in[35]
port 58 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 la_data_in[36]
port 59 nsew signal input
rlabel metal2 s 18050 29200 18106 30000 6 la_data_in[37]
port 60 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 la_data_in[38]
port 61 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 la_data_in[39]
port 62 nsew signal input
rlabel metal2 s 1950 29200 2006 30000 6 la_data_in[3]
port 63 nsew signal input
rlabel metal3 s 29200 25168 30000 25288 6 la_data_in[40]
port 64 nsew signal input
rlabel metal2 s 3882 29200 3938 30000 6 la_data_in[41]
port 65 nsew signal input
rlabel metal2 s 10966 29200 11022 30000 6 la_data_in[42]
port 66 nsew signal input
rlabel metal2 s 13542 29200 13598 30000 6 la_data_in[43]
port 67 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 la_data_in[44]
port 68 nsew signal input
rlabel metal3 s 29200 11568 30000 11688 6 la_data_in[45]
port 69 nsew signal input
rlabel metal3 s 29200 7488 30000 7608 6 la_data_in[46]
port 70 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 la_data_in[47]
port 71 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 la_data_in[48]
port 72 nsew signal input
rlabel metal3 s 29200 8 30000 128 6 la_data_in[49]
port 73 nsew signal input
rlabel metal3 s 29200 8848 30000 8968 6 la_data_in[4]
port 74 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 la_data_in[50]
port 75 nsew signal input
rlabel metal3 s 29200 4768 30000 4888 6 la_data_in[51]
port 76 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 la_data_in[52]
port 77 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_data_in[53]
port 78 nsew signal input
rlabel metal3 s 0 688 800 808 6 la_data_in[54]
port 79 nsew signal input
rlabel metal3 s 29200 26528 30000 26648 6 la_data_in[55]
port 80 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 la_data_in[56]
port 81 nsew signal input
rlabel metal3 s 29200 2728 30000 2848 6 la_data_in[57]
port 82 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 la_data_in[58]
port 83 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[59]
port 84 nsew signal input
rlabel metal2 s 14830 29200 14886 30000 6 la_data_in[5]
port 85 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_data_in[60]
port 86 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[61]
port 87 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 la_data_in[62]
port 88 nsew signal input
rlabel metal3 s 29200 1368 30000 1488 6 la_data_in[63]
port 89 nsew signal input
rlabel metal3 s 29200 20408 30000 20528 6 la_data_in[64]
port 90 nsew signal input
rlabel metal3 s 29200 12248 30000 12368 6 la_data_in[65]
port 91 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 la_data_in[66]
port 92 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 la_data_in[67]
port 93 nsew signal input
rlabel metal3 s 29200 6128 30000 6248 6 la_data_in[68]
port 94 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 la_data_in[69]
port 95 nsew signal input
rlabel metal3 s 29200 15648 30000 15768 6 la_data_in[6]
port 96 nsew signal input
rlabel metal3 s 29200 23808 30000 23928 6 la_data_in[70]
port 97 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_data_in[71]
port 98 nsew signal input
rlabel metal3 s 29200 25848 30000 25968 6 la_data_in[72]
port 99 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 la_data_in[73]
port 100 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 la_data_in[74]
port 101 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 la_data_in[75]
port 102 nsew signal input
rlabel metal2 s 18 0 74 800 6 la_data_in[76]
port 103 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la_data_in[77]
port 104 nsew signal input
rlabel metal2 s 18 29200 74 30000 6 la_data_in[78]
port 105 nsew signal input
rlabel metal2 s 9034 29200 9090 30000 6 la_data_in[79]
port 106 nsew signal input
rlabel metal2 s 19338 29200 19394 30000 6 la_data_in[7]
port 107 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 la_data_in[80]
port 108 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 la_data_in[81]
port 109 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 la_data_in[82]
port 110 nsew signal input
rlabel metal2 s 23846 29200 23902 30000 6 la_data_in[83]
port 111 nsew signal input
rlabel metal2 s 17406 29200 17462 30000 6 la_data_in[84]
port 112 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 la_data_in[85]
port 113 nsew signal input
rlabel metal2 s 27066 29200 27122 30000 6 la_data_in[86]
port 114 nsew signal input
rlabel metal3 s 29200 4088 30000 4208 6 la_data_in[87]
port 115 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 la_data_in[88]
port 116 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_data_in[89]
port 117 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 la_data_in[8]
port 118 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 la_data_in[90]
port 119 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_data_in[91]
port 120 nsew signal input
rlabel metal3 s 29200 18368 30000 18488 6 la_data_in[92]
port 121 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 la_data_in[93]
port 122 nsew signal input
rlabel metal2 s 22558 29200 22614 30000 6 la_data_in[94]
port 123 nsew signal input
rlabel metal2 s 21914 29200 21970 30000 6 la_data_in[95]
port 124 nsew signal input
rlabel metal2 s 1306 29200 1362 30000 6 la_data_in[96]
port 125 nsew signal input
rlabel metal2 s 5814 29200 5870 30000 6 la_data_in[97]
port 126 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 la_data_in[98]
port 127 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 la_data_in[99]
port 128 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 la_data_in[9]
port 129 nsew signal input
rlabel metal3 s 29200 13608 30000 13728 6 meip
port 130 nsew signal output
rlabel metal4 s 4418 2128 4738 27792 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 11366 2128 11686 27792 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 18314 2128 18634 27792 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 25262 2128 25582 27792 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 7892 2128 8212 27792 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 14840 2128 15160 27792 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 21788 2128 22108 27792 6 vssd1
port 132 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 378226
string GDS_FILE /root/rioschip/openlane/okk/runs/22_09_12_20_58/results/signoff/okk.magic.gds
string GDS_START 35840
<< end >>

