magic
tech sky130B
magscale 1 2
timestamp 1663004140
<< obsli1 >>
rect 1104 2159 88872 27761
<< obsm1 >>
rect 14 1164 89594 27792
<< metal2 >>
rect 18 29200 74 30000
rect 662 29200 718 30000
rect 1306 29200 1362 30000
rect 2594 29200 2650 30000
rect 3238 29200 3294 30000
rect 3882 29200 3938 30000
rect 4526 29200 4582 30000
rect 5170 29200 5226 30000
rect 5814 29200 5870 30000
rect 6458 29200 6514 30000
rect 7102 29200 7158 30000
rect 7746 29200 7802 30000
rect 8390 29200 8446 30000
rect 9034 29200 9090 30000
rect 10322 29200 10378 30000
rect 10966 29200 11022 30000
rect 11610 29200 11666 30000
rect 12254 29200 12310 30000
rect 12898 29200 12954 30000
rect 13542 29200 13598 30000
rect 14186 29200 14242 30000
rect 14830 29200 14886 30000
rect 15474 29200 15530 30000
rect 16118 29200 16174 30000
rect 16762 29200 16818 30000
rect 18050 29200 18106 30000
rect 18694 29200 18750 30000
rect 19338 29200 19394 30000
rect 19982 29200 20038 30000
rect 20626 29200 20682 30000
rect 21270 29200 21326 30000
rect 21914 29200 21970 30000
rect 22558 29200 22614 30000
rect 23202 29200 23258 30000
rect 23846 29200 23902 30000
rect 24490 29200 24546 30000
rect 25778 29200 25834 30000
rect 26422 29200 26478 30000
rect 27066 29200 27122 30000
rect 27710 29200 27766 30000
rect 28354 29200 28410 30000
rect 28998 29200 29054 30000
rect 29642 29200 29698 30000
rect 30286 29200 30342 30000
rect 30930 29200 30986 30000
rect 31574 29200 31630 30000
rect 32862 29200 32918 30000
rect 33506 29200 33562 30000
rect 34150 29200 34206 30000
rect 34794 29200 34850 30000
rect 35438 29200 35494 30000
rect 36082 29200 36138 30000
rect 36726 29200 36782 30000
rect 37370 29200 37426 30000
rect 38014 29200 38070 30000
rect 38658 29200 38714 30000
rect 39302 29200 39358 30000
rect 40590 29200 40646 30000
rect 41234 29200 41290 30000
rect 41878 29200 41934 30000
rect 42522 29200 42578 30000
rect 43166 29200 43222 30000
rect 43810 29200 43866 30000
rect 44454 29200 44510 30000
rect 45098 29200 45154 30000
rect 45742 29200 45798 30000
rect 46386 29200 46442 30000
rect 47030 29200 47086 30000
rect 48318 29200 48374 30000
rect 48962 29200 49018 30000
rect 49606 29200 49662 30000
rect 50250 29200 50306 30000
rect 50894 29200 50950 30000
rect 51538 29200 51594 30000
rect 52182 29200 52238 30000
rect 52826 29200 52882 30000
rect 53470 29200 53526 30000
rect 54114 29200 54170 30000
rect 54758 29200 54814 30000
rect 56046 29200 56102 30000
rect 56690 29200 56746 30000
rect 57334 29200 57390 30000
rect 57978 29200 58034 30000
rect 58622 29200 58678 30000
rect 59266 29200 59322 30000
rect 59910 29200 59966 30000
rect 60554 29200 60610 30000
rect 61198 29200 61254 30000
rect 61842 29200 61898 30000
rect 62486 29200 62542 30000
rect 63774 29200 63830 30000
rect 64418 29200 64474 30000
rect 65062 29200 65118 30000
rect 65706 29200 65762 30000
rect 66350 29200 66406 30000
rect 66994 29200 67050 30000
rect 67638 29200 67694 30000
rect 68282 29200 68338 30000
rect 68926 29200 68982 30000
rect 69570 29200 69626 30000
rect 70214 29200 70270 30000
rect 71502 29200 71558 30000
rect 72146 29200 72202 30000
rect 72790 29200 72846 30000
rect 73434 29200 73490 30000
rect 74078 29200 74134 30000
rect 74722 29200 74778 30000
rect 75366 29200 75422 30000
rect 76010 29200 76066 30000
rect 76654 29200 76710 30000
rect 77298 29200 77354 30000
rect 77942 29200 77998 30000
rect 79230 29200 79286 30000
rect 79874 29200 79930 30000
rect 80518 29200 80574 30000
rect 81162 29200 81218 30000
rect 81806 29200 81862 30000
rect 82450 29200 82506 30000
rect 83094 29200 83150 30000
rect 83738 29200 83794 30000
rect 84382 29200 84438 30000
rect 85026 29200 85082 30000
rect 85670 29200 85726 30000
rect 86958 29200 87014 30000
rect 87602 29200 87658 30000
rect 88246 29200 88302 30000
rect 88890 29200 88946 30000
rect 89534 29200 89590 30000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 84382 0 84438 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 89534 0 89590 800
<< obsm2 >>
rect 130 29144 606 29345
rect 774 29144 1250 29345
rect 1418 29144 2538 29345
rect 2706 29144 3182 29345
rect 3350 29144 3826 29345
rect 3994 29144 4470 29345
rect 4638 29144 5114 29345
rect 5282 29144 5758 29345
rect 5926 29144 6402 29345
rect 6570 29144 7046 29345
rect 7214 29144 7690 29345
rect 7858 29144 8334 29345
rect 8502 29144 8978 29345
rect 9146 29144 10266 29345
rect 10434 29144 10910 29345
rect 11078 29144 11554 29345
rect 11722 29144 12198 29345
rect 12366 29144 12842 29345
rect 13010 29144 13486 29345
rect 13654 29144 14130 29345
rect 14298 29144 14774 29345
rect 14942 29144 15418 29345
rect 15586 29144 16062 29345
rect 16230 29144 16706 29345
rect 16874 29144 17994 29345
rect 18162 29144 18638 29345
rect 18806 29144 19282 29345
rect 19450 29144 19926 29345
rect 20094 29144 20570 29345
rect 20738 29144 21214 29345
rect 21382 29144 21858 29345
rect 22026 29144 22502 29345
rect 22670 29144 23146 29345
rect 23314 29144 23790 29345
rect 23958 29144 24434 29345
rect 24602 29144 25722 29345
rect 25890 29144 26366 29345
rect 26534 29144 27010 29345
rect 27178 29144 27654 29345
rect 27822 29144 28298 29345
rect 28466 29144 28942 29345
rect 29110 29144 29586 29345
rect 29754 29144 30230 29345
rect 30398 29144 30874 29345
rect 31042 29144 31518 29345
rect 31686 29144 32806 29345
rect 32974 29144 33450 29345
rect 33618 29144 34094 29345
rect 34262 29144 34738 29345
rect 34906 29144 35382 29345
rect 35550 29144 36026 29345
rect 36194 29144 36670 29345
rect 36838 29144 37314 29345
rect 37482 29144 37958 29345
rect 38126 29144 38602 29345
rect 38770 29144 39246 29345
rect 39414 29144 40534 29345
rect 40702 29144 41178 29345
rect 41346 29144 41822 29345
rect 41990 29144 42466 29345
rect 42634 29144 43110 29345
rect 43278 29144 43754 29345
rect 43922 29144 44398 29345
rect 44566 29144 45042 29345
rect 45210 29144 45686 29345
rect 45854 29144 46330 29345
rect 46498 29144 46974 29345
rect 47142 29144 48262 29345
rect 48430 29144 48906 29345
rect 49074 29144 49550 29345
rect 49718 29144 50194 29345
rect 50362 29144 50838 29345
rect 51006 29144 51482 29345
rect 51650 29144 52126 29345
rect 52294 29144 52770 29345
rect 52938 29144 53414 29345
rect 53582 29144 54058 29345
rect 54226 29144 54702 29345
rect 54870 29144 55990 29345
rect 56158 29144 56634 29345
rect 56802 29144 57278 29345
rect 57446 29144 57922 29345
rect 58090 29144 58566 29345
rect 58734 29144 59210 29345
rect 59378 29144 59854 29345
rect 60022 29144 60498 29345
rect 60666 29144 61142 29345
rect 61310 29144 61786 29345
rect 61954 29144 62430 29345
rect 62598 29144 63718 29345
rect 63886 29144 64362 29345
rect 64530 29144 65006 29345
rect 65174 29144 65650 29345
rect 65818 29144 66294 29345
rect 66462 29144 66938 29345
rect 67106 29144 67582 29345
rect 67750 29144 68226 29345
rect 68394 29144 68870 29345
rect 69038 29144 69514 29345
rect 69682 29144 70158 29345
rect 70326 29144 71446 29345
rect 71614 29144 72090 29345
rect 72258 29144 72734 29345
rect 72902 29144 73378 29345
rect 73546 29144 74022 29345
rect 74190 29144 74666 29345
rect 74834 29144 75310 29345
rect 75478 29144 75954 29345
rect 76122 29144 76598 29345
rect 76766 29144 77242 29345
rect 77410 29144 77886 29345
rect 78054 29144 79174 29345
rect 79342 29144 79818 29345
rect 79986 29144 80462 29345
rect 80630 29144 81106 29345
rect 81274 29144 81750 29345
rect 81918 29144 82394 29345
rect 82562 29144 83038 29345
rect 83206 29144 83682 29345
rect 83850 29144 84326 29345
rect 84494 29144 84970 29345
rect 85138 29144 85614 29345
rect 85782 29144 86902 29345
rect 87070 29144 87546 29345
rect 87714 29144 88190 29345
rect 88358 29144 88834 29345
rect 89002 29144 89478 29345
rect 20 856 89588 29144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 2538 856
rect 2706 31 3182 856
rect 3350 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7690 856
rect 7858 31 8334 856
rect 8502 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14130 856
rect 14298 31 15418 856
rect 15586 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17350 856
rect 17518 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 20570 856
rect 20738 31 21214 856
rect 21382 31 21858 856
rect 22026 31 23146 856
rect 23314 31 23790 856
rect 23958 31 24434 856
rect 24602 31 25078 856
rect 25246 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28298 856
rect 28466 31 28942 856
rect 29110 31 29586 856
rect 29754 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32162 856
rect 32330 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34094 856
rect 34262 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36026 856
rect 36194 31 36670 856
rect 36838 31 37314 856
rect 37482 31 38602 856
rect 38770 31 39246 856
rect 39414 31 39890 856
rect 40058 31 40534 856
rect 40702 31 41178 856
rect 41346 31 41822 856
rect 41990 31 42466 856
rect 42634 31 43110 856
rect 43278 31 43754 856
rect 43922 31 44398 856
rect 44566 31 45042 856
rect 45210 31 46330 856
rect 46498 31 46974 856
rect 47142 31 47618 856
rect 47786 31 48262 856
rect 48430 31 48906 856
rect 49074 31 49550 856
rect 49718 31 50194 856
rect 50362 31 50838 856
rect 51006 31 51482 856
rect 51650 31 52126 856
rect 52294 31 52770 856
rect 52938 31 54058 856
rect 54226 31 54702 856
rect 54870 31 55346 856
rect 55514 31 55990 856
rect 56158 31 56634 856
rect 56802 31 57278 856
rect 57446 31 57922 856
rect 58090 31 58566 856
rect 58734 31 59210 856
rect 59378 31 59854 856
rect 60022 31 61142 856
rect 61310 31 61786 856
rect 61954 31 62430 856
rect 62598 31 63074 856
rect 63242 31 63718 856
rect 63886 31 64362 856
rect 64530 31 65006 856
rect 65174 31 65650 856
rect 65818 31 66294 856
rect 66462 31 66938 856
rect 67106 31 67582 856
rect 67750 31 68870 856
rect 69038 31 69514 856
rect 69682 31 70158 856
rect 70326 31 70802 856
rect 70970 31 71446 856
rect 71614 31 72090 856
rect 72258 31 72734 856
rect 72902 31 73378 856
rect 73546 31 74022 856
rect 74190 31 74666 856
rect 74834 31 75310 856
rect 75478 31 76598 856
rect 76766 31 77242 856
rect 77410 31 77886 856
rect 78054 31 78530 856
rect 78698 31 79174 856
rect 79342 31 79818 856
rect 79986 31 80462 856
rect 80630 31 81106 856
rect 81274 31 81750 856
rect 81918 31 82394 856
rect 82562 31 83038 856
rect 83206 31 84326 856
rect 84494 31 84970 856
rect 85138 31 85614 856
rect 85782 31 86258 856
rect 86426 31 86902 856
rect 87070 31 87546 856
rect 87714 31 88190 856
rect 88358 31 88834 856
rect 89002 31 89478 856
<< metal3 >>
rect 0 29248 800 29368
rect 89200 29248 90000 29368
rect 0 28568 800 28688
rect 89200 28568 90000 28688
rect 0 27888 800 28008
rect 89200 27888 90000 28008
rect 0 27208 800 27328
rect 89200 27208 90000 27328
rect 0 26528 800 26648
rect 89200 26528 90000 26648
rect 0 25848 800 25968
rect 0 25168 800 25288
rect 89200 25168 90000 25288
rect 0 24488 800 24608
rect 89200 24488 90000 24608
rect 89200 23808 90000 23928
rect 0 23128 800 23248
rect 89200 23128 90000 23248
rect 0 22448 800 22568
rect 89200 22448 90000 22568
rect 0 21768 800 21888
rect 89200 21768 90000 21888
rect 0 21088 800 21208
rect 89200 21088 90000 21208
rect 0 20408 800 20528
rect 89200 20408 90000 20528
rect 0 19728 800 19848
rect 89200 19728 90000 19848
rect 0 19048 800 19168
rect 89200 19048 90000 19168
rect 0 18368 800 18488
rect 89200 18368 90000 18488
rect 0 17688 800 17808
rect 0 17008 800 17128
rect 89200 17008 90000 17128
rect 0 16328 800 16448
rect 89200 16328 90000 16448
rect 89200 15648 90000 15768
rect 0 14968 800 15088
rect 89200 14968 90000 15088
rect 0 14288 800 14408
rect 89200 14288 90000 14408
rect 0 13608 800 13728
rect 89200 13608 90000 13728
rect 0 12928 800 13048
rect 89200 12928 90000 13048
rect 0 12248 800 12368
rect 89200 12248 90000 12368
rect 0 11568 800 11688
rect 89200 11568 90000 11688
rect 0 10888 800 11008
rect 89200 10888 90000 11008
rect 0 10208 800 10328
rect 89200 10208 90000 10328
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 89200 8848 90000 8968
rect 0 8168 800 8288
rect 89200 8168 90000 8288
rect 89200 7488 90000 7608
rect 0 6808 800 6928
rect 89200 6808 90000 6928
rect 0 6128 800 6248
rect 89200 6128 90000 6248
rect 0 5448 800 5568
rect 89200 5448 90000 5568
rect 0 4768 800 4888
rect 89200 4768 90000 4888
rect 0 4088 800 4208
rect 89200 4088 90000 4208
rect 0 3408 800 3528
rect 89200 3408 90000 3528
rect 0 2728 800 2848
rect 89200 2728 90000 2848
rect 0 2048 800 2168
rect 89200 2048 90000 2168
rect 0 1368 800 1488
rect 0 688 800 808
rect 89200 688 90000 808
rect 89200 8 90000 128
<< obsm3 >>
rect 880 29168 89120 29341
rect 800 28768 89200 29168
rect 880 28488 89120 28768
rect 800 28088 89200 28488
rect 880 27808 89120 28088
rect 800 27408 89200 27808
rect 880 27128 89120 27408
rect 800 26728 89200 27128
rect 880 26448 89120 26728
rect 800 26048 89200 26448
rect 880 25768 89200 26048
rect 800 25368 89200 25768
rect 880 25088 89120 25368
rect 800 24688 89200 25088
rect 880 24408 89120 24688
rect 800 24008 89200 24408
rect 800 23728 89120 24008
rect 800 23328 89200 23728
rect 880 23048 89120 23328
rect 800 22648 89200 23048
rect 880 22368 89120 22648
rect 800 21968 89200 22368
rect 880 21688 89120 21968
rect 800 21288 89200 21688
rect 880 21008 89120 21288
rect 800 20608 89200 21008
rect 880 20328 89120 20608
rect 800 19928 89200 20328
rect 880 19648 89120 19928
rect 800 19248 89200 19648
rect 880 18968 89120 19248
rect 800 18568 89200 18968
rect 880 18288 89120 18568
rect 800 17888 89200 18288
rect 880 17608 89200 17888
rect 800 17208 89200 17608
rect 880 16928 89120 17208
rect 800 16528 89200 16928
rect 880 16248 89120 16528
rect 800 15848 89200 16248
rect 800 15568 89120 15848
rect 800 15168 89200 15568
rect 880 14888 89120 15168
rect 800 14488 89200 14888
rect 880 14208 89120 14488
rect 800 13808 89200 14208
rect 880 13528 89120 13808
rect 800 13128 89200 13528
rect 880 12848 89120 13128
rect 800 12448 89200 12848
rect 880 12168 89120 12448
rect 800 11768 89200 12168
rect 880 11488 89120 11768
rect 800 11088 89200 11488
rect 880 10808 89120 11088
rect 800 10408 89200 10808
rect 880 10128 89120 10408
rect 800 9728 89200 10128
rect 880 9448 89200 9728
rect 800 9048 89200 9448
rect 880 8768 89120 9048
rect 800 8368 89200 8768
rect 880 8088 89120 8368
rect 800 7688 89200 8088
rect 800 7408 89120 7688
rect 800 7008 89200 7408
rect 880 6728 89120 7008
rect 800 6328 89200 6728
rect 880 6048 89120 6328
rect 800 5648 89200 6048
rect 880 5368 89120 5648
rect 800 4968 89200 5368
rect 880 4688 89120 4968
rect 800 4288 89200 4688
rect 880 4008 89120 4288
rect 800 3608 89200 4008
rect 880 3328 89120 3608
rect 800 2928 89200 3328
rect 880 2648 89120 2928
rect 800 2248 89200 2648
rect 880 1968 89120 2248
rect 800 1568 89200 1968
rect 880 1288 89200 1568
rect 800 888 89200 1288
rect 880 608 89120 888
rect 800 208 89200 608
rect 800 35 89120 208
<< metal4 >>
rect 11918 2128 12238 27792
rect 22892 2128 23212 27792
rect 33866 2128 34186 27792
rect 44840 2128 45160 27792
rect 55814 2128 56134 27792
rect 66788 2128 67108 27792
rect 77762 2128 78082 27792
<< obsm4 >>
rect 26555 10235 33786 25805
rect 34266 10235 44760 25805
rect 45240 10235 55734 25805
rect 56214 10235 64341 25805
<< labels >>
rlabel metal2 s 41234 0 41290 800 6 clk
port 1 nsew signal input
rlabel metal2 s 5170 29200 5226 30000 6 data_chip_en
port 2 nsew signal output
rlabel metal3 s 89200 7488 90000 7608 6 data_in[0]
port 3 nsew signal output
rlabel metal2 s 35438 29200 35494 30000 6 data_in[10]
port 4 nsew signal output
rlabel metal3 s 89200 11568 90000 11688 6 data_in[11]
port 5 nsew signal output
rlabel metal2 s 14830 29200 14886 30000 6 data_in[12]
port 6 nsew signal output
rlabel metal2 s 72146 29200 72202 30000 6 data_in[13]
port 7 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 data_in[14]
port 8 nsew signal output
rlabel metal2 s 42522 29200 42578 30000 6 data_in[15]
port 9 nsew signal output
rlabel metal2 s 34794 29200 34850 30000 6 data_in[16]
port 10 nsew signal output
rlabel metal2 s 10322 29200 10378 30000 6 data_in[17]
port 11 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 data_in[18]
port 12 nsew signal output
rlabel metal2 s 52182 29200 52238 30000 6 data_in[19]
port 13 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 data_in[1]
port 14 nsew signal output
rlabel metal2 s 662 29200 718 30000 6 data_in[20]
port 15 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 data_in[21]
port 16 nsew signal output
rlabel metal2 s 18 29200 74 30000 6 data_in[22]
port 17 nsew signal output
rlabel metal2 s 61842 29200 61898 30000 6 data_in[23]
port 18 nsew signal output
rlabel metal2 s 45742 29200 45798 30000 6 data_in[24]
port 19 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 data_in[25]
port 20 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 data_in[26]
port 21 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 data_in[27]
port 22 nsew signal output
rlabel metal2 s 71502 29200 71558 30000 6 data_in[28]
port 23 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 data_in[29]
port 24 nsew signal output
rlabel metal2 s 33506 29200 33562 30000 6 data_in[2]
port 25 nsew signal output
rlabel metal2 s 19982 29200 20038 30000 6 data_in[30]
port 26 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 data_in[31]
port 27 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 data_in[3]
port 28 nsew signal output
rlabel metal2 s 65062 29200 65118 30000 6 data_in[4]
port 29 nsew signal output
rlabel metal2 s 7102 29200 7158 30000 6 data_in[5]
port 30 nsew signal output
rlabel metal2 s 38658 29200 38714 30000 6 data_in[6]
port 31 nsew signal output
rlabel metal2 s 39302 29200 39358 30000 6 data_in[7]
port 32 nsew signal output
rlabel metal2 s 77298 29200 77354 30000 6 data_in[8]
port 33 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 data_in[9]
port 34 nsew signal output
rlabel metal2 s 36082 29200 36138 30000 6 data_index[0]
port 35 nsew signal output
rlabel metal3 s 89200 21088 90000 21208 6 data_index[1]
port 36 nsew signal output
rlabel metal2 s 81806 29200 81862 30000 6 data_index[2]
port 37 nsew signal output
rlabel metal3 s 89200 28568 90000 28688 6 data_index[3]
port 38 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 data_index[4]
port 39 nsew signal output
rlabel metal2 s 15474 29200 15530 30000 6 data_index[5]
port 40 nsew signal output
rlabel metal2 s 74078 29200 74134 30000 6 data_index[6]
port 41 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 data_index[7]
port 42 nsew signal output
rlabel metal2 s 16118 29200 16174 30000 6 data_out[0]
port 43 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 data_out[10]
port 44 nsew signal input
rlabel metal3 s 89200 26528 90000 26648 6 data_out[11]
port 45 nsew signal input
rlabel metal2 s 12898 29200 12954 30000 6 data_out[12]
port 46 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 data_out[13]
port 47 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 data_out[14]
port 48 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 data_out[15]
port 49 nsew signal input
rlabel metal2 s 41878 29200 41934 30000 6 data_out[16]
port 50 nsew signal input
rlabel metal3 s 89200 8848 90000 8968 6 data_out[17]
port 51 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 data_out[18]
port 52 nsew signal input
rlabel metal2 s 6458 29200 6514 30000 6 data_out[19]
port 53 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 data_out[1]
port 54 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 data_out[20]
port 55 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 data_out[21]
port 56 nsew signal input
rlabel metal2 s 11610 29200 11666 30000 6 data_out[22]
port 57 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 data_out[23]
port 58 nsew signal input
rlabel metal2 s 87602 29200 87658 30000 6 data_out[24]
port 59 nsew signal input
rlabel metal3 s 89200 8168 90000 8288 6 data_out[25]
port 60 nsew signal input
rlabel metal2 s 83738 29200 83794 30000 6 data_out[26]
port 61 nsew signal input
rlabel metal2 s 23846 29200 23902 30000 6 data_out[27]
port 62 nsew signal input
rlabel metal2 s 21270 29200 21326 30000 6 data_out[28]
port 63 nsew signal input
rlabel metal2 s 85026 29200 85082 30000 6 data_out[29]
port 64 nsew signal input
rlabel metal2 s 4526 29200 4582 30000 6 data_out[2]
port 65 nsew signal input
rlabel metal3 s 89200 6808 90000 6928 6 data_out[30]
port 66 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 data_out[31]
port 67 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 data_out[3]
port 68 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 data_out[4]
port 69 nsew signal input
rlabel metal2 s 51538 29200 51594 30000 6 data_out[5]
port 70 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 data_out[6]
port 71 nsew signal input
rlabel metal3 s 89200 10888 90000 11008 6 data_out[7]
port 72 nsew signal input
rlabel metal2 s 30930 29200 30986 30000 6 data_out[8]
port 73 nsew signal input
rlabel metal2 s 54114 29200 54170 30000 6 data_out[9]
port 74 nsew signal input
rlabel metal2 s 88246 29200 88302 30000 6 data_write_en
port 75 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 ld_data_o[0]
port 76 nsew signal output
rlabel metal2 s 74722 29200 74778 30000 6 ld_data_o[10]
port 77 nsew signal output
rlabel metal3 s 89200 2728 90000 2848 6 ld_data_o[11]
port 78 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 ld_data_o[12]
port 79 nsew signal output
rlabel metal2 s 43810 29200 43866 30000 6 ld_data_o[13]
port 80 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 ld_data_o[14]
port 81 nsew signal output
rlabel metal3 s 89200 19048 90000 19168 6 ld_data_o[15]
port 82 nsew signal output
rlabel metal2 s 45098 29200 45154 30000 6 ld_data_o[16]
port 83 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 ld_data_o[17]
port 84 nsew signal output
rlabel metal2 s 9034 29200 9090 30000 6 ld_data_o[18]
port 85 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 ld_data_o[19]
port 86 nsew signal output
rlabel metal3 s 89200 13608 90000 13728 6 ld_data_o[1]
port 87 nsew signal output
rlabel metal2 s 72790 29200 72846 30000 6 ld_data_o[20]
port 88 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 ld_data_o[21]
port 89 nsew signal output
rlabel metal3 s 89200 4768 90000 4888 6 ld_data_o[22]
port 90 nsew signal output
rlabel metal2 s 88890 29200 88946 30000 6 ld_data_o[23]
port 91 nsew signal output
rlabel metal2 s 69570 29200 69626 30000 6 ld_data_o[24]
port 92 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 ld_data_o[25]
port 93 nsew signal output
rlabel metal2 s 59266 29200 59322 30000 6 ld_data_o[26]
port 94 nsew signal output
rlabel metal3 s 89200 4088 90000 4208 6 ld_data_o[27]
port 95 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 ld_data_o[28]
port 96 nsew signal output
rlabel metal2 s 86958 29200 87014 30000 6 ld_data_o[29]
port 97 nsew signal output
rlabel metal2 s 62486 29200 62542 30000 6 ld_data_o[2]
port 98 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 ld_data_o[30]
port 99 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 ld_data_o[31]
port 100 nsew signal output
rlabel metal3 s 89200 8 90000 128 6 ld_data_o[3]
port 101 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 ld_data_o[4]
port 102 nsew signal output
rlabel metal2 s 50894 29200 50950 30000 6 ld_data_o[5]
port 103 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 ld_data_o[6]
port 104 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 ld_data_o[7]
port 105 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 ld_data_o[8]
port 106 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 ld_data_o[9]
port 107 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 req_addr_i[0]
port 108 nsew signal input
rlabel metal2 s 79874 29200 79930 30000 6 req_addr_i[10]
port 109 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 req_addr_i[11]
port 110 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 req_addr_i[12]
port 111 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 req_addr_i[13]
port 112 nsew signal input
rlabel metal2 s 44454 29200 44510 30000 6 req_addr_i[14]
port 113 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 req_addr_i[15]
port 114 nsew signal input
rlabel metal2 s 28998 29200 29054 30000 6 req_addr_i[16]
port 115 nsew signal input
rlabel metal2 s 22558 29200 22614 30000 6 req_addr_i[17]
port 116 nsew signal input
rlabel metal2 s 66994 29200 67050 30000 6 req_addr_i[18]
port 117 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 req_addr_i[19]
port 118 nsew signal input
rlabel metal2 s 53470 29200 53526 30000 6 req_addr_i[1]
port 119 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 req_addr_i[20]
port 120 nsew signal input
rlabel metal3 s 89200 6128 90000 6248 6 req_addr_i[21]
port 121 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 req_addr_i[22]
port 122 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 req_addr_i[23]
port 123 nsew signal input
rlabel metal3 s 89200 18368 90000 18488 6 req_addr_i[24]
port 124 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 req_addr_i[25]
port 125 nsew signal input
rlabel metal2 s 36726 29200 36782 30000 6 req_addr_i[26]
port 126 nsew signal input
rlabel metal2 s 28354 29200 28410 30000 6 req_addr_i[27]
port 127 nsew signal input
rlabel metal2 s 16762 29200 16818 30000 6 req_addr_i[28]
port 128 nsew signal input
rlabel metal2 s 82450 29200 82506 30000 6 req_addr_i[29]
port 129 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 req_addr_i[2]
port 130 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 req_addr_i[30]
port 131 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 req_addr_i[31]
port 132 nsew signal input
rlabel metal2 s 1306 29200 1362 30000 6 req_addr_i[3]
port 133 nsew signal input
rlabel metal2 s 89534 29200 89590 30000 6 req_addr_i[4]
port 134 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 req_addr_i[5]
port 135 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 req_addr_i[6]
port 136 nsew signal input
rlabel metal2 s 23202 29200 23258 30000 6 req_addr_i[7]
port 137 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 req_addr_i[8]
port 138 nsew signal input
rlabel metal2 s 67638 29200 67694 30000 6 req_addr_i[9]
port 139 nsew signal input
rlabel metal3 s 89200 23128 90000 23248 6 req_ready_o
port 140 nsew signal output
rlabel metal2 s 68282 29200 68338 30000 6 req_valid_i
port 141 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 resp_addr_o[0]
port 142 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 resp_addr_o[10]
port 143 nsew signal output
rlabel metal2 s 21914 29200 21970 30000 6 resp_addr_o[11]
port 144 nsew signal output
rlabel metal3 s 89200 21768 90000 21888 6 resp_addr_o[12]
port 145 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 resp_addr_o[13]
port 146 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 resp_addr_o[14]
port 147 nsew signal output
rlabel metal2 s 75366 29200 75422 30000 6 resp_addr_o[15]
port 148 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 resp_addr_o[16]
port 149 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 resp_addr_o[17]
port 150 nsew signal output
rlabel metal2 s 56690 29200 56746 30000 6 resp_addr_o[18]
port 151 nsew signal output
rlabel metal2 s 85670 29200 85726 30000 6 resp_addr_o[19]
port 152 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 resp_addr_o[1]
port 153 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 resp_addr_o[20]
port 154 nsew signal output
rlabel metal2 s 48962 29200 49018 30000 6 resp_addr_o[21]
port 155 nsew signal output
rlabel metal3 s 89200 16328 90000 16448 6 resp_addr_o[22]
port 156 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 resp_addr_o[23]
port 157 nsew signal output
rlabel metal2 s 65706 29200 65762 30000 6 resp_addr_o[24]
port 158 nsew signal output
rlabel metal2 s 60554 29200 60610 30000 6 resp_addr_o[25]
port 159 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 resp_addr_o[26]
port 160 nsew signal output
rlabel metal2 s 56046 29200 56102 30000 6 resp_addr_o[27]
port 161 nsew signal output
rlabel metal2 s 41234 29200 41290 30000 6 resp_addr_o[28]
port 162 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 resp_addr_o[29]
port 163 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 resp_addr_o[2]
port 164 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 resp_addr_o[30]
port 165 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 resp_addr_o[31]
port 166 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 resp_addr_o[3]
port 167 nsew signal output
rlabel metal2 s 46386 29200 46442 30000 6 resp_addr_o[4]
port 168 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 resp_addr_o[5]
port 169 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 resp_addr_o[6]
port 170 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 resp_addr_o[7]
port 171 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 resp_addr_o[8]
port 172 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 resp_addr_o[9]
port 173 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 resp_ready_i
port 174 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 resp_valid_o
port 175 nsew signal output
rlabel metal3 s 89200 14968 90000 15088 6 rstn
port 176 nsew signal input
rlabel metal2 s 43166 29200 43222 30000 6 tag_chip_en
port 177 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 tag_data_in[0]
port 178 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 tag_data_in[10]
port 179 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 tag_data_in[11]
port 180 nsew signal output
rlabel metal2 s 34150 29200 34206 30000 6 tag_data_in[12]
port 181 nsew signal output
rlabel metal2 s 14186 29200 14242 30000 6 tag_data_in[13]
port 182 nsew signal output
rlabel metal2 s 2594 29200 2650 30000 6 tag_data_in[14]
port 183 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 tag_data_in[15]
port 184 nsew signal output
rlabel metal3 s 89200 10208 90000 10328 6 tag_data_in[16]
port 185 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 tag_data_in[17]
port 186 nsew signal output
rlabel metal2 s 32862 29200 32918 30000 6 tag_data_in[18]
port 187 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 tag_data_in[19]
port 188 nsew signal output
rlabel metal3 s 89200 3408 90000 3528 6 tag_data_in[1]
port 189 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 tag_data_in[20]
port 190 nsew signal output
rlabel metal3 s 89200 19728 90000 19848 6 tag_data_in[21]
port 191 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 tag_data_in[22]
port 192 nsew signal output
rlabel metal2 s 662 0 718 800 6 tag_data_in[23]
port 193 nsew signal output
rlabel metal2 s 64418 29200 64474 30000 6 tag_data_in[24]
port 194 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 tag_data_in[25]
port 195 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 tag_data_in[26]
port 196 nsew signal output
rlabel metal3 s 89200 17008 90000 17128 6 tag_data_in[27]
port 197 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 tag_data_in[28]
port 198 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 tag_data_in[29]
port 199 nsew signal output
rlabel metal2 s 18050 29200 18106 30000 6 tag_data_in[2]
port 200 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 tag_data_in[30]
port 201 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 tag_data_in[31]
port 202 nsew signal output
rlabel metal3 s 89200 24488 90000 24608 6 tag_data_in[3]
port 203 nsew signal output
rlabel metal2 s 24490 29200 24546 30000 6 tag_data_in[4]
port 204 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 tag_data_in[5]
port 205 nsew signal output
rlabel metal2 s 3882 29200 3938 30000 6 tag_data_in[6]
port 206 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 tag_data_in[7]
port 207 nsew signal output
rlabel metal2 s 38014 29200 38070 30000 6 tag_data_in[8]
port 208 nsew signal output
rlabel metal2 s 57978 29200 58034 30000 6 tag_data_in[9]
port 209 nsew signal output
rlabel metal2 s 66350 29200 66406 30000 6 tag_index[0]
port 210 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 tag_index[1]
port 211 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 tag_index[2]
port 212 nsew signal output
rlabel metal2 s 18694 29200 18750 30000 6 tag_index[3]
port 213 nsew signal output
rlabel metal2 s 52826 29200 52882 30000 6 tag_index[4]
port 214 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 tag_index[5]
port 215 nsew signal output
rlabel metal3 s 89200 23808 90000 23928 6 tag_index[6]
port 216 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 tag_index[7]
port 217 nsew signal output
rlabel metal2 s 79230 29200 79286 30000 6 tag_out[0]
port 218 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 tag_out[10]
port 219 nsew signal input
rlabel metal2 s 30286 29200 30342 30000 6 tag_out[11]
port 220 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 tag_out[12]
port 221 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 tag_out[13]
port 222 nsew signal input
rlabel metal2 s 31574 29200 31630 30000 6 tag_out[14]
port 223 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 tag_out[15]
port 224 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 tag_out[16]
port 225 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 tag_out[17]
port 226 nsew signal input
rlabel metal2 s 61198 29200 61254 30000 6 tag_out[18]
port 227 nsew signal input
rlabel metal3 s 89200 27208 90000 27328 6 tag_out[19]
port 228 nsew signal input
rlabel metal2 s 10966 29200 11022 30000 6 tag_out[1]
port 229 nsew signal input
rlabel metal2 s 58622 29200 58678 30000 6 tag_out[20]
port 230 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 tag_out[21]
port 231 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 tag_out[22]
port 232 nsew signal input
rlabel metal2 s 54758 29200 54814 30000 6 tag_out[23]
port 233 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 tag_out[24]
port 234 nsew signal input
rlabel metal2 s 80518 29200 80574 30000 6 tag_out[25]
port 235 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 tag_out[26]
port 236 nsew signal input
rlabel metal2 s 47030 29200 47086 30000 6 tag_out[27]
port 237 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 tag_out[28]
port 238 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 tag_out[29]
port 239 nsew signal input
rlabel metal3 s 89200 5448 90000 5568 6 tag_out[2]
port 240 nsew signal input
rlabel metal2 s 5814 29200 5870 30000 6 tag_out[30]
port 241 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 tag_out[31]
port 242 nsew signal input
rlabel metal2 s 19338 29200 19394 30000 6 tag_out[3]
port 243 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 tag_out[4]
port 244 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 tag_out[5]
port 245 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 tag_out[6]
port 246 nsew signal input
rlabel metal3 s 89200 25168 90000 25288 6 tag_out[7]
port 247 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 tag_out[8]
port 248 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 tag_out[9]
port 249 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 tag_write_en
port 250 nsew signal output
rlabel metal4 s 11918 2128 12238 27792 6 vccd1
port 251 nsew power bidirectional
rlabel metal4 s 33866 2128 34186 27792 6 vccd1
port 251 nsew power bidirectional
rlabel metal4 s 55814 2128 56134 27792 6 vccd1
port 251 nsew power bidirectional
rlabel metal4 s 77762 2128 78082 27792 6 vccd1
port 251 nsew power bidirectional
rlabel metal4 s 22892 2128 23212 27792 6 vssd1
port 252 nsew ground bidirectional
rlabel metal4 s 44840 2128 45160 27792 6 vssd1
port 252 nsew ground bidirectional
rlabel metal4 s 66788 2128 67108 27792 6 vssd1
port 252 nsew ground bidirectional
rlabel metal2 s 48318 29200 48374 30000 6 wb_ack_i
port 253 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wb_adr_o[0]
port 254 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 wb_adr_o[10]
port 255 nsew signal output
rlabel metal2 s 59910 29200 59966 30000 6 wb_adr_o[11]
port 256 nsew signal output
rlabel metal3 s 0 688 800 808 6 wb_adr_o[12]
port 257 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 wb_adr_o[13]
port 258 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 wb_adr_o[14]
port 259 nsew signal output
rlabel metal2 s 7746 29200 7802 30000 6 wb_adr_o[15]
port 260 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 wb_adr_o[16]
port 261 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 wb_adr_o[17]
port 262 nsew signal output
rlabel metal2 s 83094 29200 83150 30000 6 wb_adr_o[18]
port 263 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 wb_adr_o[19]
port 264 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wb_adr_o[1]
port 265 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wb_adr_o[20]
port 266 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 wb_adr_o[21]
port 267 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 wb_adr_o[22]
port 268 nsew signal output
rlabel metal2 s 57334 29200 57390 30000 6 wb_adr_o[23]
port 269 nsew signal output
rlabel metal3 s 89200 15648 90000 15768 6 wb_adr_o[24]
port 270 nsew signal output
rlabel metal2 s 26422 29200 26478 30000 6 wb_adr_o[25]
port 271 nsew signal output
rlabel metal2 s 29642 29200 29698 30000 6 wb_adr_o[26]
port 272 nsew signal output
rlabel metal2 s 27710 29200 27766 30000 6 wb_adr_o[27]
port 273 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 wb_adr_o[28]
port 274 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 wb_adr_o[29]
port 275 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 wb_adr_o[2]
port 276 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wb_adr_o[30]
port 277 nsew signal output
rlabel metal2 s 76654 29200 76710 30000 6 wb_adr_o[31]
port 278 nsew signal output
rlabel metal3 s 89200 29248 90000 29368 6 wb_adr_o[3]
port 279 nsew signal output
rlabel metal2 s 40590 29200 40646 30000 6 wb_adr_o[4]
port 280 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wb_adr_o[5]
port 281 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 wb_adr_o[6]
port 282 nsew signal output
rlabel metal3 s 89200 27888 90000 28008 6 wb_adr_o[7]
port 283 nsew signal output
rlabel metal2 s 13542 29200 13598 30000 6 wb_adr_o[8]
port 284 nsew signal output
rlabel metal3 s 89200 12248 90000 12368 6 wb_adr_o[9]
port 285 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 wb_bl_o[0]
port 286 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 wb_bl_o[1]
port 287 nsew signal output
rlabel metal2 s 84382 29200 84438 30000 6 wb_bl_o[2]
port 288 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 wb_bl_o[3]
port 289 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wb_bl_o[4]
port 290 nsew signal output
rlabel metal3 s 89200 2048 90000 2168 6 wb_bl_o[5]
port 291 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 wb_bl_o[6]
port 292 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 wb_bl_o[7]
port 293 nsew signal output
rlabel metal2 s 8390 29200 8446 30000 6 wb_bl_o[8]
port 294 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 wb_bl_o[9]
port 295 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wb_bry_o
port 296 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wb_cyc_o
port 297 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 wb_dat_i[0]
port 298 nsew signal input
rlabel metal2 s 81162 29200 81218 30000 6 wb_dat_i[10]
port 299 nsew signal input
rlabel metal3 s 89200 20408 90000 20528 6 wb_dat_i[11]
port 300 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wb_dat_i[12]
port 301 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 wb_dat_i[13]
port 302 nsew signal input
rlabel metal3 s 89200 688 90000 808 6 wb_dat_i[14]
port 303 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wb_dat_i[15]
port 304 nsew signal input
rlabel metal3 s 89200 22448 90000 22568 6 wb_dat_i[16]
port 305 nsew signal input
rlabel metal2 s 77942 29200 77998 30000 6 wb_dat_i[17]
port 306 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wb_dat_i[18]
port 307 nsew signal input
rlabel metal2 s 76010 29200 76066 30000 6 wb_dat_i[19]
port 308 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 wb_dat_i[1]
port 309 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wb_dat_i[20]
port 310 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wb_dat_i[21]
port 311 nsew signal input
rlabel metal2 s 18 0 74 800 6 wb_dat_i[22]
port 312 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wb_dat_i[23]
port 313 nsew signal input
rlabel metal2 s 3238 29200 3294 30000 6 wb_dat_i[24]
port 314 nsew signal input
rlabel metal2 s 25778 29200 25834 30000 6 wb_dat_i[25]
port 315 nsew signal input
rlabel metal2 s 49606 29200 49662 30000 6 wb_dat_i[26]
port 316 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_dat_i[27]
port 317 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wb_dat_i[28]
port 318 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wb_dat_i[29]
port 319 nsew signal input
rlabel metal2 s 63774 29200 63830 30000 6 wb_dat_i[2]
port 320 nsew signal input
rlabel metal2 s 50250 29200 50306 30000 6 wb_dat_i[30]
port 321 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wb_dat_i[31]
port 322 nsew signal input
rlabel metal2 s 73434 29200 73490 30000 6 wb_dat_i[3]
port 323 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 wb_dat_i[4]
port 324 nsew signal input
rlabel metal2 s 12254 29200 12310 30000 6 wb_dat_i[5]
port 325 nsew signal input
rlabel metal3 s 89200 14288 90000 14408 6 wb_dat_i[6]
port 326 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wb_dat_i[7]
port 327 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wb_dat_i[8]
port 328 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wb_dat_i[9]
port 329 nsew signal input
rlabel metal3 s 89200 12928 90000 13048 6 wb_stb_o
port 330 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wb_we_o
port 331 nsew signal output
rlabel metal2 s 70214 29200 70270 30000 6 write_data_mask[0]
port 332 nsew signal output
rlabel metal2 s 68926 29200 68982 30000 6 write_data_mask[1]
port 333 nsew signal output
rlabel metal2 s 27066 29200 27122 30000 6 write_data_mask[2]
port 334 nsew signal output
rlabel metal2 s 37370 29200 37426 30000 6 write_data_mask[3]
port 335 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 write_tag_mask[0]
port 336 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 write_tag_mask[1]
port 337 nsew signal output
rlabel metal2 s 20626 29200 20682 30000 6 write_tag_mask[2]
port 338 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 write_tag_mask[3]
port 339 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 90000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3631518
string GDS_FILE /root/hellochip/openlane/l1iinterface/runs/22_09_13_01_32/results/signoff/l1icache_32.magic.gds
string GDS_START 303802
<< end >>

