magic
tech sky130B
magscale 1 2
timestamp 1663004689
<< obsli1 >>
rect 1104 2159 138828 87601
<< obsm1 >>
rect 14 1232 139826 88256
<< metal2 >>
rect 18 89200 74 90000
rect 662 89200 718 90000
rect 1950 89200 2006 90000
rect 2594 89200 2650 90000
rect 3238 89200 3294 90000
rect 4526 89200 4582 90000
rect 5170 89200 5226 90000
rect 5814 89200 5870 90000
rect 7102 89200 7158 90000
rect 7746 89200 7802 90000
rect 8390 89200 8446 90000
rect 9678 89200 9734 90000
rect 10322 89200 10378 90000
rect 10966 89200 11022 90000
rect 12254 89200 12310 90000
rect 12898 89200 12954 90000
rect 13542 89200 13598 90000
rect 14830 89200 14886 90000
rect 15474 89200 15530 90000
rect 16118 89200 16174 90000
rect 17406 89200 17462 90000
rect 18050 89200 18106 90000
rect 19338 89200 19394 90000
rect 19982 89200 20038 90000
rect 20626 89200 20682 90000
rect 21914 89200 21970 90000
rect 22558 89200 22614 90000
rect 23202 89200 23258 90000
rect 24490 89200 24546 90000
rect 25134 89200 25190 90000
rect 25778 89200 25834 90000
rect 27066 89200 27122 90000
rect 27710 89200 27766 90000
rect 28354 89200 28410 90000
rect 29642 89200 29698 90000
rect 30286 89200 30342 90000
rect 30930 89200 30986 90000
rect 32218 89200 32274 90000
rect 32862 89200 32918 90000
rect 33506 89200 33562 90000
rect 34794 89200 34850 90000
rect 35438 89200 35494 90000
rect 36082 89200 36138 90000
rect 37370 89200 37426 90000
rect 38014 89200 38070 90000
rect 39302 89200 39358 90000
rect 39946 89200 40002 90000
rect 40590 89200 40646 90000
rect 41878 89200 41934 90000
rect 42522 89200 42578 90000
rect 43166 89200 43222 90000
rect 44454 89200 44510 90000
rect 45098 89200 45154 90000
rect 45742 89200 45798 90000
rect 47030 89200 47086 90000
rect 47674 89200 47730 90000
rect 48318 89200 48374 90000
rect 49606 89200 49662 90000
rect 50250 89200 50306 90000
rect 50894 89200 50950 90000
rect 52182 89200 52238 90000
rect 52826 89200 52882 90000
rect 53470 89200 53526 90000
rect 54758 89200 54814 90000
rect 55402 89200 55458 90000
rect 56046 89200 56102 90000
rect 57334 89200 57390 90000
rect 57978 89200 58034 90000
rect 59266 89200 59322 90000
rect 59910 89200 59966 90000
rect 60554 89200 60610 90000
rect 61842 89200 61898 90000
rect 62486 89200 62542 90000
rect 63130 89200 63186 90000
rect 64418 89200 64474 90000
rect 65062 89200 65118 90000
rect 65706 89200 65762 90000
rect 66994 89200 67050 90000
rect 67638 89200 67694 90000
rect 68282 89200 68338 90000
rect 69570 89200 69626 90000
rect 70214 89200 70270 90000
rect 70858 89200 70914 90000
rect 72146 89200 72202 90000
rect 72790 89200 72846 90000
rect 73434 89200 73490 90000
rect 74722 89200 74778 90000
rect 75366 89200 75422 90000
rect 76010 89200 76066 90000
rect 77298 89200 77354 90000
rect 77942 89200 77998 90000
rect 79230 89200 79286 90000
rect 79874 89200 79930 90000
rect 80518 89200 80574 90000
rect 81806 89200 81862 90000
rect 82450 89200 82506 90000
rect 83094 89200 83150 90000
rect 84382 89200 84438 90000
rect 85026 89200 85082 90000
rect 85670 89200 85726 90000
rect 86958 89200 87014 90000
rect 87602 89200 87658 90000
rect 88246 89200 88302 90000
rect 89534 89200 89590 90000
rect 90178 89200 90234 90000
rect 90822 89200 90878 90000
rect 92110 89200 92166 90000
rect 92754 89200 92810 90000
rect 93398 89200 93454 90000
rect 94686 89200 94742 90000
rect 95330 89200 95386 90000
rect 95974 89200 96030 90000
rect 97262 89200 97318 90000
rect 97906 89200 97962 90000
rect 98550 89200 98606 90000
rect 99838 89200 99894 90000
rect 100482 89200 100538 90000
rect 101770 89200 101826 90000
rect 102414 89200 102470 90000
rect 103058 89200 103114 90000
rect 104346 89200 104402 90000
rect 104990 89200 105046 90000
rect 105634 89200 105690 90000
rect 106922 89200 106978 90000
rect 107566 89200 107622 90000
rect 108210 89200 108266 90000
rect 109498 89200 109554 90000
rect 110142 89200 110198 90000
rect 110786 89200 110842 90000
rect 112074 89200 112130 90000
rect 112718 89200 112774 90000
rect 113362 89200 113418 90000
rect 114650 89200 114706 90000
rect 115294 89200 115350 90000
rect 115938 89200 115994 90000
rect 117226 89200 117282 90000
rect 117870 89200 117926 90000
rect 118514 89200 118570 90000
rect 119802 89200 119858 90000
rect 120446 89200 120502 90000
rect 121734 89200 121790 90000
rect 122378 89200 122434 90000
rect 123022 89200 123078 90000
rect 124310 89200 124366 90000
rect 124954 89200 125010 90000
rect 125598 89200 125654 90000
rect 126886 89200 126942 90000
rect 127530 89200 127586 90000
rect 128174 89200 128230 90000
rect 129462 89200 129518 90000
rect 130106 89200 130162 90000
rect 130750 89200 130806 90000
rect 132038 89200 132094 90000
rect 132682 89200 132738 90000
rect 133326 89200 133382 90000
rect 134614 89200 134670 90000
rect 135258 89200 135314 90000
rect 135902 89200 135958 90000
rect 137190 89200 137246 90000
rect 137834 89200 137890 90000
rect 138478 89200 138534 90000
rect 139766 89200 139822 90000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92754 0 92810 800
rect 93398 0 93454 800
rect 94042 0 94098 800
rect 95330 0 95386 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 100482 0 100538 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 103058 0 103114 800
rect 103702 0 103758 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106278 0 106334 800
rect 107566 0 107622 800
rect 108210 0 108266 800
rect 108854 0 108910 800
rect 110142 0 110198 800
rect 110786 0 110842 800
rect 111430 0 111486 800
rect 112718 0 112774 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 115294 0 115350 800
rect 115938 0 115994 800
rect 116582 0 116638 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119158 0 119214 800
rect 120446 0 120502 800
rect 121090 0 121146 800
rect 121734 0 121790 800
rect 123022 0 123078 800
rect 123666 0 123722 800
rect 124954 0 125010 800
rect 125598 0 125654 800
rect 126242 0 126298 800
rect 127530 0 127586 800
rect 128174 0 128230 800
rect 128818 0 128874 800
rect 130106 0 130162 800
rect 130750 0 130806 800
rect 131394 0 131450 800
rect 132682 0 132738 800
rect 133326 0 133382 800
rect 133970 0 134026 800
rect 135258 0 135314 800
rect 135902 0 135958 800
rect 136546 0 136602 800
rect 137834 0 137890 800
rect 138478 0 138534 800
rect 139122 0 139178 800
<< obsm2 >>
rect 130 89144 606 89865
rect 774 89144 1894 89865
rect 2062 89144 2538 89865
rect 2706 89144 3182 89865
rect 3350 89144 4470 89865
rect 4638 89144 5114 89865
rect 5282 89144 5758 89865
rect 5926 89144 7046 89865
rect 7214 89144 7690 89865
rect 7858 89144 8334 89865
rect 8502 89144 9622 89865
rect 9790 89144 10266 89865
rect 10434 89144 10910 89865
rect 11078 89144 12198 89865
rect 12366 89144 12842 89865
rect 13010 89144 13486 89865
rect 13654 89144 14774 89865
rect 14942 89144 15418 89865
rect 15586 89144 16062 89865
rect 16230 89144 17350 89865
rect 17518 89144 17994 89865
rect 18162 89144 19282 89865
rect 19450 89144 19926 89865
rect 20094 89144 20570 89865
rect 20738 89144 21858 89865
rect 22026 89144 22502 89865
rect 22670 89144 23146 89865
rect 23314 89144 24434 89865
rect 24602 89144 25078 89865
rect 25246 89144 25722 89865
rect 25890 89144 27010 89865
rect 27178 89144 27654 89865
rect 27822 89144 28298 89865
rect 28466 89144 29586 89865
rect 29754 89144 30230 89865
rect 30398 89144 30874 89865
rect 31042 89144 32162 89865
rect 32330 89144 32806 89865
rect 32974 89144 33450 89865
rect 33618 89144 34738 89865
rect 34906 89144 35382 89865
rect 35550 89144 36026 89865
rect 36194 89144 37314 89865
rect 37482 89144 37958 89865
rect 38126 89144 39246 89865
rect 39414 89144 39890 89865
rect 40058 89144 40534 89865
rect 40702 89144 41822 89865
rect 41990 89144 42466 89865
rect 42634 89144 43110 89865
rect 43278 89144 44398 89865
rect 44566 89144 45042 89865
rect 45210 89144 45686 89865
rect 45854 89144 46974 89865
rect 47142 89144 47618 89865
rect 47786 89144 48262 89865
rect 48430 89144 49550 89865
rect 49718 89144 50194 89865
rect 50362 89144 50838 89865
rect 51006 89144 52126 89865
rect 52294 89144 52770 89865
rect 52938 89144 53414 89865
rect 53582 89144 54702 89865
rect 54870 89144 55346 89865
rect 55514 89144 55990 89865
rect 56158 89144 57278 89865
rect 57446 89144 57922 89865
rect 58090 89144 59210 89865
rect 59378 89144 59854 89865
rect 60022 89144 60498 89865
rect 60666 89144 61786 89865
rect 61954 89144 62430 89865
rect 62598 89144 63074 89865
rect 63242 89144 64362 89865
rect 64530 89144 65006 89865
rect 65174 89144 65650 89865
rect 65818 89144 66938 89865
rect 67106 89144 67582 89865
rect 67750 89144 68226 89865
rect 68394 89144 69514 89865
rect 69682 89144 70158 89865
rect 70326 89144 70802 89865
rect 70970 89144 72090 89865
rect 72258 89144 72734 89865
rect 72902 89144 73378 89865
rect 73546 89144 74666 89865
rect 74834 89144 75310 89865
rect 75478 89144 75954 89865
rect 76122 89144 77242 89865
rect 77410 89144 77886 89865
rect 78054 89144 79174 89865
rect 79342 89144 79818 89865
rect 79986 89144 80462 89865
rect 80630 89144 81750 89865
rect 81918 89144 82394 89865
rect 82562 89144 83038 89865
rect 83206 89144 84326 89865
rect 84494 89144 84970 89865
rect 85138 89144 85614 89865
rect 85782 89144 86902 89865
rect 87070 89144 87546 89865
rect 87714 89144 88190 89865
rect 88358 89144 89478 89865
rect 89646 89144 90122 89865
rect 90290 89144 90766 89865
rect 90934 89144 92054 89865
rect 92222 89144 92698 89865
rect 92866 89144 93342 89865
rect 93510 89144 94630 89865
rect 94798 89144 95274 89865
rect 95442 89144 95918 89865
rect 96086 89144 97206 89865
rect 97374 89144 97850 89865
rect 98018 89144 98494 89865
rect 98662 89144 99782 89865
rect 99950 89144 100426 89865
rect 100594 89144 101714 89865
rect 101882 89144 102358 89865
rect 102526 89144 103002 89865
rect 103170 89144 104290 89865
rect 104458 89144 104934 89865
rect 105102 89144 105578 89865
rect 105746 89144 106866 89865
rect 107034 89144 107510 89865
rect 107678 89144 108154 89865
rect 108322 89144 109442 89865
rect 109610 89144 110086 89865
rect 110254 89144 110730 89865
rect 110898 89144 112018 89865
rect 112186 89144 112662 89865
rect 112830 89144 113306 89865
rect 113474 89144 114594 89865
rect 114762 89144 115238 89865
rect 115406 89144 115882 89865
rect 116050 89144 117170 89865
rect 117338 89144 117814 89865
rect 117982 89144 118458 89865
rect 118626 89144 119746 89865
rect 119914 89144 120390 89865
rect 120558 89144 121678 89865
rect 121846 89144 122322 89865
rect 122490 89144 122966 89865
rect 123134 89144 124254 89865
rect 124422 89144 124898 89865
rect 125066 89144 125542 89865
rect 125710 89144 126830 89865
rect 126998 89144 127474 89865
rect 127642 89144 128118 89865
rect 128286 89144 129406 89865
rect 129574 89144 130050 89865
rect 130218 89144 130694 89865
rect 130862 89144 131982 89865
rect 132150 89144 132626 89865
rect 132794 89144 133270 89865
rect 133438 89144 134558 89865
rect 134726 89144 135202 89865
rect 135370 89144 135846 89865
rect 136014 89144 137134 89865
rect 137302 89144 137778 89865
rect 137946 89144 138422 89865
rect 138590 89144 139710 89865
rect 20 856 139820 89144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 2538 856
rect 2706 31 3182 856
rect 3350 31 3826 856
rect 3994 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7690 856
rect 7858 31 8334 856
rect 8502 31 8978 856
rect 9146 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14130 856
rect 14298 31 15418 856
rect 15586 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19282 856
rect 19450 31 20570 856
rect 20738 31 21214 856
rect 21382 31 22502 856
rect 22670 31 23146 856
rect 23314 31 23790 856
rect 23958 31 25078 856
rect 25246 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27654 856
rect 27822 31 28298 856
rect 28466 31 28942 856
rect 29110 31 30230 856
rect 30398 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34094 856
rect 34262 31 35382 856
rect 35550 31 36026 856
rect 36194 31 36670 856
rect 36838 31 37958 856
rect 38126 31 38602 856
rect 38770 31 39246 856
rect 39414 31 40534 856
rect 40702 31 41178 856
rect 41346 31 42466 856
rect 42634 31 43110 856
rect 43278 31 43754 856
rect 43922 31 45042 856
rect 45210 31 45686 856
rect 45854 31 46330 856
rect 46498 31 47618 856
rect 47786 31 48262 856
rect 48430 31 48906 856
rect 49074 31 50194 856
rect 50362 31 50838 856
rect 51006 31 51482 856
rect 51650 31 52770 856
rect 52938 31 53414 856
rect 53582 31 54058 856
rect 54226 31 55346 856
rect 55514 31 55990 856
rect 56158 31 56634 856
rect 56802 31 57922 856
rect 58090 31 58566 856
rect 58734 31 59210 856
rect 59378 31 60498 856
rect 60666 31 61142 856
rect 61310 31 62430 856
rect 62598 31 63074 856
rect 63242 31 63718 856
rect 63886 31 65006 856
rect 65174 31 65650 856
rect 65818 31 66294 856
rect 66462 31 67582 856
rect 67750 31 68226 856
rect 68394 31 68870 856
rect 69038 31 70158 856
rect 70326 31 70802 856
rect 70970 31 71446 856
rect 71614 31 72734 856
rect 72902 31 73378 856
rect 73546 31 74022 856
rect 74190 31 75310 856
rect 75478 31 75954 856
rect 76122 31 76598 856
rect 76766 31 77886 856
rect 78054 31 78530 856
rect 78698 31 79174 856
rect 79342 31 80462 856
rect 80630 31 81106 856
rect 81274 31 82394 856
rect 82562 31 83038 856
rect 83206 31 83682 856
rect 83850 31 84970 856
rect 85138 31 85614 856
rect 85782 31 86258 856
rect 86426 31 87546 856
rect 87714 31 88190 856
rect 88358 31 88834 856
rect 89002 31 90122 856
rect 90290 31 90766 856
rect 90934 31 91410 856
rect 91578 31 92698 856
rect 92866 31 93342 856
rect 93510 31 93986 856
rect 94154 31 95274 856
rect 95442 31 95918 856
rect 96086 31 96562 856
rect 96730 31 97850 856
rect 98018 31 98494 856
rect 98662 31 99138 856
rect 99306 31 100426 856
rect 100594 31 101070 856
rect 101238 31 101714 856
rect 101882 31 103002 856
rect 103170 31 103646 856
rect 103814 31 104934 856
rect 105102 31 105578 856
rect 105746 31 106222 856
rect 106390 31 107510 856
rect 107678 31 108154 856
rect 108322 31 108798 856
rect 108966 31 110086 856
rect 110254 31 110730 856
rect 110898 31 111374 856
rect 111542 31 112662 856
rect 112830 31 113306 856
rect 113474 31 113950 856
rect 114118 31 115238 856
rect 115406 31 115882 856
rect 116050 31 116526 856
rect 116694 31 117814 856
rect 117982 31 118458 856
rect 118626 31 119102 856
rect 119270 31 120390 856
rect 120558 31 121034 856
rect 121202 31 121678 856
rect 121846 31 122966 856
rect 123134 31 123610 856
rect 123778 31 124898 856
rect 125066 31 125542 856
rect 125710 31 126186 856
rect 126354 31 127474 856
rect 127642 31 128118 856
rect 128286 31 128762 856
rect 128930 31 130050 856
rect 130218 31 130694 856
rect 130862 31 131338 856
rect 131506 31 132626 856
rect 132794 31 133270 856
rect 133438 31 133914 856
rect 134082 31 135202 856
rect 135370 31 135846 856
rect 136014 31 136490 856
rect 136658 31 137778 856
rect 137946 31 138422 856
rect 138590 31 139066 856
rect 139234 31 139820 856
<< metal3 >>
rect 0 89768 800 89888
rect 139200 89768 140000 89888
rect 0 88408 800 88528
rect 139200 88408 140000 88528
rect 0 87728 800 87848
rect 139200 87728 140000 87848
rect 0 87048 800 87168
rect 139200 87048 140000 87168
rect 0 85688 800 85808
rect 139200 85688 140000 85808
rect 0 85008 800 85128
rect 139200 85008 140000 85128
rect 139200 84328 140000 84448
rect 0 83648 800 83768
rect 0 82968 800 83088
rect 139200 82968 140000 83088
rect 0 82288 800 82408
rect 139200 82288 140000 82408
rect 139200 81608 140000 81728
rect 0 80928 800 81048
rect 0 80248 800 80368
rect 139200 80248 140000 80368
rect 0 79568 800 79688
rect 139200 79568 140000 79688
rect 139200 78888 140000 79008
rect 0 78208 800 78328
rect 0 77528 800 77648
rect 139200 77528 140000 77648
rect 0 76848 800 76968
rect 139200 76848 140000 76968
rect 139200 76168 140000 76288
rect 0 75488 800 75608
rect 0 74808 800 74928
rect 139200 74808 140000 74928
rect 0 74128 800 74248
rect 139200 74128 140000 74248
rect 139200 73448 140000 73568
rect 0 72768 800 72888
rect 0 72088 800 72208
rect 139200 72088 140000 72208
rect 0 71408 800 71528
rect 139200 71408 140000 71528
rect 139200 70728 140000 70848
rect 0 70048 800 70168
rect 0 69368 800 69488
rect 139200 69368 140000 69488
rect 0 68688 800 68808
rect 139200 68688 140000 68808
rect 0 67328 800 67448
rect 139200 67328 140000 67448
rect 0 66648 800 66768
rect 139200 66648 140000 66768
rect 0 65968 800 66088
rect 139200 65968 140000 66088
rect 0 64608 800 64728
rect 139200 64608 140000 64728
rect 0 63928 800 64048
rect 139200 63928 140000 64048
rect 139200 63248 140000 63368
rect 0 62568 800 62688
rect 0 61888 800 62008
rect 139200 61888 140000 62008
rect 0 61208 800 61328
rect 139200 61208 140000 61328
rect 139200 60528 140000 60648
rect 0 59848 800 59968
rect 0 59168 800 59288
rect 139200 59168 140000 59288
rect 0 58488 800 58608
rect 139200 58488 140000 58608
rect 139200 57808 140000 57928
rect 0 57128 800 57248
rect 0 56448 800 56568
rect 139200 56448 140000 56568
rect 0 55768 800 55888
rect 139200 55768 140000 55888
rect 139200 55088 140000 55208
rect 0 54408 800 54528
rect 0 53728 800 53848
rect 139200 53728 140000 53848
rect 0 53048 800 53168
rect 139200 53048 140000 53168
rect 139200 52368 140000 52488
rect 0 51688 800 51808
rect 0 51008 800 51128
rect 139200 51008 140000 51128
rect 0 50328 800 50448
rect 139200 50328 140000 50448
rect 139200 49648 140000 49768
rect 0 48968 800 49088
rect 0 48288 800 48408
rect 139200 48288 140000 48408
rect 0 47608 800 47728
rect 139200 47608 140000 47728
rect 0 46248 800 46368
rect 139200 46248 140000 46368
rect 0 45568 800 45688
rect 139200 45568 140000 45688
rect 0 44888 800 45008
rect 139200 44888 140000 45008
rect 0 43528 800 43648
rect 139200 43528 140000 43648
rect 0 42848 800 42968
rect 139200 42848 140000 42968
rect 139200 42168 140000 42288
rect 0 41488 800 41608
rect 0 40808 800 40928
rect 139200 40808 140000 40928
rect 0 40128 800 40248
rect 139200 40128 140000 40248
rect 139200 39448 140000 39568
rect 0 38768 800 38888
rect 0 38088 800 38208
rect 139200 38088 140000 38208
rect 0 37408 800 37528
rect 139200 37408 140000 37528
rect 139200 36728 140000 36848
rect 0 36048 800 36168
rect 0 35368 800 35488
rect 139200 35368 140000 35488
rect 0 34688 800 34808
rect 139200 34688 140000 34808
rect 139200 34008 140000 34128
rect 0 33328 800 33448
rect 0 32648 800 32768
rect 139200 32648 140000 32768
rect 0 31968 800 32088
rect 139200 31968 140000 32088
rect 139200 31288 140000 31408
rect 0 30608 800 30728
rect 0 29928 800 30048
rect 139200 29928 140000 30048
rect 0 29248 800 29368
rect 139200 29248 140000 29368
rect 139200 28568 140000 28688
rect 0 27888 800 28008
rect 0 27208 800 27328
rect 139200 27208 140000 27328
rect 0 26528 800 26648
rect 139200 26528 140000 26648
rect 139200 25848 140000 25968
rect 0 25168 800 25288
rect 0 24488 800 24608
rect 139200 24488 140000 24608
rect 0 23808 800 23928
rect 139200 23808 140000 23928
rect 0 22448 800 22568
rect 139200 22448 140000 22568
rect 0 21768 800 21888
rect 139200 21768 140000 21888
rect 139200 21088 140000 21208
rect 0 20408 800 20528
rect 0 19728 800 19848
rect 139200 19728 140000 19848
rect 0 19048 800 19168
rect 139200 19048 140000 19168
rect 139200 18368 140000 18488
rect 0 17688 800 17808
rect 0 17008 800 17128
rect 139200 17008 140000 17128
rect 0 16328 800 16448
rect 139200 16328 140000 16448
rect 139200 15648 140000 15768
rect 0 14968 800 15088
rect 0 14288 800 14408
rect 139200 14288 140000 14408
rect 0 13608 800 13728
rect 139200 13608 140000 13728
rect 139200 12928 140000 13048
rect 0 12248 800 12368
rect 0 11568 800 11688
rect 139200 11568 140000 11688
rect 0 10888 800 11008
rect 139200 10888 140000 11008
rect 139200 10208 140000 10328
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 139200 8848 140000 8968
rect 0 8168 800 8288
rect 139200 8168 140000 8288
rect 139200 7488 140000 7608
rect 0 6808 800 6928
rect 0 6128 800 6248
rect 139200 6128 140000 6248
rect 0 5448 800 5568
rect 139200 5448 140000 5568
rect 139200 4768 140000 4888
rect 0 4088 800 4208
rect 0 3408 800 3528
rect 139200 3408 140000 3528
rect 0 2728 800 2848
rect 139200 2728 140000 2848
rect 0 1368 800 1488
rect 139200 1368 140000 1488
rect 0 688 800 808
rect 139200 688 140000 808
rect 139200 8 140000 128
<< obsm3 >>
rect 880 89688 139120 89861
rect 800 88608 139200 89688
rect 880 88328 139120 88608
rect 800 87928 139200 88328
rect 880 87648 139120 87928
rect 800 87248 139200 87648
rect 880 86968 139120 87248
rect 800 85888 139200 86968
rect 880 85608 139120 85888
rect 800 85208 139200 85608
rect 880 84928 139120 85208
rect 800 84528 139200 84928
rect 800 84248 139120 84528
rect 800 83848 139200 84248
rect 880 83568 139200 83848
rect 800 83168 139200 83568
rect 880 82888 139120 83168
rect 800 82488 139200 82888
rect 880 82208 139120 82488
rect 800 81808 139200 82208
rect 800 81528 139120 81808
rect 800 81128 139200 81528
rect 880 80848 139200 81128
rect 800 80448 139200 80848
rect 880 80168 139120 80448
rect 800 79768 139200 80168
rect 880 79488 139120 79768
rect 800 79088 139200 79488
rect 800 78808 139120 79088
rect 800 78408 139200 78808
rect 880 78128 139200 78408
rect 800 77728 139200 78128
rect 880 77448 139120 77728
rect 800 77048 139200 77448
rect 880 76768 139120 77048
rect 800 76368 139200 76768
rect 800 76088 139120 76368
rect 800 75688 139200 76088
rect 880 75408 139200 75688
rect 800 75008 139200 75408
rect 880 74728 139120 75008
rect 800 74328 139200 74728
rect 880 74048 139120 74328
rect 800 73648 139200 74048
rect 800 73368 139120 73648
rect 800 72968 139200 73368
rect 880 72688 139200 72968
rect 800 72288 139200 72688
rect 880 72008 139120 72288
rect 800 71608 139200 72008
rect 880 71328 139120 71608
rect 800 70928 139200 71328
rect 800 70648 139120 70928
rect 800 70248 139200 70648
rect 880 69968 139200 70248
rect 800 69568 139200 69968
rect 880 69288 139120 69568
rect 800 68888 139200 69288
rect 880 68608 139120 68888
rect 800 67528 139200 68608
rect 880 67248 139120 67528
rect 800 66848 139200 67248
rect 880 66568 139120 66848
rect 800 66168 139200 66568
rect 880 65888 139120 66168
rect 800 64808 139200 65888
rect 880 64528 139120 64808
rect 800 64128 139200 64528
rect 880 63848 139120 64128
rect 800 63448 139200 63848
rect 800 63168 139120 63448
rect 800 62768 139200 63168
rect 880 62488 139200 62768
rect 800 62088 139200 62488
rect 880 61808 139120 62088
rect 800 61408 139200 61808
rect 880 61128 139120 61408
rect 800 60728 139200 61128
rect 800 60448 139120 60728
rect 800 60048 139200 60448
rect 880 59768 139200 60048
rect 800 59368 139200 59768
rect 880 59088 139120 59368
rect 800 58688 139200 59088
rect 880 58408 139120 58688
rect 800 58008 139200 58408
rect 800 57728 139120 58008
rect 800 57328 139200 57728
rect 880 57048 139200 57328
rect 800 56648 139200 57048
rect 880 56368 139120 56648
rect 800 55968 139200 56368
rect 880 55688 139120 55968
rect 800 55288 139200 55688
rect 800 55008 139120 55288
rect 800 54608 139200 55008
rect 880 54328 139200 54608
rect 800 53928 139200 54328
rect 880 53648 139120 53928
rect 800 53248 139200 53648
rect 880 52968 139120 53248
rect 800 52568 139200 52968
rect 800 52288 139120 52568
rect 800 51888 139200 52288
rect 880 51608 139200 51888
rect 800 51208 139200 51608
rect 880 50928 139120 51208
rect 800 50528 139200 50928
rect 880 50248 139120 50528
rect 800 49848 139200 50248
rect 800 49568 139120 49848
rect 800 49168 139200 49568
rect 880 48888 139200 49168
rect 800 48488 139200 48888
rect 880 48208 139120 48488
rect 800 47808 139200 48208
rect 880 47528 139120 47808
rect 800 46448 139200 47528
rect 880 46168 139120 46448
rect 800 45768 139200 46168
rect 880 45488 139120 45768
rect 800 45088 139200 45488
rect 880 44808 139120 45088
rect 800 43728 139200 44808
rect 880 43448 139120 43728
rect 800 43048 139200 43448
rect 880 42768 139120 43048
rect 800 42368 139200 42768
rect 800 42088 139120 42368
rect 800 41688 139200 42088
rect 880 41408 139200 41688
rect 800 41008 139200 41408
rect 880 40728 139120 41008
rect 800 40328 139200 40728
rect 880 40048 139120 40328
rect 800 39648 139200 40048
rect 800 39368 139120 39648
rect 800 38968 139200 39368
rect 880 38688 139200 38968
rect 800 38288 139200 38688
rect 880 38008 139120 38288
rect 800 37608 139200 38008
rect 880 37328 139120 37608
rect 800 36928 139200 37328
rect 800 36648 139120 36928
rect 800 36248 139200 36648
rect 880 35968 139200 36248
rect 800 35568 139200 35968
rect 880 35288 139120 35568
rect 800 34888 139200 35288
rect 880 34608 139120 34888
rect 800 34208 139200 34608
rect 800 33928 139120 34208
rect 800 33528 139200 33928
rect 880 33248 139200 33528
rect 800 32848 139200 33248
rect 880 32568 139120 32848
rect 800 32168 139200 32568
rect 880 31888 139120 32168
rect 800 31488 139200 31888
rect 800 31208 139120 31488
rect 800 30808 139200 31208
rect 880 30528 139200 30808
rect 800 30128 139200 30528
rect 880 29848 139120 30128
rect 800 29448 139200 29848
rect 880 29168 139120 29448
rect 800 28768 139200 29168
rect 800 28488 139120 28768
rect 800 28088 139200 28488
rect 880 27808 139200 28088
rect 800 27408 139200 27808
rect 880 27128 139120 27408
rect 800 26728 139200 27128
rect 880 26448 139120 26728
rect 800 26048 139200 26448
rect 800 25768 139120 26048
rect 800 25368 139200 25768
rect 880 25088 139200 25368
rect 800 24688 139200 25088
rect 880 24408 139120 24688
rect 800 24008 139200 24408
rect 880 23728 139120 24008
rect 800 22648 139200 23728
rect 880 22368 139120 22648
rect 800 21968 139200 22368
rect 880 21688 139120 21968
rect 800 21288 139200 21688
rect 800 21008 139120 21288
rect 800 20608 139200 21008
rect 880 20328 139200 20608
rect 800 19928 139200 20328
rect 880 19648 139120 19928
rect 800 19248 139200 19648
rect 880 18968 139120 19248
rect 800 18568 139200 18968
rect 800 18288 139120 18568
rect 800 17888 139200 18288
rect 880 17608 139200 17888
rect 800 17208 139200 17608
rect 880 16928 139120 17208
rect 800 16528 139200 16928
rect 880 16248 139120 16528
rect 800 15848 139200 16248
rect 800 15568 139120 15848
rect 800 15168 139200 15568
rect 880 14888 139200 15168
rect 800 14488 139200 14888
rect 880 14208 139120 14488
rect 800 13808 139200 14208
rect 880 13528 139120 13808
rect 800 13128 139200 13528
rect 800 12848 139120 13128
rect 800 12448 139200 12848
rect 880 12168 139200 12448
rect 800 11768 139200 12168
rect 880 11488 139120 11768
rect 800 11088 139200 11488
rect 880 10808 139120 11088
rect 800 10408 139200 10808
rect 800 10128 139120 10408
rect 800 9728 139200 10128
rect 880 9448 139200 9728
rect 800 9048 139200 9448
rect 880 8768 139120 9048
rect 800 8368 139200 8768
rect 880 8088 139120 8368
rect 800 7688 139200 8088
rect 800 7408 139120 7688
rect 800 7008 139200 7408
rect 880 6728 139200 7008
rect 800 6328 139200 6728
rect 880 6048 139120 6328
rect 800 5648 139200 6048
rect 880 5368 139120 5648
rect 800 4968 139200 5368
rect 800 4688 139120 4968
rect 800 4288 139200 4688
rect 880 4008 139200 4288
rect 800 3608 139200 4008
rect 880 3328 139120 3608
rect 800 2928 139200 3328
rect 880 2648 139120 2928
rect 800 1568 139200 2648
rect 880 1288 139120 1568
rect 800 888 139200 1288
rect 880 608 139120 888
rect 800 208 139200 608
rect 800 35 139120 208
<< metal4 >>
rect 4208 2128 4528 87632
rect 19568 2128 19888 87632
rect 34928 2128 35248 87632
rect 50288 2128 50608 87632
rect 65648 2128 65968 87632
rect 81008 2128 81328 87632
rect 96368 2128 96688 87632
rect 111728 2128 112048 87632
rect 127088 2128 127408 87632
<< obsm4 >>
rect 18827 2347 19488 86189
rect 19968 2347 34848 86189
rect 35328 2347 50208 86189
rect 50688 2347 65568 86189
rect 66048 2347 80928 86189
rect 81408 2347 96288 86189
rect 96768 2347 111648 86189
rect 112128 2347 115861 86189
<< labels >>
rlabel metal2 s 126242 0 126298 800 6 clk
port 1 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 data_chip_en_1
port 2 nsew signal output
rlabel metal3 s 0 688 800 808 6 data_chip_en_2
port 3 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 data_in_1[0]
port 4 nsew signal output
rlabel metal2 s 70214 89200 70270 90000 6 data_in_1[10]
port 5 nsew signal output
rlabel metal2 s 40590 89200 40646 90000 6 data_in_1[11]
port 6 nsew signal output
rlabel metal3 s 139200 43528 140000 43648 6 data_in_1[12]
port 7 nsew signal output
rlabel metal2 s 69570 89200 69626 90000 6 data_in_1[13]
port 8 nsew signal output
rlabel metal3 s 139200 61888 140000 62008 6 data_in_1[14]
port 9 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 data_in_1[15]
port 10 nsew signal output
rlabel metal2 s 8390 89200 8446 90000 6 data_in_1[16]
port 11 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 data_in_1[17]
port 12 nsew signal output
rlabel metal3 s 139200 87048 140000 87168 6 data_in_1[18]
port 13 nsew signal output
rlabel metal3 s 139200 35368 140000 35488 6 data_in_1[19]
port 14 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 data_in_1[1]
port 15 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 data_in_1[20]
port 16 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 data_in_1[21]
port 17 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 data_in_1[22]
port 18 nsew signal output
rlabel metal3 s 139200 52368 140000 52488 6 data_in_1[23]
port 19 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 data_in_1[24]
port 20 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 data_in_1[25]
port 21 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 data_in_1[26]
port 22 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 data_in_1[27]
port 23 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 data_in_1[28]
port 24 nsew signal output
rlabel metal2 s 90178 89200 90234 90000 6 data_in_1[29]
port 25 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 data_in_1[2]
port 26 nsew signal output
rlabel metal2 s 135258 89200 135314 90000 6 data_in_1[30]
port 27 nsew signal output
rlabel metal2 s 105634 89200 105690 90000 6 data_in_1[31]
port 28 nsew signal output
rlabel metal3 s 139200 11568 140000 11688 6 data_in_1[3]
port 29 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 data_in_1[4]
port 30 nsew signal output
rlabel metal2 s 109498 89200 109554 90000 6 data_in_1[5]
port 31 nsew signal output
rlabel metal2 s 77942 89200 77998 90000 6 data_in_1[6]
port 32 nsew signal output
rlabel metal3 s 139200 31968 140000 32088 6 data_in_1[7]
port 33 nsew signal output
rlabel metal2 s 10966 89200 11022 90000 6 data_in_1[8]
port 34 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 data_in_1[9]
port 35 nsew signal output
rlabel metal2 s 108210 89200 108266 90000 6 data_in_2[0]
port 36 nsew signal output
rlabel metal3 s 139200 19048 140000 19168 6 data_in_2[10]
port 37 nsew signal output
rlabel metal2 s 94686 89200 94742 90000 6 data_in_2[11]
port 38 nsew signal output
rlabel metal2 s 19338 89200 19394 90000 6 data_in_2[12]
port 39 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 data_in_2[13]
port 40 nsew signal output
rlabel metal3 s 139200 36728 140000 36848 6 data_in_2[14]
port 41 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 data_in_2[15]
port 42 nsew signal output
rlabel metal2 s 92754 89200 92810 90000 6 data_in_2[16]
port 43 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 data_in_2[17]
port 44 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 data_in_2[18]
port 45 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 data_in_2[19]
port 46 nsew signal output
rlabel metal2 s 45098 89200 45154 90000 6 data_in_2[1]
port 47 nsew signal output
rlabel metal2 s 93398 89200 93454 90000 6 data_in_2[20]
port 48 nsew signal output
rlabel metal2 s 9678 89200 9734 90000 6 data_in_2[21]
port 49 nsew signal output
rlabel metal2 s 13542 89200 13598 90000 6 data_in_2[22]
port 50 nsew signal output
rlabel metal2 s 2594 89200 2650 90000 6 data_in_2[23]
port 51 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 data_in_2[24]
port 52 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 data_in_2[25]
port 53 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 data_in_2[26]
port 54 nsew signal output
rlabel metal2 s 129462 89200 129518 90000 6 data_in_2[27]
port 55 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 data_in_2[28]
port 56 nsew signal output
rlabel metal3 s 139200 8848 140000 8968 6 data_in_2[29]
port 57 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 data_in_2[2]
port 58 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 data_in_2[30]
port 59 nsew signal output
rlabel metal2 s 130750 89200 130806 90000 6 data_in_2[31]
port 60 nsew signal output
rlabel metal2 s 37370 89200 37426 90000 6 data_in_2[3]
port 61 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 data_in_2[4]
port 62 nsew signal output
rlabel metal2 s 121734 89200 121790 90000 6 data_in_2[5]
port 63 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 data_in_2[6]
port 64 nsew signal output
rlabel metal3 s 139200 87728 140000 87848 6 data_in_2[7]
port 65 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 data_in_2[8]
port 66 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 data_in_2[9]
port 67 nsew signal output
rlabel metal3 s 139200 57808 140000 57928 6 data_index_1[0]
port 68 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 data_index_1[1]
port 69 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 data_index_1[2]
port 70 nsew signal output
rlabel metal3 s 139200 27208 140000 27328 6 data_index_1[3]
port 71 nsew signal output
rlabel metal2 s 61842 89200 61898 90000 6 data_index_1[4]
port 72 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 data_index_1[5]
port 73 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 data_index_1[6]
port 74 nsew signal output
rlabel metal2 s 48318 89200 48374 90000 6 data_index_1[7]
port 75 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 data_index_2[0]
port 76 nsew signal output
rlabel metal2 s 110142 89200 110198 90000 6 data_index_2[1]
port 77 nsew signal output
rlabel metal3 s 139200 81608 140000 81728 6 data_index_2[2]
port 78 nsew signal output
rlabel metal3 s 139200 74808 140000 74928 6 data_index_2[3]
port 79 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 data_index_2[4]
port 80 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 data_index_2[5]
port 81 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 data_index_2[6]
port 82 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 data_index_2[7]
port 83 nsew signal output
rlabel metal3 s 139200 59168 140000 59288 6 data_out_1[0]
port 84 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 data_out_1[10]
port 85 nsew signal input
rlabel metal3 s 139200 32648 140000 32768 6 data_out_1[11]
port 86 nsew signal input
rlabel metal2 s 99838 89200 99894 90000 6 data_out_1[12]
port 87 nsew signal input
rlabel metal3 s 139200 74128 140000 74248 6 data_out_1[13]
port 88 nsew signal input
rlabel metal3 s 139200 24488 140000 24608 6 data_out_1[14]
port 89 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 data_out_1[15]
port 90 nsew signal input
rlabel metal3 s 139200 34008 140000 34128 6 data_out_1[16]
port 91 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 data_out_1[17]
port 92 nsew signal input
rlabel metal3 s 139200 4768 140000 4888 6 data_out_1[18]
port 93 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 data_out_1[19]
port 94 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 data_out_1[1]
port 95 nsew signal input
rlabel metal2 s 104990 89200 105046 90000 6 data_out_1[20]
port 96 nsew signal input
rlabel metal2 s 32218 89200 32274 90000 6 data_out_1[21]
port 97 nsew signal input
rlabel metal2 s 43166 89200 43222 90000 6 data_out_1[22]
port 98 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 data_out_1[23]
port 99 nsew signal input
rlabel metal3 s 139200 38088 140000 38208 6 data_out_1[24]
port 100 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 data_out_1[25]
port 101 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 data_out_1[26]
port 102 nsew signal input
rlabel metal2 s 81806 89200 81862 90000 6 data_out_1[27]
port 103 nsew signal input
rlabel metal3 s 139200 7488 140000 7608 6 data_out_1[28]
port 104 nsew signal input
rlabel metal2 s 132682 89200 132738 90000 6 data_out_1[29]
port 105 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 data_out_1[2]
port 106 nsew signal input
rlabel metal3 s 139200 65968 140000 66088 6 data_out_1[30]
port 107 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 data_out_1[31]
port 108 nsew signal input
rlabel metal3 s 139200 56448 140000 56568 6 data_out_1[3]
port 109 nsew signal input
rlabel metal2 s 70858 89200 70914 90000 6 data_out_1[4]
port 110 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 data_out_1[5]
port 111 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 data_out_1[6]
port 112 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 data_out_1[7]
port 113 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 data_out_1[8]
port 114 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 data_out_1[9]
port 115 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 data_out_2[0]
port 116 nsew signal input
rlabel metal2 s 68282 89200 68338 90000 6 data_out_2[10]
port 117 nsew signal input
rlabel metal3 s 139200 77528 140000 77648 6 data_out_2[11]
port 118 nsew signal input
rlabel metal2 s 88246 89200 88302 90000 6 data_out_2[12]
port 119 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 data_out_2[13]
port 120 nsew signal input
rlabel metal2 s 49606 89200 49662 90000 6 data_out_2[14]
port 121 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 data_out_2[15]
port 122 nsew signal input
rlabel metal2 s 97906 89200 97962 90000 6 data_out_2[16]
port 123 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 data_out_2[17]
port 124 nsew signal input
rlabel metal2 s 34794 89200 34850 90000 6 data_out_2[18]
port 125 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 data_out_2[19]
port 126 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 data_out_2[1]
port 127 nsew signal input
rlabel metal3 s 139200 18368 140000 18488 6 data_out_2[20]
port 128 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 data_out_2[21]
port 129 nsew signal input
rlabel metal2 s 122378 89200 122434 90000 6 data_out_2[22]
port 130 nsew signal input
rlabel metal2 s 115294 89200 115350 90000 6 data_out_2[23]
port 131 nsew signal input
rlabel metal2 s 84382 89200 84438 90000 6 data_out_2[24]
port 132 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 data_out_2[25]
port 133 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 data_out_2[26]
port 134 nsew signal input
rlabel metal2 s 5170 89200 5226 90000 6 data_out_2[27]
port 135 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 data_out_2[28]
port 136 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 data_out_2[29]
port 137 nsew signal input
rlabel metal2 s 30930 89200 30986 90000 6 data_out_2[2]
port 138 nsew signal input
rlabel metal3 s 139200 31288 140000 31408 6 data_out_2[30]
port 139 nsew signal input
rlabel metal2 s 5814 89200 5870 90000 6 data_out_2[31]
port 140 nsew signal input
rlabel metal2 s 22558 89200 22614 90000 6 data_out_2[3]
port 141 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 data_out_2[4]
port 142 nsew signal input
rlabel metal2 s 90822 89200 90878 90000 6 data_out_2[5]
port 143 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 data_out_2[6]
port 144 nsew signal input
rlabel metal2 s 65062 89200 65118 90000 6 data_out_2[7]
port 145 nsew signal input
rlabel metal2 s 10322 89200 10378 90000 6 data_out_2[8]
port 146 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 data_out_2[9]
port 147 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 data_write_en_1
port 148 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 data_write_en_2
port 149 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 ld_data_o[0]
port 150 nsew signal output
rlabel metal3 s 139200 76168 140000 76288 6 ld_data_o[10]
port 151 nsew signal output
rlabel metal3 s 139200 21768 140000 21888 6 ld_data_o[11]
port 152 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 ld_data_o[12]
port 153 nsew signal output
rlabel metal2 s 28354 89200 28410 90000 6 ld_data_o[13]
port 154 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 ld_data_o[14]
port 155 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 ld_data_o[15]
port 156 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 ld_data_o[16]
port 157 nsew signal output
rlabel metal2 s 57978 89200 58034 90000 6 ld_data_o[17]
port 158 nsew signal output
rlabel metal2 s 15474 89200 15530 90000 6 ld_data_o[18]
port 159 nsew signal output
rlabel metal2 s 14830 89200 14886 90000 6 ld_data_o[19]
port 160 nsew signal output
rlabel metal3 s 139200 79568 140000 79688 6 ld_data_o[1]
port 161 nsew signal output
rlabel metal2 s 60554 89200 60610 90000 6 ld_data_o[20]
port 162 nsew signal output
rlabel metal2 s 59266 89200 59322 90000 6 ld_data_o[21]
port 163 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 ld_data_o[22]
port 164 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 ld_data_o[23]
port 165 nsew signal output
rlabel metal2 s 52826 89200 52882 90000 6 ld_data_o[24]
port 166 nsew signal output
rlabel metal2 s 87602 89200 87658 90000 6 ld_data_o[25]
port 167 nsew signal output
rlabel metal2 s 115938 89200 115994 90000 6 ld_data_o[26]
port 168 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 ld_data_o[27]
port 169 nsew signal output
rlabel metal3 s 139200 25848 140000 25968 6 ld_data_o[28]
port 170 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 ld_data_o[29]
port 171 nsew signal output
rlabel metal3 s 139200 40808 140000 40928 6 ld_data_o[2]
port 172 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 ld_data_o[30]
port 173 nsew signal output
rlabel metal2 s 76010 89200 76066 90000 6 ld_data_o[31]
port 174 nsew signal output
rlabel metal3 s 139200 15648 140000 15768 6 ld_data_o[32]
port 175 nsew signal output
rlabel metal2 s 85670 89200 85726 90000 6 ld_data_o[33]
port 176 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 ld_data_o[34]
port 177 nsew signal output
rlabel metal3 s 139200 88408 140000 88528 6 ld_data_o[35]
port 178 nsew signal output
rlabel metal2 s 39946 89200 40002 90000 6 ld_data_o[36]
port 179 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 ld_data_o[37]
port 180 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 ld_data_o[38]
port 181 nsew signal output
rlabel metal3 s 139200 70728 140000 70848 6 ld_data_o[39]
port 182 nsew signal output
rlabel metal3 s 139200 89768 140000 89888 6 ld_data_o[3]
port 183 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 ld_data_o[40]
port 184 nsew signal output
rlabel metal2 s 55402 89200 55458 90000 6 ld_data_o[41]
port 185 nsew signal output
rlabel metal3 s 139200 78888 140000 79008 6 ld_data_o[42]
port 186 nsew signal output
rlabel metal2 s 82450 89200 82506 90000 6 ld_data_o[43]
port 187 nsew signal output
rlabel metal3 s 139200 46248 140000 46368 6 ld_data_o[44]
port 188 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 ld_data_o[45]
port 189 nsew signal output
rlabel metal2 s 32862 89200 32918 90000 6 ld_data_o[46]
port 190 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 ld_data_o[47]
port 191 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 ld_data_o[48]
port 192 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 ld_data_o[49]
port 193 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 ld_data_o[4]
port 194 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 ld_data_o[50]
port 195 nsew signal output
rlabel metal2 s 77298 89200 77354 90000 6 ld_data_o[51]
port 196 nsew signal output
rlabel metal2 s 27710 89200 27766 90000 6 ld_data_o[52]
port 197 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 ld_data_o[53]
port 198 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 ld_data_o[54]
port 199 nsew signal output
rlabel metal2 s 134614 89200 134670 90000 6 ld_data_o[55]
port 200 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 ld_data_o[56]
port 201 nsew signal output
rlabel metal3 s 139200 8 140000 128 6 ld_data_o[57]
port 202 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 ld_data_o[58]
port 203 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 ld_data_o[59]
port 204 nsew signal output
rlabel metal2 s 19982 89200 20038 90000 6 ld_data_o[5]
port 205 nsew signal output
rlabel metal2 s 65706 89200 65762 90000 6 ld_data_o[60]
port 206 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 ld_data_o[61]
port 207 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 ld_data_o[62]
port 208 nsew signal output
rlabel metal2 s 24490 89200 24546 90000 6 ld_data_o[63]
port 209 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 ld_data_o[6]
port 210 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 ld_data_o[7]
port 211 nsew signal output
rlabel metal2 s 75366 89200 75422 90000 6 ld_data_o[8]
port 212 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 ld_data_o[9]
port 213 nsew signal output
rlabel metal2 s 66994 89200 67050 90000 6 opcode
port 214 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 req_addr_i[0]
port 215 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 req_addr_i[10]
port 216 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 req_addr_i[11]
port 217 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 req_addr_i[12]
port 218 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 req_addr_i[13]
port 219 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 req_addr_i[14]
port 220 nsew signal input
rlabel metal3 s 139200 34688 140000 34808 6 req_addr_i[15]
port 221 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 req_addr_i[16]
port 222 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 req_addr_i[17]
port 223 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 req_addr_i[18]
port 224 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 req_addr_i[19]
port 225 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 req_addr_i[1]
port 226 nsew signal input
rlabel metal2 s 62486 89200 62542 90000 6 req_addr_i[20]
port 227 nsew signal input
rlabel metal2 s 47674 89200 47730 90000 6 req_addr_i[21]
port 228 nsew signal input
rlabel metal2 s 139766 89200 139822 90000 6 req_addr_i[22]
port 229 nsew signal input
rlabel metal2 s 72790 89200 72846 90000 6 req_addr_i[23]
port 230 nsew signal input
rlabel metal2 s 3238 89200 3294 90000 6 req_addr_i[24]
port 231 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 req_addr_i[25]
port 232 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 req_addr_i[26]
port 233 nsew signal input
rlabel metal2 s 124310 89200 124366 90000 6 req_addr_i[27]
port 234 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 req_addr_i[28]
port 235 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 req_addr_i[29]
port 236 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 req_addr_i[2]
port 237 nsew signal input
rlabel metal3 s 139200 2728 140000 2848 6 req_addr_i[30]
port 238 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 req_addr_i[31]
port 239 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 req_addr_i[3]
port 240 nsew signal input
rlabel metal2 s 67638 89200 67694 90000 6 req_addr_i[4]
port 241 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 req_addr_i[5]
port 242 nsew signal input
rlabel metal2 s 50894 89200 50950 90000 6 req_addr_i[6]
port 243 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 req_addr_i[7]
port 244 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 req_addr_i[8]
port 245 nsew signal input
rlabel metal2 s 125598 89200 125654 90000 6 req_addr_i[9]
port 246 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 req_ready_o
port 247 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 req_valid_i
port 248 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 resp_ready_i
port 249 nsew signal input
rlabel metal2 s 16118 89200 16174 90000 6 resp_valid_o
port 250 nsew signal output
rlabel metal2 s 135902 89200 135958 90000 6 rob_index_i
port 251 nsew signal input
rlabel metal2 s 52182 89200 52238 90000 6 rob_index_o
port 252 nsew signal output
rlabel metal2 s 25134 89200 25190 90000 6 rstn
port 253 nsew signal input
rlabel metal2 s 130106 89200 130162 90000 6 st_data_i[0]
port 254 nsew signal input
rlabel metal2 s 112074 89200 112130 90000 6 st_data_i[10]
port 255 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 st_data_i[11]
port 256 nsew signal input
rlabel metal2 s 128174 89200 128230 90000 6 st_data_i[12]
port 257 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 st_data_i[13]
port 258 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 st_data_i[14]
port 259 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 st_data_i[15]
port 260 nsew signal input
rlabel metal2 s 20626 89200 20682 90000 6 st_data_i[16]
port 261 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 st_data_i[17]
port 262 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 st_data_i[18]
port 263 nsew signal input
rlabel metal2 s 53470 89200 53526 90000 6 st_data_i[19]
port 264 nsew signal input
rlabel metal2 s 662 0 718 800 6 st_data_i[1]
port 265 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 st_data_i[20]
port 266 nsew signal input
rlabel metal3 s 139200 61208 140000 61328 6 st_data_i[21]
port 267 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 st_data_i[22]
port 268 nsew signal input
rlabel metal3 s 139200 53048 140000 53168 6 st_data_i[23]
port 269 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 st_data_i[24]
port 270 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 st_data_i[25]
port 271 nsew signal input
rlabel metal3 s 139200 12928 140000 13048 6 st_data_i[26]
port 272 nsew signal input
rlabel metal2 s 117226 89200 117282 90000 6 st_data_i[27]
port 273 nsew signal input
rlabel metal2 s 42522 89200 42578 90000 6 st_data_i[28]
port 274 nsew signal input
rlabel metal2 s 113362 89200 113418 90000 6 st_data_i[29]
port 275 nsew signal input
rlabel metal2 s 124954 89200 125010 90000 6 st_data_i[2]
port 276 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 st_data_i[30]
port 277 nsew signal input
rlabel metal2 s 92110 89200 92166 90000 6 st_data_i[31]
port 278 nsew signal input
rlabel metal2 s 120446 89200 120502 90000 6 st_data_i[32]
port 279 nsew signal input
rlabel metal2 s 86958 89200 87014 90000 6 st_data_i[33]
port 280 nsew signal input
rlabel metal3 s 139200 58488 140000 58608 6 st_data_i[34]
port 281 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 st_data_i[35]
port 282 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 st_data_i[36]
port 283 nsew signal input
rlabel metal3 s 139200 80248 140000 80368 6 st_data_i[37]
port 284 nsew signal input
rlabel metal2 s 64418 89200 64474 90000 6 st_data_i[38]
port 285 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 st_data_i[39]
port 286 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 st_data_i[3]
port 287 nsew signal input
rlabel metal2 s 41878 89200 41934 90000 6 st_data_i[40]
port 288 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 st_data_i[41]
port 289 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 st_data_i[42]
port 290 nsew signal input
rlabel metal3 s 139200 82968 140000 83088 6 st_data_i[43]
port 291 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 st_data_i[44]
port 292 nsew signal input
rlabel metal3 s 139200 21088 140000 21208 6 st_data_i[45]
port 293 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 st_data_i[46]
port 294 nsew signal input
rlabel metal3 s 139200 69368 140000 69488 6 st_data_i[47]
port 295 nsew signal input
rlabel metal3 s 139200 19728 140000 19848 6 st_data_i[48]
port 296 nsew signal input
rlabel metal2 s 126886 89200 126942 90000 6 st_data_i[49]
port 297 nsew signal input
rlabel metal2 s 138478 89200 138534 90000 6 st_data_i[4]
port 298 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 st_data_i[50]
port 299 nsew signal input
rlabel metal3 s 139200 42168 140000 42288 6 st_data_i[51]
port 300 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 st_data_i[52]
port 301 nsew signal input
rlabel metal3 s 139200 16328 140000 16448 6 st_data_i[53]
port 302 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 st_data_i[54]
port 303 nsew signal input
rlabel metal2 s 89534 89200 89590 90000 6 st_data_i[55]
port 304 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 st_data_i[56]
port 305 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 st_data_i[57]
port 306 nsew signal input
rlabel metal3 s 139200 63248 140000 63368 6 st_data_i[58]
port 307 nsew signal input
rlabel metal3 s 139200 3408 140000 3528 6 st_data_i[59]
port 308 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 st_data_i[5]
port 309 nsew signal input
rlabel metal2 s 4526 89200 4582 90000 6 st_data_i[60]
port 310 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 st_data_i[61]
port 311 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 st_data_i[62]
port 312 nsew signal input
rlabel metal2 s 47030 89200 47086 90000 6 st_data_i[63]
port 313 nsew signal input
rlabel metal3 s 139200 51008 140000 51128 6 st_data_i[6]
port 314 nsew signal input
rlabel metal2 s 56046 89200 56102 90000 6 st_data_i[7]
port 315 nsew signal input
rlabel metal3 s 139200 13608 140000 13728 6 st_data_i[8]
port 316 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 st_data_i[9]
port 317 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 tag_chip_en
port 318 nsew signal output
rlabel metal3 s 139200 37408 140000 37528 6 tag_data_in[0]
port 319 nsew signal output
rlabel metal2 s 73434 89200 73490 90000 6 tag_data_in[10]
port 320 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 tag_data_in[11]
port 321 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 tag_data_in[12]
port 322 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 tag_data_in[13]
port 323 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 tag_data_in[14]
port 324 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 tag_data_in[15]
port 325 nsew signal output
rlabel metal2 s 1950 89200 2006 90000 6 tag_data_in[16]
port 326 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 tag_data_in[17]
port 327 nsew signal output
rlabel metal2 s 63130 89200 63186 90000 6 tag_data_in[18]
port 328 nsew signal output
rlabel metal3 s 139200 8168 140000 8288 6 tag_data_in[19]
port 329 nsew signal output
rlabel metal2 s 662 89200 718 90000 6 tag_data_in[1]
port 330 nsew signal output
rlabel metal3 s 139200 688 140000 808 6 tag_data_in[20]
port 331 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 tag_data_in[21]
port 332 nsew signal output
rlabel metal2 s 74722 89200 74778 90000 6 tag_data_in[22]
port 333 nsew signal output
rlabel metal2 s 18 89200 74 90000 6 tag_data_in[23]
port 334 nsew signal output
rlabel metal3 s 139200 23808 140000 23928 6 tag_data_in[24]
port 335 nsew signal output
rlabel metal3 s 139200 73448 140000 73568 6 tag_data_in[25]
port 336 nsew signal output
rlabel metal3 s 139200 85688 140000 85808 6 tag_data_in[26]
port 337 nsew signal output
rlabel metal2 s 117870 89200 117926 90000 6 tag_data_in[27]
port 338 nsew signal output
rlabel metal3 s 139200 72088 140000 72208 6 tag_data_in[28]
port 339 nsew signal output
rlabel metal2 s 79874 89200 79930 90000 6 tag_data_in[29]
port 340 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 tag_data_in[2]
port 341 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 tag_data_in[30]
port 342 nsew signal output
rlabel metal2 s 35438 89200 35494 90000 6 tag_data_in[31]
port 343 nsew signal output
rlabel metal3 s 139200 28568 140000 28688 6 tag_data_in[3]
port 344 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 tag_data_in[4]
port 345 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 tag_data_in[5]
port 346 nsew signal output
rlabel metal3 s 139200 53728 140000 53848 6 tag_data_in[6]
port 347 nsew signal output
rlabel metal3 s 139200 39448 140000 39568 6 tag_data_in[7]
port 348 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 tag_data_in[8]
port 349 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 tag_data_in[9]
port 350 nsew signal output
rlabel metal2 s 30286 89200 30342 90000 6 tag_index[0]
port 351 nsew signal output
rlabel metal3 s 139200 66648 140000 66768 6 tag_index[1]
port 352 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 tag_index[2]
port 353 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 tag_index[3]
port 354 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 tag_index[4]
port 355 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 tag_index[5]
port 356 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 tag_index[6]
port 357 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 tag_index[7]
port 358 nsew signal output
rlabel metal3 s 139200 55768 140000 55888 6 tag_out[0]
port 359 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 tag_out[10]
port 360 nsew signal input
rlabel metal2 s 95974 89200 96030 90000 6 tag_out[11]
port 361 nsew signal input
rlabel metal2 s 79230 89200 79286 90000 6 tag_out[12]
port 362 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 tag_out[13]
port 363 nsew signal input
rlabel metal3 s 139200 67328 140000 67448 6 tag_out[14]
port 364 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 tag_out[15]
port 365 nsew signal input
rlabel metal2 s 18050 89200 18106 90000 6 tag_out[16]
port 366 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 tag_out[17]
port 367 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 tag_out[18]
port 368 nsew signal input
rlabel metal2 s 119802 89200 119858 90000 6 tag_out[19]
port 369 nsew signal input
rlabel metal2 s 112718 89200 112774 90000 6 tag_out[1]
port 370 nsew signal input
rlabel metal2 s 132038 89200 132094 90000 6 tag_out[20]
port 371 nsew signal input
rlabel metal2 s 137190 89200 137246 90000 6 tag_out[21]
port 372 nsew signal input
rlabel metal2 s 137834 89200 137890 90000 6 tag_out[22]
port 373 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 tag_out[23]
port 374 nsew signal input
rlabel metal2 s 101770 89200 101826 90000 6 tag_out[24]
port 375 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 tag_out[25]
port 376 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 tag_out[26]
port 377 nsew signal input
rlabel metal2 s 25778 89200 25834 90000 6 tag_out[27]
port 378 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 tag_out[28]
port 379 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 tag_out[29]
port 380 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 tag_out[2]
port 381 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 tag_out[30]
port 382 nsew signal input
rlabel metal2 s 39302 89200 39358 90000 6 tag_out[31]
port 383 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 tag_out[3]
port 384 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 tag_out[4]
port 385 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 tag_out[5]
port 386 nsew signal input
rlabel metal2 s 97262 89200 97318 90000 6 tag_out[6]
port 387 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 tag_out[7]
port 388 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 tag_out[8]
port 389 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 tag_out[9]
port 390 nsew signal input
rlabel metal3 s 139200 45568 140000 45688 6 tag_write_en
port 391 nsew signal output
rlabel metal3 s 139200 68688 140000 68808 6 type_i[0]
port 392 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 type_i[1]
port 393 nsew signal input
rlabel metal2 s 36082 89200 36138 90000 6 type_i[2]
port 394 nsew signal input
rlabel metal4 s 4208 2128 4528 87632 6 vccd1
port 395 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 87632 6 vccd1
port 395 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 87632 6 vccd1
port 395 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 87632 6 vccd1
port 395 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 87632 6 vccd1
port 395 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 87632 6 vssd1
port 396 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 87632 6 vssd1
port 396 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 87632 6 vssd1
port 396 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 87632 6 vssd1
port 396 nsew ground bidirectional
rlabel metal3 s 0 35368 800 35488 6 wb_ack_i
port 397 nsew signal input
rlabel metal2 s 12898 89200 12954 90000 6 wb_adr_o[0]
port 398 nsew signal output
rlabel metal2 s 80518 89200 80574 90000 6 wb_adr_o[10]
port 399 nsew signal output
rlabel metal3 s 139200 47608 140000 47728 6 wb_adr_o[11]
port 400 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 wb_adr_o[12]
port 401 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 wb_adr_o[13]
port 402 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 wb_adr_o[14]
port 403 nsew signal output
rlabel metal2 s 72146 89200 72202 90000 6 wb_adr_o[15]
port 404 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 wb_adr_o[16]
port 405 nsew signal output
rlabel metal2 s 29642 89200 29698 90000 6 wb_adr_o[17]
port 406 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wb_adr_o[18]
port 407 nsew signal output
rlabel metal3 s 139200 44888 140000 45008 6 wb_adr_o[19]
port 408 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 wb_adr_o[1]
port 409 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 wb_adr_o[20]
port 410 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 wb_adr_o[21]
port 411 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 wb_adr_o[22]
port 412 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 wb_adr_o[23]
port 413 nsew signal output
rlabel metal2 s 106922 89200 106978 90000 6 wb_adr_o[24]
port 414 nsew signal output
rlabel metal3 s 139200 76848 140000 76968 6 wb_adr_o[25]
port 415 nsew signal output
rlabel metal2 s 33506 89200 33562 90000 6 wb_adr_o[26]
port 416 nsew signal output
rlabel metal2 s 44454 89200 44510 90000 6 wb_adr_o[27]
port 417 nsew signal output
rlabel metal3 s 139200 1368 140000 1488 6 wb_adr_o[28]
port 418 nsew signal output
rlabel metal2 s 27066 89200 27122 90000 6 wb_adr_o[29]
port 419 nsew signal output
rlabel metal3 s 139200 22448 140000 22568 6 wb_adr_o[2]
port 420 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 wb_adr_o[30]
port 421 nsew signal output
rlabel metal2 s 59910 89200 59966 90000 6 wb_adr_o[31]
port 422 nsew signal output
rlabel metal2 s 12254 89200 12310 90000 6 wb_adr_o[3]
port 423 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wb_adr_o[4]
port 424 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 wb_adr_o[5]
port 425 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 wb_adr_o[6]
port 426 nsew signal output
rlabel metal3 s 139200 63928 140000 64048 6 wb_adr_o[7]
port 427 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 wb_adr_o[8]
port 428 nsew signal output
rlabel metal3 s 139200 55088 140000 55208 6 wb_adr_o[9]
port 429 nsew signal output
rlabel metal3 s 139200 17008 140000 17128 6 wb_bl_o[0]
port 430 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 wb_bl_o[1]
port 431 nsew signal output
rlabel metal2 s 85026 89200 85082 90000 6 wb_bl_o[2]
port 432 nsew signal output
rlabel metal2 s 118514 89200 118570 90000 6 wb_bl_o[3]
port 433 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 wb_bl_o[4]
port 434 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 wb_bl_o[5]
port 435 nsew signal output
rlabel metal3 s 139200 6128 140000 6248 6 wb_bl_o[6]
port 436 nsew signal output
rlabel metal2 s 23202 89200 23258 90000 6 wb_bl_o[7]
port 437 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 wb_bl_o[8]
port 438 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wb_bl_o[9]
port 439 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 wb_bry_o
port 440 nsew signal output
rlabel metal3 s 139200 50328 140000 50448 6 wb_cyc_o
port 441 nsew signal output
rlabel metal2 s 133326 89200 133382 90000 6 wb_dat_i[0]
port 442 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wb_dat_i[10]
port 443 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 wb_dat_i[11]
port 444 nsew signal input
rlabel metal3 s 139200 29248 140000 29368 6 wb_dat_i[12]
port 445 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 wb_dat_i[13]
port 446 nsew signal input
rlabel metal2 s 102414 89200 102470 90000 6 wb_dat_i[14]
port 447 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 wb_dat_i[15]
port 448 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wb_dat_i[16]
port 449 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wb_dat_i[17]
port 450 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 wb_dat_i[18]
port 451 nsew signal input
rlabel metal3 s 139200 10208 140000 10328 6 wb_dat_i[19]
port 452 nsew signal input
rlabel metal2 s 50250 89200 50306 90000 6 wb_dat_i[1]
port 453 nsew signal input
rlabel metal3 s 139200 84328 140000 84448 6 wb_dat_i[20]
port 454 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 wb_dat_i[21]
port 455 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 wb_dat_i[22]
port 456 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 wb_dat_i[23]
port 457 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wb_dat_i[24]
port 458 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wb_dat_i[25]
port 459 nsew signal input
rlabel metal3 s 139200 40128 140000 40248 6 wb_dat_i[26]
port 460 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 wb_dat_i[27]
port 461 nsew signal input
rlabel metal2 s 95330 89200 95386 90000 6 wb_dat_i[28]
port 462 nsew signal input
rlabel metal2 s 123022 89200 123078 90000 6 wb_dat_i[29]
port 463 nsew signal input
rlabel metal2 s 21914 89200 21970 90000 6 wb_dat_i[2]
port 464 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wb_dat_i[30]
port 465 nsew signal input
rlabel metal3 s 139200 49648 140000 49768 6 wb_dat_i[31]
port 466 nsew signal input
rlabel metal2 s 127530 89200 127586 90000 6 wb_dat_i[3]
port 467 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 wb_dat_i[4]
port 468 nsew signal input
rlabel metal3 s 139200 71408 140000 71528 6 wb_dat_i[5]
port 469 nsew signal input
rlabel metal3 s 139200 14288 140000 14408 6 wb_dat_i[6]
port 470 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 wb_dat_i[7]
port 471 nsew signal input
rlabel metal2 s 114650 89200 114706 90000 6 wb_dat_i[8]
port 472 nsew signal input
rlabel metal2 s 45742 89200 45798 90000 6 wb_dat_i[9]
port 473 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wb_dat_o[0]
port 474 nsew signal output
rlabel metal3 s 139200 48288 140000 48408 6 wb_dat_o[10]
port 475 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 wb_dat_o[11]
port 476 nsew signal output
rlabel metal3 s 139200 10888 140000 11008 6 wb_dat_o[12]
port 477 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 wb_dat_o[13]
port 478 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 wb_dat_o[14]
port 479 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wb_dat_o[15]
port 480 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 wb_dat_o[16]
port 481 nsew signal output
rlabel metal3 s 139200 26528 140000 26648 6 wb_dat_o[17]
port 482 nsew signal output
rlabel metal2 s 110786 89200 110842 90000 6 wb_dat_o[18]
port 483 nsew signal output
rlabel metal3 s 139200 82288 140000 82408 6 wb_dat_o[19]
port 484 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 wb_dat_o[1]
port 485 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wb_dat_o[20]
port 486 nsew signal output
rlabel metal3 s 139200 42848 140000 42968 6 wb_dat_o[21]
port 487 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wb_dat_o[22]
port 488 nsew signal output
rlabel metal3 s 139200 85008 140000 85128 6 wb_dat_o[23]
port 489 nsew signal output
rlabel metal2 s 107566 89200 107622 90000 6 wb_dat_o[24]
port 490 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 wb_dat_o[25]
port 491 nsew signal output
rlabel metal2 s 104346 89200 104402 90000 6 wb_dat_o[26]
port 492 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 wb_dat_o[27]
port 493 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 wb_dat_o[28]
port 494 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 wb_dat_o[29]
port 495 nsew signal output
rlabel metal2 s 18 0 74 800 6 wb_dat_o[2]
port 496 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 wb_dat_o[30]
port 497 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 wb_dat_o[31]
port 498 nsew signal output
rlabel metal2 s 7746 89200 7802 90000 6 wb_dat_o[3]
port 499 nsew signal output
rlabel metal2 s 54758 89200 54814 90000 6 wb_dat_o[4]
port 500 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 wb_dat_o[5]
port 501 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wb_dat_o[6]
port 502 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wb_dat_o[7]
port 503 nsew signal output
rlabel metal2 s 83094 89200 83150 90000 6 wb_dat_o[8]
port 504 nsew signal output
rlabel metal2 s 57334 89200 57390 90000 6 wb_dat_o[9]
port 505 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 wb_sel_o[0]
port 506 nsew signal output
rlabel metal2 s 103058 89200 103114 90000 6 wb_sel_o[1]
port 507 nsew signal output
rlabel metal3 s 139200 5448 140000 5568 6 wb_sel_o[2]
port 508 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 wb_sel_o[3]
port 509 nsew signal output
rlabel metal3 s 139200 64608 140000 64728 6 wb_stb_o
port 510 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wb_we_o
port 511 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 write_data_mask_1[0]
port 512 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 write_data_mask_1[1]
port 513 nsew signal output
rlabel metal3 s 139200 60528 140000 60648 6 write_data_mask_1[2]
port 514 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 write_data_mask_1[3]
port 515 nsew signal output
rlabel metal2 s 100482 89200 100538 90000 6 write_data_mask_2[0]
port 516 nsew signal output
rlabel metal2 s 98550 89200 98606 90000 6 write_data_mask_2[1]
port 517 nsew signal output
rlabel metal2 s 17406 89200 17462 90000 6 write_data_mask_2[2]
port 518 nsew signal output
rlabel metal2 s 38014 89200 38070 90000 6 write_data_mask_2[3]
port 519 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 write_tag_mask[0]
port 520 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 write_tag_mask[1]
port 521 nsew signal output
rlabel metal2 s 7102 89200 7158 90000 6 write_tag_mask[2]
port 522 nsew signal output
rlabel metal3 s 139200 29928 140000 30048 6 write_tag_mask[3]
port 523 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 140000 90000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23104550
string GDS_FILE /root/hellochip/openlane/lidinterface/runs/22_09_13_01_32/results/signoff/l1dcache.magic.gds
string GDS_START 1130078
<< end >>

