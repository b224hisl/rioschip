VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_function_generator
  CLASS BLOCK ;
  FOREIGN wrapped_function_generator ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 260.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 159.840 250.000 160.440 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 256.000 125.950 260.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 78.240 250.000 78.840 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 256.000 106.630 260.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 10.240 250.000 10.840 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 91.840 250.000 92.440 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 105.440 250.000 106.040 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 163.240 250.000 163.840 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 115.640 250.000 116.240 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 256.000 13.250 260.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 256.000 232.210 260.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 256.000 45.450 260.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 256.000 158.150 260.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 238.040 250.000 238.640 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 102.040 250.000 102.640 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 256.000 177.470 260.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 13.640 250.000 14.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 256.000 19.690 260.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 122.440 250.000 123.040 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 256.000 39.010 260.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 217.640 250.000 218.240 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 23.840 250.000 24.440 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 256.000 216.110 260.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 234.640 250.000 235.240 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 256.000 225.770 260.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 258.440 250.000 259.040 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 256.000 122.730 260.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 142.840 250.000 143.440 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 256.000 6.810 260.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 256.000 248.310 260.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 256.000 113.070 260.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 227.840 250.000 228.440 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 183.640 250.000 184.240 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 85.040 250.000 85.640 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 248.240 250.000 248.840 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 81.640 250.000 82.240 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 256.000 180.690 260.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 221.040 250.000 221.640 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 47.640 250.000 48.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 61.240 250.000 61.840 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 256.000 187.130 260.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 256.000 193.570 260.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 256.000 77.650 260.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 17.040 250.000 17.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 256.000 174.250 260.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 256.000 74.430 260.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 37.440 250.000 38.040 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 176.840 250.000 177.440 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 256.000 142.050 260.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 231.240 250.000 231.840 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 54.440 250.000 55.040 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 256.000 135.610 260.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 256.000 241.870 260.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 256.000 228.990 260.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 256.000 200.010 260.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 256.000 51.890 260.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 256.000 35.790 260.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 170.040 250.000 170.640 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 256.000 42.230 260.000 ;
    END
  END io_out[9]
  PIN rambus_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END rambus_wb_ack_i
  PIN rambus_wb_adr_o[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 200.640 250.000 201.240 ;
    END
  END rambus_wb_adr_o[0]
  PIN rambus_wb_adr_o[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END rambus_wb_adr_o[1]
  PIN rambus_wb_adr_o[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 256.000 55.110 260.000 ;
    END
  END rambus_wb_adr_o[2]
  PIN rambus_wb_adr_o[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 30.640 250.000 31.240 ;
    END
  END rambus_wb_adr_o[3]
  PIN rambus_wb_adr_o[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 255.040 250.000 255.640 ;
    END
  END rambus_wb_adr_o[4]
  PIN rambus_wb_adr_o[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 88.440 250.000 89.040 ;
    END
  END rambus_wb_adr_o[5]
  PIN rambus_wb_adr_o[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 34.040 250.000 34.640 ;
    END
  END rambus_wb_adr_o[6]
  PIN rambus_wb_adr_o[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 146.240 250.000 146.840 ;
    END
  END rambus_wb_adr_o[7]
  PIN rambus_wb_adr_o[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END rambus_wb_adr_o[8]
  PIN rambus_wb_adr_o[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END rambus_wb_adr_o[9]
  PIN rambus_wb_clk_o
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END rambus_wb_clk_o
  PIN rambus_wb_cyc_o
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 256.000 26.130 260.000 ;
    END
  END rambus_wb_cyc_o
  PIN rambus_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 256.000 67.990 260.000 ;
    END
  END rambus_wb_dat_i[0]
  PIN rambus_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END rambus_wb_dat_i[10]
  PIN rambus_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END rambus_wb_dat_i[11]
  PIN rambus_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 3.440 250.000 4.040 ;
    END
  END rambus_wb_dat_i[12]
  PIN rambus_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 68.040 250.000 68.640 ;
    END
  END rambus_wb_dat_i[13]
  PIN rambus_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 256.000 109.850 260.000 ;
    END
  END rambus_wb_dat_i[14]
  PIN rambus_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 256.000 64.770 260.000 ;
    END
  END rambus_wb_dat_i[15]
  PIN rambus_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 256.000 90.530 260.000 ;
    END
  END rambus_wb_dat_i[16]
  PIN rambus_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END rambus_wb_dat_i[17]
  PIN rambus_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END rambus_wb_dat_i[18]
  PIN rambus_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END rambus_wb_dat_i[19]
  PIN rambus_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END rambus_wb_dat_i[1]
  PIN rambus_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END rambus_wb_dat_i[20]
  PIN rambus_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 256.000 80.870 260.000 ;
    END
  END rambus_wb_dat_i[21]
  PIN rambus_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 40.840 250.000 41.440 ;
    END
  END rambus_wb_dat_i[22]
  PIN rambus_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 156.440 250.000 157.040 ;
    END
  END rambus_wb_dat_i[23]
  PIN rambus_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 166.640 250.000 167.240 ;
    END
  END rambus_wb_dat_i[24]
  PIN rambus_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 193.840 250.000 194.440 ;
    END
  END rambus_wb_dat_i[25]
  PIN rambus_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 256.000 119.510 260.000 ;
    END
  END rambus_wb_dat_i[26]
  PIN rambus_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END rambus_wb_dat_i[27]
  PIN rambus_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 256.000 0.370 260.000 ;
    END
  END rambus_wb_dat_i[28]
  PIN rambus_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 210.840 250.000 211.440 ;
    END
  END rambus_wb_dat_i[29]
  PIN rambus_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END rambus_wb_dat_i[2]
  PIN rambus_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 51.040 250.000 51.640 ;
    END
  END rambus_wb_dat_i[30]
  PIN rambus_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 256.000 71.210 260.000 ;
    END
  END rambus_wb_dat_i[31]
  PIN rambus_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 149.640 250.000 150.240 ;
    END
  END rambus_wb_dat_i[3]
  PIN rambus_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 119.040 250.000 119.640 ;
    END
  END rambus_wb_dat_i[4]
  PIN rambus_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END rambus_wb_dat_i[5]
  PIN rambus_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 256.000 22.910 260.000 ;
    END
  END rambus_wb_dat_i[6]
  PIN rambus_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END rambus_wb_dat_i[7]
  PIN rambus_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END rambus_wb_dat_i[8]
  PIN rambus_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 256.000 203.230 260.000 ;
    END
  END rambus_wb_dat_i[9]
  PIN rambus_wb_dat_o[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END rambus_wb_dat_o[0]
  PIN rambus_wb_dat_o[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END rambus_wb_dat_o[10]
  PIN rambus_wb_dat_o[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END rambus_wb_dat_o[11]
  PIN rambus_wb_dat_o[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END rambus_wb_dat_o[12]
  PIN rambus_wb_dat_o[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 173.440 250.000 174.040 ;
    END
  END rambus_wb_dat_o[13]
  PIN rambus_wb_dat_o[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END rambus_wb_dat_o[14]
  PIN rambus_wb_dat_o[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 256.000 212.890 260.000 ;
    END
  END rambus_wb_dat_o[15]
  PIN rambus_wb_dat_o[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END rambus_wb_dat_o[16]
  PIN rambus_wb_dat_o[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END rambus_wb_dat_o[17]
  PIN rambus_wb_dat_o[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END rambus_wb_dat_o[18]
  PIN rambus_wb_dat_o[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 256.000 103.410 260.000 ;
    END
  END rambus_wb_dat_o[19]
  PIN rambus_wb_dat_o[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END rambus_wb_dat_o[1]
  PIN rambus_wb_dat_o[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END rambus_wb_dat_o[20]
  PIN rambus_wb_dat_o[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END rambus_wb_dat_o[21]
  PIN rambus_wb_dat_o[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END rambus_wb_dat_o[22]
  PIN rambus_wb_dat_o[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 98.640 250.000 99.240 ;
    END
  END rambus_wb_dat_o[23]
  PIN rambus_wb_dat_o[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 256.000 154.930 260.000 ;
    END
  END rambus_wb_dat_o[24]
  PIN rambus_wb_dat_o[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END rambus_wb_dat_o[25]
  PIN rambus_wb_dat_o[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 256.000 116.290 260.000 ;
    END
  END rambus_wb_dat_o[26]
  PIN rambus_wb_dat_o[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END rambus_wb_dat_o[27]
  PIN rambus_wb_dat_o[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 251.640 250.000 252.240 ;
    END
  END rambus_wb_dat_o[28]
  PIN rambus_wb_dat_o[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END rambus_wb_dat_o[29]
  PIN rambus_wb_dat_o[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END rambus_wb_dat_o[2]
  PIN rambus_wb_dat_o[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 207.440 250.000 208.040 ;
    END
  END rambus_wb_dat_o[30]
  PIN rambus_wb_dat_o[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END rambus_wb_dat_o[31]
  PIN rambus_wb_dat_o[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 256.000 87.310 260.000 ;
    END
  END rambus_wb_dat_o[3]
  PIN rambus_wb_dat_o[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END rambus_wb_dat_o[4]
  PIN rambus_wb_dat_o[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 256.000 161.370 260.000 ;
    END
  END rambus_wb_dat_o[5]
  PIN rambus_wb_dat_o[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END rambus_wb_dat_o[6]
  PIN rambus_wb_dat_o[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 71.440 250.000 72.040 ;
    END
  END rambus_wb_dat_o[7]
  PIN rambus_wb_dat_o[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END rambus_wb_dat_o[8]
  PIN rambus_wb_dat_o[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 256.000 61.550 260.000 ;
    END
  END rambus_wb_dat_o[9]
  PIN rambus_wb_rst_o
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END rambus_wb_rst_o
  PIN rambus_wb_sel_o[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END rambus_wb_sel_o[0]
  PIN rambus_wb_sel_o[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 256.000 164.590 260.000 ;
    END
  END rambus_wb_sel_o[1]
  PIN rambus_wb_sel_o[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 256.000 48.670 260.000 ;
    END
  END rambus_wb_sel_o[2]
  PIN rambus_wb_sel_o[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END rambus_wb_sel_o[3]
  PIN rambus_wb_stb_o
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 256.000 148.490 260.000 ;
    END
  END rambus_wb_stb_o
  PIN rambus_wb_we_o
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END rambus_wb_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 247.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 247.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 247.760 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 6.840 250.000 7.440 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 256.000 132.390 260.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 256.000 190.350 260.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 256.000 100.190 260.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 256.000 32.570 260.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 139.440 250.000 140.040 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 256.000 222.550 260.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 27.240 250.000 27.840 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 256.000 96.970 260.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 256.000 145.270 260.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 112.240 250.000 112.840 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 204.040 250.000 204.640 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 256.000 245.090 260.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 74.840 250.000 75.440 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 256.000 238.650 260.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 44.240 250.000 44.840 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 256.000 129.170 260.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 190.440 250.000 191.040 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 256.000 3.590 260.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 256.000 16.470 260.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 256.000 10.030 260.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 108.840 250.000 109.440 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 256.000 209.670 260.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 244.840 250.000 245.440 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 256.000 58.330 260.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 129.240 250.000 129.840 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 241.440 250.000 242.040 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 180.240 250.000 180.840 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 256.000 235.430 260.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 256.000 93.750 260.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 136.040 250.000 136.640 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 57.840 250.000 58.440 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 95.240 250.000 95.840 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 256.000 219.330 260.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 214.240 250.000 214.840 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 0.040 250.000 0.640 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 132.640 250.000 133.240 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 224.440 250.000 225.040 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 256.000 206.450 260.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 20.440 250.000 21.040 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 256.000 196.790 260.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 256.000 138.830 260.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 256.000 84.090 260.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 256.000 183.910 260.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 64.640 250.000 65.240 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 197.240 250.000 197.840 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 187.040 250.000 187.640 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 256.000 171.030 260.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 256.000 167.810 260.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 256.000 29.350 260.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 125.840 250.000 126.440 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 247.605 ;
      LAYER met1 ;
        RECT 0.070 9.220 248.330 251.220 ;
      LAYER met2 ;
        RECT 0.650 255.720 3.030 258.925 ;
        RECT 3.870 255.720 6.250 258.925 ;
        RECT 7.090 255.720 9.470 258.925 ;
        RECT 10.310 255.720 12.690 258.925 ;
        RECT 13.530 255.720 15.910 258.925 ;
        RECT 16.750 255.720 19.130 258.925 ;
        RECT 19.970 255.720 22.350 258.925 ;
        RECT 23.190 255.720 25.570 258.925 ;
        RECT 26.410 255.720 28.790 258.925 ;
        RECT 29.630 255.720 32.010 258.925 ;
        RECT 32.850 255.720 35.230 258.925 ;
        RECT 36.070 255.720 38.450 258.925 ;
        RECT 39.290 255.720 41.670 258.925 ;
        RECT 42.510 255.720 44.890 258.925 ;
        RECT 45.730 255.720 48.110 258.925 ;
        RECT 48.950 255.720 51.330 258.925 ;
        RECT 52.170 255.720 54.550 258.925 ;
        RECT 55.390 255.720 57.770 258.925 ;
        RECT 58.610 255.720 60.990 258.925 ;
        RECT 61.830 255.720 64.210 258.925 ;
        RECT 65.050 255.720 67.430 258.925 ;
        RECT 68.270 255.720 70.650 258.925 ;
        RECT 71.490 255.720 73.870 258.925 ;
        RECT 74.710 255.720 77.090 258.925 ;
        RECT 77.930 255.720 80.310 258.925 ;
        RECT 81.150 255.720 83.530 258.925 ;
        RECT 84.370 255.720 86.750 258.925 ;
        RECT 87.590 255.720 89.970 258.925 ;
        RECT 90.810 255.720 93.190 258.925 ;
        RECT 94.030 255.720 96.410 258.925 ;
        RECT 97.250 255.720 99.630 258.925 ;
        RECT 100.470 255.720 102.850 258.925 ;
        RECT 103.690 255.720 106.070 258.925 ;
        RECT 106.910 255.720 109.290 258.925 ;
        RECT 110.130 255.720 112.510 258.925 ;
        RECT 113.350 255.720 115.730 258.925 ;
        RECT 116.570 255.720 118.950 258.925 ;
        RECT 119.790 255.720 122.170 258.925 ;
        RECT 123.010 255.720 125.390 258.925 ;
        RECT 126.230 255.720 128.610 258.925 ;
        RECT 129.450 255.720 131.830 258.925 ;
        RECT 132.670 255.720 135.050 258.925 ;
        RECT 135.890 255.720 138.270 258.925 ;
        RECT 139.110 255.720 141.490 258.925 ;
        RECT 142.330 255.720 144.710 258.925 ;
        RECT 145.550 255.720 147.930 258.925 ;
        RECT 148.770 255.720 154.370 258.925 ;
        RECT 155.210 255.720 157.590 258.925 ;
        RECT 158.430 255.720 160.810 258.925 ;
        RECT 161.650 255.720 164.030 258.925 ;
        RECT 164.870 255.720 167.250 258.925 ;
        RECT 168.090 255.720 170.470 258.925 ;
        RECT 171.310 255.720 173.690 258.925 ;
        RECT 174.530 255.720 176.910 258.925 ;
        RECT 177.750 255.720 180.130 258.925 ;
        RECT 180.970 255.720 183.350 258.925 ;
        RECT 184.190 255.720 186.570 258.925 ;
        RECT 187.410 255.720 189.790 258.925 ;
        RECT 190.630 255.720 193.010 258.925 ;
        RECT 193.850 255.720 196.230 258.925 ;
        RECT 197.070 255.720 199.450 258.925 ;
        RECT 200.290 255.720 202.670 258.925 ;
        RECT 203.510 255.720 205.890 258.925 ;
        RECT 206.730 255.720 209.110 258.925 ;
        RECT 209.950 255.720 212.330 258.925 ;
        RECT 213.170 255.720 215.550 258.925 ;
        RECT 216.390 255.720 218.770 258.925 ;
        RECT 219.610 255.720 221.990 258.925 ;
        RECT 222.830 255.720 225.210 258.925 ;
        RECT 226.050 255.720 228.430 258.925 ;
        RECT 229.270 255.720 231.650 258.925 ;
        RECT 232.490 255.720 234.870 258.925 ;
        RECT 235.710 255.720 238.090 258.925 ;
        RECT 238.930 255.720 241.310 258.925 ;
        RECT 242.150 255.720 244.530 258.925 ;
        RECT 245.370 255.720 247.750 258.925 ;
        RECT 0.100 4.280 248.300 255.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
        RECT 119.790 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 141.490 4.280 ;
        RECT 142.330 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.930 4.280 ;
        RECT 148.770 0.155 151.150 4.280 ;
        RECT 151.990 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 160.810 4.280 ;
        RECT 161.650 0.155 164.030 4.280 ;
        RECT 164.870 0.155 167.250 4.280 ;
        RECT 168.090 0.155 170.470 4.280 ;
        RECT 171.310 0.155 173.690 4.280 ;
        RECT 174.530 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 186.570 4.280 ;
        RECT 187.410 0.155 189.790 4.280 ;
        RECT 190.630 0.155 193.010 4.280 ;
        RECT 193.850 0.155 199.450 4.280 ;
        RECT 200.290 0.155 202.670 4.280 ;
        RECT 203.510 0.155 205.890 4.280 ;
        RECT 206.730 0.155 209.110 4.280 ;
        RECT 209.950 0.155 212.330 4.280 ;
        RECT 213.170 0.155 215.550 4.280 ;
        RECT 216.390 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.990 4.280 ;
        RECT 222.830 0.155 225.210 4.280 ;
        RECT 226.050 0.155 228.430 4.280 ;
        RECT 229.270 0.155 231.650 4.280 ;
        RECT 232.490 0.155 234.870 4.280 ;
        RECT 235.710 0.155 238.090 4.280 ;
        RECT 238.930 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 247.750 4.280 ;
      LAYER met3 ;
        RECT 4.400 258.040 245.600 258.905 ;
        RECT 4.000 256.040 246.000 258.040 ;
        RECT 4.400 254.640 245.600 256.040 ;
        RECT 4.000 252.640 246.000 254.640 ;
        RECT 4.400 251.240 245.600 252.640 ;
        RECT 4.000 249.240 246.000 251.240 ;
        RECT 4.400 247.840 245.600 249.240 ;
        RECT 4.000 245.840 246.000 247.840 ;
        RECT 4.400 244.440 245.600 245.840 ;
        RECT 4.000 242.440 246.000 244.440 ;
        RECT 4.400 241.040 245.600 242.440 ;
        RECT 4.000 239.040 246.000 241.040 ;
        RECT 4.400 237.640 245.600 239.040 ;
        RECT 4.000 235.640 246.000 237.640 ;
        RECT 4.400 234.240 245.600 235.640 ;
        RECT 4.000 232.240 246.000 234.240 ;
        RECT 4.400 230.840 245.600 232.240 ;
        RECT 4.000 228.840 246.000 230.840 ;
        RECT 4.400 227.440 245.600 228.840 ;
        RECT 4.000 225.440 246.000 227.440 ;
        RECT 4.400 224.040 245.600 225.440 ;
        RECT 4.000 222.040 246.000 224.040 ;
        RECT 4.400 220.640 245.600 222.040 ;
        RECT 4.000 218.640 246.000 220.640 ;
        RECT 4.400 217.240 245.600 218.640 ;
        RECT 4.000 215.240 246.000 217.240 ;
        RECT 4.400 213.840 245.600 215.240 ;
        RECT 4.000 211.840 246.000 213.840 ;
        RECT 4.000 210.440 245.600 211.840 ;
        RECT 4.000 208.440 246.000 210.440 ;
        RECT 4.400 207.040 245.600 208.440 ;
        RECT 4.000 205.040 246.000 207.040 ;
        RECT 4.400 203.640 245.600 205.040 ;
        RECT 4.000 201.640 246.000 203.640 ;
        RECT 4.400 200.240 245.600 201.640 ;
        RECT 4.000 198.240 246.000 200.240 ;
        RECT 4.400 196.840 245.600 198.240 ;
        RECT 4.000 194.840 246.000 196.840 ;
        RECT 4.400 193.440 245.600 194.840 ;
        RECT 4.000 191.440 246.000 193.440 ;
        RECT 4.400 190.040 245.600 191.440 ;
        RECT 4.000 188.040 246.000 190.040 ;
        RECT 4.400 186.640 245.600 188.040 ;
        RECT 4.000 184.640 246.000 186.640 ;
        RECT 4.400 183.240 245.600 184.640 ;
        RECT 4.000 181.240 246.000 183.240 ;
        RECT 4.400 179.840 245.600 181.240 ;
        RECT 4.000 177.840 246.000 179.840 ;
        RECT 4.400 176.440 245.600 177.840 ;
        RECT 4.000 174.440 246.000 176.440 ;
        RECT 4.400 173.040 245.600 174.440 ;
        RECT 4.000 171.040 246.000 173.040 ;
        RECT 4.400 169.640 245.600 171.040 ;
        RECT 4.000 167.640 246.000 169.640 ;
        RECT 4.400 166.240 245.600 167.640 ;
        RECT 4.000 164.240 246.000 166.240 ;
        RECT 4.400 162.840 245.600 164.240 ;
        RECT 4.000 160.840 246.000 162.840 ;
        RECT 4.400 159.440 245.600 160.840 ;
        RECT 4.000 157.440 246.000 159.440 ;
        RECT 4.400 156.040 245.600 157.440 ;
        RECT 4.000 154.040 246.000 156.040 ;
        RECT 4.400 152.640 246.000 154.040 ;
        RECT 4.000 150.640 246.000 152.640 ;
        RECT 4.400 149.240 245.600 150.640 ;
        RECT 4.000 147.240 246.000 149.240 ;
        RECT 4.400 145.840 245.600 147.240 ;
        RECT 4.000 143.840 246.000 145.840 ;
        RECT 4.400 142.440 245.600 143.840 ;
        RECT 4.000 140.440 246.000 142.440 ;
        RECT 4.400 139.040 245.600 140.440 ;
        RECT 4.000 137.040 246.000 139.040 ;
        RECT 4.400 135.640 245.600 137.040 ;
        RECT 4.000 133.640 246.000 135.640 ;
        RECT 4.400 132.240 245.600 133.640 ;
        RECT 4.000 130.240 246.000 132.240 ;
        RECT 4.400 128.840 245.600 130.240 ;
        RECT 4.000 126.840 246.000 128.840 ;
        RECT 4.400 125.440 245.600 126.840 ;
        RECT 4.000 123.440 246.000 125.440 ;
        RECT 4.400 122.040 245.600 123.440 ;
        RECT 4.000 120.040 246.000 122.040 ;
        RECT 4.400 118.640 245.600 120.040 ;
        RECT 4.000 116.640 246.000 118.640 ;
        RECT 4.400 115.240 245.600 116.640 ;
        RECT 4.000 113.240 246.000 115.240 ;
        RECT 4.400 111.840 245.600 113.240 ;
        RECT 4.000 109.840 246.000 111.840 ;
        RECT 4.400 108.440 245.600 109.840 ;
        RECT 4.000 106.440 246.000 108.440 ;
        RECT 4.400 105.040 245.600 106.440 ;
        RECT 4.000 103.040 246.000 105.040 ;
        RECT 4.400 101.640 245.600 103.040 ;
        RECT 4.000 99.640 246.000 101.640 ;
        RECT 4.400 98.240 245.600 99.640 ;
        RECT 4.000 96.240 246.000 98.240 ;
        RECT 4.400 94.840 245.600 96.240 ;
        RECT 4.000 92.840 246.000 94.840 ;
        RECT 4.400 91.440 245.600 92.840 ;
        RECT 4.000 89.440 246.000 91.440 ;
        RECT 4.400 88.040 245.600 89.440 ;
        RECT 4.000 86.040 246.000 88.040 ;
        RECT 4.400 84.640 245.600 86.040 ;
        RECT 4.000 82.640 246.000 84.640 ;
        RECT 4.400 81.240 245.600 82.640 ;
        RECT 4.000 79.240 246.000 81.240 ;
        RECT 4.400 77.840 245.600 79.240 ;
        RECT 4.000 75.840 246.000 77.840 ;
        RECT 4.400 74.440 245.600 75.840 ;
        RECT 4.000 72.440 246.000 74.440 ;
        RECT 4.400 71.040 245.600 72.440 ;
        RECT 4.000 69.040 246.000 71.040 ;
        RECT 4.400 67.640 245.600 69.040 ;
        RECT 4.000 65.640 246.000 67.640 ;
        RECT 4.400 64.240 245.600 65.640 ;
        RECT 4.000 62.240 246.000 64.240 ;
        RECT 4.400 60.840 245.600 62.240 ;
        RECT 4.000 58.840 246.000 60.840 ;
        RECT 4.400 57.440 245.600 58.840 ;
        RECT 4.000 55.440 246.000 57.440 ;
        RECT 4.400 54.040 245.600 55.440 ;
        RECT 4.000 52.040 246.000 54.040 ;
        RECT 4.400 50.640 245.600 52.040 ;
        RECT 4.000 48.640 246.000 50.640 ;
        RECT 4.400 47.240 245.600 48.640 ;
        RECT 4.000 45.240 246.000 47.240 ;
        RECT 4.400 43.840 245.600 45.240 ;
        RECT 4.000 41.840 246.000 43.840 ;
        RECT 4.400 40.440 245.600 41.840 ;
        RECT 4.000 38.440 246.000 40.440 ;
        RECT 4.400 37.040 245.600 38.440 ;
        RECT 4.000 35.040 246.000 37.040 ;
        RECT 4.400 33.640 245.600 35.040 ;
        RECT 4.000 31.640 246.000 33.640 ;
        RECT 4.400 30.240 245.600 31.640 ;
        RECT 4.000 28.240 246.000 30.240 ;
        RECT 4.400 26.840 245.600 28.240 ;
        RECT 4.000 24.840 246.000 26.840 ;
        RECT 4.400 23.440 245.600 24.840 ;
        RECT 4.000 21.440 246.000 23.440 ;
        RECT 4.400 20.040 245.600 21.440 ;
        RECT 4.000 18.040 246.000 20.040 ;
        RECT 4.400 16.640 245.600 18.040 ;
        RECT 4.000 14.640 246.000 16.640 ;
        RECT 4.400 13.240 245.600 14.640 ;
        RECT 4.000 11.240 246.000 13.240 ;
        RECT 4.400 9.840 245.600 11.240 ;
        RECT 4.000 7.840 246.000 9.840 ;
        RECT 4.400 6.440 245.600 7.840 ;
        RECT 4.000 4.440 246.000 6.440 ;
        RECT 4.400 3.040 245.600 4.440 ;
        RECT 4.000 1.040 246.000 3.040 ;
        RECT 4.000 0.175 245.600 1.040 ;
      LAYER met4 ;
        RECT 100.575 11.735 163.465 109.985 ;
  END
END wrapped_function_generator
END LIBRARY

