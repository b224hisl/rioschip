magic
tech sky130B
magscale 1 2
timestamp 1663004302
<< obsli1 >>
rect 1104 2159 118864 207825
<< obsm1 >>
rect 14 1368 119862 207856
<< metal2 >>
rect 18 209200 74 210000
rect 662 209200 718 210000
rect 1306 209200 1362 210000
rect 1950 209200 2006 210000
rect 2594 209200 2650 210000
rect 3238 209200 3294 210000
rect 3882 209200 3938 210000
rect 4526 209200 4582 210000
rect 5170 209200 5226 210000
rect 6458 209200 6514 210000
rect 7102 209200 7158 210000
rect 7746 209200 7802 210000
rect 8390 209200 8446 210000
rect 9034 209200 9090 210000
rect 9678 209200 9734 210000
rect 10322 209200 10378 210000
rect 10966 209200 11022 210000
rect 11610 209200 11666 210000
rect 12254 209200 12310 210000
rect 12898 209200 12954 210000
rect 13542 209200 13598 210000
rect 14186 209200 14242 210000
rect 14830 209200 14886 210000
rect 15474 209200 15530 210000
rect 16118 209200 16174 210000
rect 16762 209200 16818 210000
rect 17406 209200 17462 210000
rect 18050 209200 18106 210000
rect 18694 209200 18750 210000
rect 19338 209200 19394 210000
rect 19982 209200 20038 210000
rect 20626 209200 20682 210000
rect 21270 209200 21326 210000
rect 21914 209200 21970 210000
rect 22558 209200 22614 210000
rect 23202 209200 23258 210000
rect 23846 209200 23902 210000
rect 24490 209200 24546 210000
rect 25134 209200 25190 210000
rect 25778 209200 25834 210000
rect 26422 209200 26478 210000
rect 27066 209200 27122 210000
rect 27710 209200 27766 210000
rect 28354 209200 28410 210000
rect 29642 209200 29698 210000
rect 30286 209200 30342 210000
rect 30930 209200 30986 210000
rect 31574 209200 31630 210000
rect 32218 209200 32274 210000
rect 32862 209200 32918 210000
rect 33506 209200 33562 210000
rect 34150 209200 34206 210000
rect 34794 209200 34850 210000
rect 35438 209200 35494 210000
rect 36082 209200 36138 210000
rect 36726 209200 36782 210000
rect 37370 209200 37426 210000
rect 38014 209200 38070 210000
rect 38658 209200 38714 210000
rect 39302 209200 39358 210000
rect 39946 209200 40002 210000
rect 40590 209200 40646 210000
rect 41234 209200 41290 210000
rect 41878 209200 41934 210000
rect 42522 209200 42578 210000
rect 43166 209200 43222 210000
rect 43810 209200 43866 210000
rect 44454 209200 44510 210000
rect 45098 209200 45154 210000
rect 45742 209200 45798 210000
rect 46386 209200 46442 210000
rect 47030 209200 47086 210000
rect 47674 209200 47730 210000
rect 48318 209200 48374 210000
rect 48962 209200 49018 210000
rect 49606 209200 49662 210000
rect 50250 209200 50306 210000
rect 50894 209200 50950 210000
rect 52182 209200 52238 210000
rect 52826 209200 52882 210000
rect 53470 209200 53526 210000
rect 54114 209200 54170 210000
rect 54758 209200 54814 210000
rect 55402 209200 55458 210000
rect 56046 209200 56102 210000
rect 56690 209200 56746 210000
rect 57334 209200 57390 210000
rect 57978 209200 58034 210000
rect 58622 209200 58678 210000
rect 59266 209200 59322 210000
rect 59910 209200 59966 210000
rect 60554 209200 60610 210000
rect 61198 209200 61254 210000
rect 61842 209200 61898 210000
rect 62486 209200 62542 210000
rect 63130 209200 63186 210000
rect 63774 209200 63830 210000
rect 64418 209200 64474 210000
rect 65062 209200 65118 210000
rect 65706 209200 65762 210000
rect 66350 209200 66406 210000
rect 66994 209200 67050 210000
rect 67638 209200 67694 210000
rect 68282 209200 68338 210000
rect 68926 209200 68982 210000
rect 69570 209200 69626 210000
rect 70214 209200 70270 210000
rect 70858 209200 70914 210000
rect 71502 209200 71558 210000
rect 72146 209200 72202 210000
rect 72790 209200 72846 210000
rect 73434 209200 73490 210000
rect 74078 209200 74134 210000
rect 75366 209200 75422 210000
rect 76010 209200 76066 210000
rect 76654 209200 76710 210000
rect 77298 209200 77354 210000
rect 77942 209200 77998 210000
rect 78586 209200 78642 210000
rect 79230 209200 79286 210000
rect 79874 209200 79930 210000
rect 80518 209200 80574 210000
rect 81162 209200 81218 210000
rect 81806 209200 81862 210000
rect 82450 209200 82506 210000
rect 83094 209200 83150 210000
rect 83738 209200 83794 210000
rect 84382 209200 84438 210000
rect 85026 209200 85082 210000
rect 85670 209200 85726 210000
rect 86314 209200 86370 210000
rect 86958 209200 87014 210000
rect 87602 209200 87658 210000
rect 88246 209200 88302 210000
rect 88890 209200 88946 210000
rect 89534 209200 89590 210000
rect 90178 209200 90234 210000
rect 90822 209200 90878 210000
rect 91466 209200 91522 210000
rect 92110 209200 92166 210000
rect 92754 209200 92810 210000
rect 93398 209200 93454 210000
rect 94042 209200 94098 210000
rect 94686 209200 94742 210000
rect 95330 209200 95386 210000
rect 95974 209200 96030 210000
rect 96618 209200 96674 210000
rect 97906 209200 97962 210000
rect 98550 209200 98606 210000
rect 99194 209200 99250 210000
rect 99838 209200 99894 210000
rect 100482 209200 100538 210000
rect 101126 209200 101182 210000
rect 101770 209200 101826 210000
rect 102414 209200 102470 210000
rect 103058 209200 103114 210000
rect 103702 209200 103758 210000
rect 104346 209200 104402 210000
rect 104990 209200 105046 210000
rect 105634 209200 105690 210000
rect 106278 209200 106334 210000
rect 106922 209200 106978 210000
rect 107566 209200 107622 210000
rect 108210 209200 108266 210000
rect 108854 209200 108910 210000
rect 109498 209200 109554 210000
rect 110142 209200 110198 210000
rect 110786 209200 110842 210000
rect 111430 209200 111486 210000
rect 112074 209200 112130 210000
rect 112718 209200 112774 210000
rect 113362 209200 113418 210000
rect 114006 209200 114062 210000
rect 114650 209200 114706 210000
rect 115294 209200 115350 210000
rect 115938 209200 115994 210000
rect 116582 209200 116638 210000
rect 117226 209200 117282 210000
rect 117870 209200 117926 210000
rect 118514 209200 118570 210000
rect 119158 209200 119214 210000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 84382 0 84438 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92754 0 92810 800
rect 93398 0 93454 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97262 0 97318 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99838 0 99894 800
rect 100482 0 100538 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 103702 0 103758 800
rect 104346 0 104402 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106278 0 106334 800
rect 106922 0 106978 800
rect 107566 0 107622 800
rect 108210 0 108266 800
rect 108854 0 108910 800
rect 109498 0 109554 800
rect 110142 0 110198 800
rect 110786 0 110842 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 112718 0 112774 800
rect 113362 0 113418 800
rect 114650 0 114706 800
rect 115294 0 115350 800
rect 115938 0 115994 800
rect 116582 0 116638 800
rect 117226 0 117282 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119158 0 119214 800
rect 119802 0 119858 800
<< obsm2 >>
rect 130 209144 606 209250
rect 774 209144 1250 209250
rect 1418 209144 1894 209250
rect 2062 209144 2538 209250
rect 2706 209144 3182 209250
rect 3350 209144 3826 209250
rect 3994 209144 4470 209250
rect 4638 209144 5114 209250
rect 5282 209144 6402 209250
rect 6570 209144 7046 209250
rect 7214 209144 7690 209250
rect 7858 209144 8334 209250
rect 8502 209144 8978 209250
rect 9146 209144 9622 209250
rect 9790 209144 10266 209250
rect 10434 209144 10910 209250
rect 11078 209144 11554 209250
rect 11722 209144 12198 209250
rect 12366 209144 12842 209250
rect 13010 209144 13486 209250
rect 13654 209144 14130 209250
rect 14298 209144 14774 209250
rect 14942 209144 15418 209250
rect 15586 209144 16062 209250
rect 16230 209144 16706 209250
rect 16874 209144 17350 209250
rect 17518 209144 17994 209250
rect 18162 209144 18638 209250
rect 18806 209144 19282 209250
rect 19450 209144 19926 209250
rect 20094 209144 20570 209250
rect 20738 209144 21214 209250
rect 21382 209144 21858 209250
rect 22026 209144 22502 209250
rect 22670 209144 23146 209250
rect 23314 209144 23790 209250
rect 23958 209144 24434 209250
rect 24602 209144 25078 209250
rect 25246 209144 25722 209250
rect 25890 209144 26366 209250
rect 26534 209144 27010 209250
rect 27178 209144 27654 209250
rect 27822 209144 28298 209250
rect 28466 209144 29586 209250
rect 29754 209144 30230 209250
rect 30398 209144 30874 209250
rect 31042 209144 31518 209250
rect 31686 209144 32162 209250
rect 32330 209144 32806 209250
rect 32974 209144 33450 209250
rect 33618 209144 34094 209250
rect 34262 209144 34738 209250
rect 34906 209144 35382 209250
rect 35550 209144 36026 209250
rect 36194 209144 36670 209250
rect 36838 209144 37314 209250
rect 37482 209144 37958 209250
rect 38126 209144 38602 209250
rect 38770 209144 39246 209250
rect 39414 209144 39890 209250
rect 40058 209144 40534 209250
rect 40702 209144 41178 209250
rect 41346 209144 41822 209250
rect 41990 209144 42466 209250
rect 42634 209144 43110 209250
rect 43278 209144 43754 209250
rect 43922 209144 44398 209250
rect 44566 209144 45042 209250
rect 45210 209144 45686 209250
rect 45854 209144 46330 209250
rect 46498 209144 46974 209250
rect 47142 209144 47618 209250
rect 47786 209144 48262 209250
rect 48430 209144 48906 209250
rect 49074 209144 49550 209250
rect 49718 209144 50194 209250
rect 50362 209144 50838 209250
rect 51006 209144 52126 209250
rect 52294 209144 52770 209250
rect 52938 209144 53414 209250
rect 53582 209144 54058 209250
rect 54226 209144 54702 209250
rect 54870 209144 55346 209250
rect 55514 209144 55990 209250
rect 56158 209144 56634 209250
rect 56802 209144 57278 209250
rect 57446 209144 57922 209250
rect 58090 209144 58566 209250
rect 58734 209144 59210 209250
rect 59378 209144 59854 209250
rect 60022 209144 60498 209250
rect 60666 209144 61142 209250
rect 61310 209144 61786 209250
rect 61954 209144 62430 209250
rect 62598 209144 63074 209250
rect 63242 209144 63718 209250
rect 63886 209144 64362 209250
rect 64530 209144 65006 209250
rect 65174 209144 65650 209250
rect 65818 209144 66294 209250
rect 66462 209144 66938 209250
rect 67106 209144 67582 209250
rect 67750 209144 68226 209250
rect 68394 209144 68870 209250
rect 69038 209144 69514 209250
rect 69682 209144 70158 209250
rect 70326 209144 70802 209250
rect 70970 209144 71446 209250
rect 71614 209144 72090 209250
rect 72258 209144 72734 209250
rect 72902 209144 73378 209250
rect 73546 209144 74022 209250
rect 74190 209144 75310 209250
rect 75478 209144 75954 209250
rect 76122 209144 76598 209250
rect 76766 209144 77242 209250
rect 77410 209144 77886 209250
rect 78054 209144 78530 209250
rect 78698 209144 79174 209250
rect 79342 209144 79818 209250
rect 79986 209144 80462 209250
rect 80630 209144 81106 209250
rect 81274 209144 81750 209250
rect 81918 209144 82394 209250
rect 82562 209144 83038 209250
rect 83206 209144 83682 209250
rect 83850 209144 84326 209250
rect 84494 209144 84970 209250
rect 85138 209144 85614 209250
rect 85782 209144 86258 209250
rect 86426 209144 86902 209250
rect 87070 209144 87546 209250
rect 87714 209144 88190 209250
rect 88358 209144 88834 209250
rect 89002 209144 89478 209250
rect 89646 209144 90122 209250
rect 90290 209144 90766 209250
rect 90934 209144 91410 209250
rect 91578 209144 92054 209250
rect 92222 209144 92698 209250
rect 92866 209144 93342 209250
rect 93510 209144 93986 209250
rect 94154 209144 94630 209250
rect 94798 209144 95274 209250
rect 95442 209144 95918 209250
rect 96086 209144 96562 209250
rect 96730 209144 97850 209250
rect 98018 209144 98494 209250
rect 98662 209144 99138 209250
rect 99306 209144 99782 209250
rect 99950 209144 100426 209250
rect 100594 209144 101070 209250
rect 101238 209144 101714 209250
rect 101882 209144 102358 209250
rect 102526 209144 103002 209250
rect 103170 209144 103646 209250
rect 103814 209144 104290 209250
rect 104458 209144 104934 209250
rect 105102 209144 105578 209250
rect 105746 209144 106222 209250
rect 106390 209144 106866 209250
rect 107034 209144 107510 209250
rect 107678 209144 108154 209250
rect 108322 209144 108798 209250
rect 108966 209144 109442 209250
rect 109610 209144 110086 209250
rect 110254 209144 110730 209250
rect 110898 209144 111374 209250
rect 111542 209144 112018 209250
rect 112186 209144 112662 209250
rect 112830 209144 113306 209250
rect 113474 209144 113950 209250
rect 114118 209144 114594 209250
rect 114762 209144 115238 209250
rect 115406 209144 115882 209250
rect 116050 209144 116526 209250
rect 116694 209144 117170 209250
rect 117338 209144 117814 209250
rect 117982 209144 118458 209250
rect 118626 209144 119102 209250
rect 119270 209144 119856 209250
rect 20 856 119856 209144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 2538 856
rect 2706 31 3182 856
rect 3350 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7046 856
rect 7214 31 7690 856
rect 7858 31 8334 856
rect 8502 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14130 856
rect 14298 31 14774 856
rect 14942 31 15418 856
rect 15586 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17350 856
rect 17518 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 20570 856
rect 20738 31 21214 856
rect 21382 31 21858 856
rect 22026 31 23146 856
rect 23314 31 23790 856
rect 23958 31 24434 856
rect 24602 31 25078 856
rect 25246 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28298 856
rect 28466 31 28942 856
rect 29110 31 29586 856
rect 29754 31 30230 856
rect 30398 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32162 856
rect 32330 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34094 856
rect 34262 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36026 856
rect 36194 31 36670 856
rect 36838 31 37314 856
rect 37482 31 37958 856
rect 38126 31 38602 856
rect 38770 31 39246 856
rect 39414 31 39890 856
rect 40058 31 40534 856
rect 40702 31 41178 856
rect 41346 31 41822 856
rect 41990 31 42466 856
rect 42634 31 43110 856
rect 43278 31 43754 856
rect 43922 31 44398 856
rect 44566 31 45686 856
rect 45854 31 46330 856
rect 46498 31 46974 856
rect 47142 31 47618 856
rect 47786 31 48262 856
rect 48430 31 48906 856
rect 49074 31 49550 856
rect 49718 31 50194 856
rect 50362 31 50838 856
rect 51006 31 51482 856
rect 51650 31 52126 856
rect 52294 31 52770 856
rect 52938 31 53414 856
rect 53582 31 54058 856
rect 54226 31 54702 856
rect 54870 31 55346 856
rect 55514 31 55990 856
rect 56158 31 56634 856
rect 56802 31 57278 856
rect 57446 31 57922 856
rect 58090 31 58566 856
rect 58734 31 59210 856
rect 59378 31 59854 856
rect 60022 31 60498 856
rect 60666 31 61142 856
rect 61310 31 61786 856
rect 61954 31 62430 856
rect 62598 31 63074 856
rect 63242 31 63718 856
rect 63886 31 64362 856
rect 64530 31 65006 856
rect 65174 31 65650 856
rect 65818 31 66294 856
rect 66462 31 66938 856
rect 67106 31 67582 856
rect 67750 31 68870 856
rect 69038 31 69514 856
rect 69682 31 70158 856
rect 70326 31 70802 856
rect 70970 31 71446 856
rect 71614 31 72090 856
rect 72258 31 72734 856
rect 72902 31 73378 856
rect 73546 31 74022 856
rect 74190 31 74666 856
rect 74834 31 75310 856
rect 75478 31 75954 856
rect 76122 31 76598 856
rect 76766 31 77242 856
rect 77410 31 77886 856
rect 78054 31 78530 856
rect 78698 31 79174 856
rect 79342 31 79818 856
rect 79986 31 80462 856
rect 80630 31 81106 856
rect 81274 31 81750 856
rect 81918 31 82394 856
rect 82562 31 83038 856
rect 83206 31 83682 856
rect 83850 31 84326 856
rect 84494 31 84970 856
rect 85138 31 85614 856
rect 85782 31 86258 856
rect 86426 31 86902 856
rect 87070 31 87546 856
rect 87714 31 88190 856
rect 88358 31 88834 856
rect 89002 31 89478 856
rect 89646 31 90122 856
rect 90290 31 91410 856
rect 91578 31 92054 856
rect 92222 31 92698 856
rect 92866 31 93342 856
rect 93510 31 93986 856
rect 94154 31 94630 856
rect 94798 31 95274 856
rect 95442 31 95918 856
rect 96086 31 96562 856
rect 96730 31 97206 856
rect 97374 31 97850 856
rect 98018 31 98494 856
rect 98662 31 99138 856
rect 99306 31 99782 856
rect 99950 31 100426 856
rect 100594 31 101070 856
rect 101238 31 101714 856
rect 101882 31 102358 856
rect 102526 31 103002 856
rect 103170 31 103646 856
rect 103814 31 104290 856
rect 104458 31 104934 856
rect 105102 31 105578 856
rect 105746 31 106222 856
rect 106390 31 106866 856
rect 107034 31 107510 856
rect 107678 31 108154 856
rect 108322 31 108798 856
rect 108966 31 109442 856
rect 109610 31 110086 856
rect 110254 31 110730 856
rect 110898 31 111374 856
rect 111542 31 112018 856
rect 112186 31 112662 856
rect 112830 31 113306 856
rect 113474 31 114594 856
rect 114762 31 115238 856
rect 115406 31 115882 856
rect 116050 31 116526 856
rect 116694 31 117170 856
rect 117338 31 117814 856
rect 117982 31 118458 856
rect 118626 31 119102 856
rect 119270 31 119746 856
<< metal3 >>
rect 0 209448 800 209568
rect 119200 209448 120000 209568
rect 0 208768 800 208888
rect 119200 208768 120000 208888
rect 0 208088 800 208208
rect 119200 208088 120000 208208
rect 0 207408 800 207528
rect 119200 207408 120000 207528
rect 0 206728 800 206848
rect 119200 206728 120000 206848
rect 0 206048 800 206168
rect 119200 206048 120000 206168
rect 0 205368 800 205488
rect 119200 205368 120000 205488
rect 0 204688 800 204808
rect 119200 204688 120000 204808
rect 0 204008 800 204128
rect 119200 204008 120000 204128
rect 0 203328 800 203448
rect 119200 203328 120000 203448
rect 0 202648 800 202768
rect 119200 202648 120000 202768
rect 0 201968 800 202088
rect 119200 201968 120000 202088
rect 0 201288 800 201408
rect 119200 201288 120000 201408
rect 0 200608 800 200728
rect 119200 200608 120000 200728
rect 0 199928 800 200048
rect 119200 199928 120000 200048
rect 0 199248 800 199368
rect 119200 199248 120000 199368
rect 0 198568 800 198688
rect 119200 198568 120000 198688
rect 0 197888 800 198008
rect 119200 197888 120000 198008
rect 0 197208 800 197328
rect 119200 197208 120000 197328
rect 0 196528 800 196648
rect 119200 196528 120000 196648
rect 0 195848 800 195968
rect 119200 195848 120000 195968
rect 0 195168 800 195288
rect 119200 195168 120000 195288
rect 0 194488 800 194608
rect 119200 194488 120000 194608
rect 0 193808 800 193928
rect 119200 193808 120000 193928
rect 0 193128 800 193248
rect 119200 193128 120000 193248
rect 119200 192448 120000 192568
rect 0 191768 800 191888
rect 119200 191768 120000 191888
rect 0 191088 800 191208
rect 119200 191088 120000 191208
rect 0 190408 800 190528
rect 119200 190408 120000 190528
rect 0 189728 800 189848
rect 119200 189728 120000 189848
rect 0 189048 800 189168
rect 119200 189048 120000 189168
rect 0 188368 800 188488
rect 119200 188368 120000 188488
rect 0 187688 800 187808
rect 119200 187688 120000 187808
rect 0 187008 800 187128
rect 119200 187008 120000 187128
rect 0 186328 800 186448
rect 119200 186328 120000 186448
rect 0 185648 800 185768
rect 0 184968 800 185088
rect 119200 184968 120000 185088
rect 0 184288 800 184408
rect 119200 184288 120000 184408
rect 0 183608 800 183728
rect 119200 183608 120000 183728
rect 0 182928 800 183048
rect 119200 182928 120000 183048
rect 0 182248 800 182368
rect 119200 182248 120000 182368
rect 0 181568 800 181688
rect 119200 181568 120000 181688
rect 0 180888 800 181008
rect 119200 180888 120000 181008
rect 0 180208 800 180328
rect 119200 180208 120000 180328
rect 0 179528 800 179648
rect 119200 179528 120000 179648
rect 0 178848 800 178968
rect 119200 178848 120000 178968
rect 0 178168 800 178288
rect 119200 178168 120000 178288
rect 0 177488 800 177608
rect 119200 177488 120000 177608
rect 0 176808 800 176928
rect 119200 176808 120000 176928
rect 0 176128 800 176248
rect 119200 176128 120000 176248
rect 0 175448 800 175568
rect 119200 175448 120000 175568
rect 0 174768 800 174888
rect 119200 174768 120000 174888
rect 0 174088 800 174208
rect 119200 174088 120000 174208
rect 0 173408 800 173528
rect 119200 173408 120000 173528
rect 0 172728 800 172848
rect 119200 172728 120000 172848
rect 0 172048 800 172168
rect 119200 172048 120000 172168
rect 0 171368 800 171488
rect 119200 171368 120000 171488
rect 0 170688 800 170808
rect 119200 170688 120000 170808
rect 0 170008 800 170128
rect 119200 170008 120000 170128
rect 0 169328 800 169448
rect 119200 169328 120000 169448
rect 0 168648 800 168768
rect 119200 168648 120000 168768
rect 119200 167968 120000 168088
rect 0 167288 800 167408
rect 119200 167288 120000 167408
rect 0 166608 800 166728
rect 119200 166608 120000 166728
rect 0 165928 800 166048
rect 119200 165928 120000 166048
rect 0 165248 800 165368
rect 119200 165248 120000 165368
rect 0 164568 800 164688
rect 119200 164568 120000 164688
rect 0 163888 800 164008
rect 119200 163888 120000 164008
rect 0 163208 800 163328
rect 119200 163208 120000 163328
rect 0 162528 800 162648
rect 119200 162528 120000 162648
rect 0 161848 800 161968
rect 0 161168 800 161288
rect 119200 161168 120000 161288
rect 0 160488 800 160608
rect 119200 160488 120000 160608
rect 0 159808 800 159928
rect 119200 159808 120000 159928
rect 0 159128 800 159248
rect 119200 159128 120000 159248
rect 0 158448 800 158568
rect 119200 158448 120000 158568
rect 0 157768 800 157888
rect 119200 157768 120000 157888
rect 0 157088 800 157208
rect 119200 157088 120000 157208
rect 0 156408 800 156528
rect 119200 156408 120000 156528
rect 0 155728 800 155848
rect 119200 155728 120000 155848
rect 0 155048 800 155168
rect 119200 155048 120000 155168
rect 0 154368 800 154488
rect 119200 154368 120000 154488
rect 0 153688 800 153808
rect 119200 153688 120000 153808
rect 0 153008 800 153128
rect 119200 153008 120000 153128
rect 0 152328 800 152448
rect 119200 152328 120000 152448
rect 0 151648 800 151768
rect 119200 151648 120000 151768
rect 0 150968 800 151088
rect 119200 150968 120000 151088
rect 0 150288 800 150408
rect 119200 150288 120000 150408
rect 0 149608 800 149728
rect 119200 149608 120000 149728
rect 0 148928 800 149048
rect 119200 148928 120000 149048
rect 0 148248 800 148368
rect 119200 148248 120000 148368
rect 0 147568 800 147688
rect 119200 147568 120000 147688
rect 0 146888 800 147008
rect 119200 146888 120000 147008
rect 0 146208 800 146328
rect 119200 146208 120000 146328
rect 0 145528 800 145648
rect 119200 145528 120000 145648
rect 0 144848 800 144968
rect 119200 144848 120000 144968
rect 119200 144168 120000 144288
rect 0 143488 800 143608
rect 119200 143488 120000 143608
rect 0 142808 800 142928
rect 119200 142808 120000 142928
rect 0 142128 800 142248
rect 119200 142128 120000 142248
rect 0 141448 800 141568
rect 119200 141448 120000 141568
rect 0 140768 800 140888
rect 119200 140768 120000 140888
rect 0 140088 800 140208
rect 119200 140088 120000 140208
rect 0 139408 800 139528
rect 119200 139408 120000 139528
rect 0 138728 800 138848
rect 119200 138728 120000 138848
rect 0 138048 800 138168
rect 119200 138048 120000 138168
rect 0 137368 800 137488
rect 0 136688 800 136808
rect 119200 136688 120000 136808
rect 0 136008 800 136128
rect 119200 136008 120000 136128
rect 0 135328 800 135448
rect 119200 135328 120000 135448
rect 0 134648 800 134768
rect 119200 134648 120000 134768
rect 0 133968 800 134088
rect 119200 133968 120000 134088
rect 0 133288 800 133408
rect 119200 133288 120000 133408
rect 0 132608 800 132728
rect 119200 132608 120000 132728
rect 0 131928 800 132048
rect 119200 131928 120000 132048
rect 0 131248 800 131368
rect 119200 131248 120000 131368
rect 0 130568 800 130688
rect 119200 130568 120000 130688
rect 0 129888 800 130008
rect 119200 129888 120000 130008
rect 0 129208 800 129328
rect 119200 129208 120000 129328
rect 0 128528 800 128648
rect 119200 128528 120000 128648
rect 0 127848 800 127968
rect 119200 127848 120000 127968
rect 0 127168 800 127288
rect 119200 127168 120000 127288
rect 0 126488 800 126608
rect 119200 126488 120000 126608
rect 0 125808 800 125928
rect 119200 125808 120000 125928
rect 0 125128 800 125248
rect 119200 125128 120000 125248
rect 0 124448 800 124568
rect 119200 124448 120000 124568
rect 0 123768 800 123888
rect 119200 123768 120000 123888
rect 0 123088 800 123208
rect 119200 123088 120000 123208
rect 0 122408 800 122528
rect 119200 122408 120000 122528
rect 0 121728 800 121848
rect 119200 121728 120000 121848
rect 0 121048 800 121168
rect 119200 121048 120000 121168
rect 119200 120368 120000 120488
rect 0 119688 800 119808
rect 119200 119688 120000 119808
rect 0 119008 800 119128
rect 119200 119008 120000 119128
rect 0 118328 800 118448
rect 119200 118328 120000 118448
rect 0 117648 800 117768
rect 119200 117648 120000 117768
rect 0 116968 800 117088
rect 119200 116968 120000 117088
rect 0 116288 800 116408
rect 119200 116288 120000 116408
rect 0 115608 800 115728
rect 119200 115608 120000 115728
rect 0 114928 800 115048
rect 119200 114928 120000 115048
rect 0 114248 800 114368
rect 119200 114248 120000 114368
rect 0 113568 800 113688
rect 0 112888 800 113008
rect 119200 112888 120000 113008
rect 0 112208 800 112328
rect 119200 112208 120000 112328
rect 0 111528 800 111648
rect 119200 111528 120000 111648
rect 0 110848 800 110968
rect 119200 110848 120000 110968
rect 0 110168 800 110288
rect 119200 110168 120000 110288
rect 0 109488 800 109608
rect 119200 109488 120000 109608
rect 0 108808 800 108928
rect 119200 108808 120000 108928
rect 0 108128 800 108248
rect 119200 108128 120000 108248
rect 0 107448 800 107568
rect 119200 107448 120000 107568
rect 0 106768 800 106888
rect 119200 106768 120000 106888
rect 0 106088 800 106208
rect 119200 106088 120000 106208
rect 0 105408 800 105528
rect 119200 105408 120000 105528
rect 0 104728 800 104848
rect 119200 104728 120000 104848
rect 0 104048 800 104168
rect 119200 104048 120000 104168
rect 0 103368 800 103488
rect 119200 103368 120000 103488
rect 0 102688 800 102808
rect 119200 102688 120000 102808
rect 0 102008 800 102128
rect 119200 102008 120000 102128
rect 0 101328 800 101448
rect 119200 101328 120000 101448
rect 0 100648 800 100768
rect 119200 100648 120000 100768
rect 0 99968 800 100088
rect 119200 99968 120000 100088
rect 0 99288 800 99408
rect 119200 99288 120000 99408
rect 0 98608 800 98728
rect 119200 98608 120000 98728
rect 0 97928 800 98048
rect 119200 97928 120000 98048
rect 0 97248 800 97368
rect 119200 97248 120000 97368
rect 0 96568 800 96688
rect 119200 96568 120000 96688
rect 119200 95888 120000 96008
rect 0 95208 800 95328
rect 119200 95208 120000 95328
rect 0 94528 800 94648
rect 119200 94528 120000 94648
rect 0 93848 800 93968
rect 119200 93848 120000 93968
rect 0 93168 800 93288
rect 119200 93168 120000 93288
rect 0 92488 800 92608
rect 119200 92488 120000 92608
rect 0 91808 800 91928
rect 119200 91808 120000 91928
rect 0 91128 800 91248
rect 119200 91128 120000 91248
rect 0 90448 800 90568
rect 119200 90448 120000 90568
rect 0 89768 800 89888
rect 119200 89768 120000 89888
rect 0 89088 800 89208
rect 0 88408 800 88528
rect 119200 88408 120000 88528
rect 0 87728 800 87848
rect 119200 87728 120000 87848
rect 0 87048 800 87168
rect 119200 87048 120000 87168
rect 0 86368 800 86488
rect 119200 86368 120000 86488
rect 0 85688 800 85808
rect 119200 85688 120000 85808
rect 0 85008 800 85128
rect 119200 85008 120000 85128
rect 0 84328 800 84448
rect 119200 84328 120000 84448
rect 0 83648 800 83768
rect 119200 83648 120000 83768
rect 0 82968 800 83088
rect 119200 82968 120000 83088
rect 0 82288 800 82408
rect 119200 82288 120000 82408
rect 0 81608 800 81728
rect 119200 81608 120000 81728
rect 0 80928 800 81048
rect 119200 80928 120000 81048
rect 0 80248 800 80368
rect 119200 80248 120000 80368
rect 0 79568 800 79688
rect 119200 79568 120000 79688
rect 0 78888 800 79008
rect 119200 78888 120000 79008
rect 0 78208 800 78328
rect 119200 78208 120000 78328
rect 0 77528 800 77648
rect 119200 77528 120000 77648
rect 0 76848 800 76968
rect 119200 76848 120000 76968
rect 0 76168 800 76288
rect 119200 76168 120000 76288
rect 0 75488 800 75608
rect 119200 75488 120000 75608
rect 0 74808 800 74928
rect 119200 74808 120000 74928
rect 0 74128 800 74248
rect 119200 74128 120000 74248
rect 0 73448 800 73568
rect 119200 73448 120000 73568
rect 0 72768 800 72888
rect 119200 72768 120000 72888
rect 119200 72088 120000 72208
rect 0 71408 800 71528
rect 119200 71408 120000 71528
rect 0 70728 800 70848
rect 119200 70728 120000 70848
rect 0 70048 800 70168
rect 119200 70048 120000 70168
rect 0 69368 800 69488
rect 119200 69368 120000 69488
rect 0 68688 800 68808
rect 119200 68688 120000 68808
rect 0 68008 800 68128
rect 119200 68008 120000 68128
rect 0 67328 800 67448
rect 119200 67328 120000 67448
rect 0 66648 800 66768
rect 119200 66648 120000 66768
rect 0 65968 800 66088
rect 119200 65968 120000 66088
rect 0 65288 800 65408
rect 0 64608 800 64728
rect 119200 64608 120000 64728
rect 0 63928 800 64048
rect 119200 63928 120000 64048
rect 0 63248 800 63368
rect 119200 63248 120000 63368
rect 0 62568 800 62688
rect 119200 62568 120000 62688
rect 0 61888 800 62008
rect 119200 61888 120000 62008
rect 0 61208 800 61328
rect 119200 61208 120000 61328
rect 0 60528 800 60648
rect 119200 60528 120000 60648
rect 0 59848 800 59968
rect 119200 59848 120000 59968
rect 0 59168 800 59288
rect 119200 59168 120000 59288
rect 0 58488 800 58608
rect 119200 58488 120000 58608
rect 0 57808 800 57928
rect 119200 57808 120000 57928
rect 0 57128 800 57248
rect 119200 57128 120000 57248
rect 0 56448 800 56568
rect 119200 56448 120000 56568
rect 0 55768 800 55888
rect 119200 55768 120000 55888
rect 0 55088 800 55208
rect 119200 55088 120000 55208
rect 0 54408 800 54528
rect 119200 54408 120000 54528
rect 0 53728 800 53848
rect 119200 53728 120000 53848
rect 0 53048 800 53168
rect 119200 53048 120000 53168
rect 0 52368 800 52488
rect 119200 52368 120000 52488
rect 0 51688 800 51808
rect 119200 51688 120000 51808
rect 0 51008 800 51128
rect 119200 51008 120000 51128
rect 0 50328 800 50448
rect 119200 50328 120000 50448
rect 0 49648 800 49768
rect 119200 49648 120000 49768
rect 0 48968 800 49088
rect 119200 48968 120000 49088
rect 0 48288 800 48408
rect 119200 48288 120000 48408
rect 119200 47608 120000 47728
rect 0 46928 800 47048
rect 119200 46928 120000 47048
rect 0 46248 800 46368
rect 119200 46248 120000 46368
rect 0 45568 800 45688
rect 119200 45568 120000 45688
rect 0 44888 800 45008
rect 119200 44888 120000 45008
rect 0 44208 800 44328
rect 119200 44208 120000 44328
rect 0 43528 800 43648
rect 119200 43528 120000 43648
rect 0 42848 800 42968
rect 119200 42848 120000 42968
rect 0 42168 800 42288
rect 119200 42168 120000 42288
rect 0 41488 800 41608
rect 0 40808 800 40928
rect 119200 40808 120000 40928
rect 0 40128 800 40248
rect 119200 40128 120000 40248
rect 0 39448 800 39568
rect 119200 39448 120000 39568
rect 0 38768 800 38888
rect 119200 38768 120000 38888
rect 0 38088 800 38208
rect 119200 38088 120000 38208
rect 0 37408 800 37528
rect 119200 37408 120000 37528
rect 0 36728 800 36848
rect 119200 36728 120000 36848
rect 0 36048 800 36168
rect 119200 36048 120000 36168
rect 0 35368 800 35488
rect 119200 35368 120000 35488
rect 0 34688 800 34808
rect 119200 34688 120000 34808
rect 0 34008 800 34128
rect 119200 34008 120000 34128
rect 0 33328 800 33448
rect 119200 33328 120000 33448
rect 0 32648 800 32768
rect 119200 32648 120000 32768
rect 0 31968 800 32088
rect 119200 31968 120000 32088
rect 0 31288 800 31408
rect 119200 31288 120000 31408
rect 0 30608 800 30728
rect 119200 30608 120000 30728
rect 0 29928 800 30048
rect 119200 29928 120000 30048
rect 0 29248 800 29368
rect 119200 29248 120000 29368
rect 0 28568 800 28688
rect 119200 28568 120000 28688
rect 0 27888 800 28008
rect 119200 27888 120000 28008
rect 0 27208 800 27328
rect 119200 27208 120000 27328
rect 0 26528 800 26648
rect 119200 26528 120000 26648
rect 0 25848 800 25968
rect 119200 25848 120000 25968
rect 0 25168 800 25288
rect 119200 25168 120000 25288
rect 0 24488 800 24608
rect 119200 24488 120000 24608
rect 119200 23808 120000 23928
rect 0 23128 800 23248
rect 119200 23128 120000 23248
rect 0 22448 800 22568
rect 119200 22448 120000 22568
rect 0 21768 800 21888
rect 119200 21768 120000 21888
rect 0 21088 800 21208
rect 119200 21088 120000 21208
rect 0 20408 800 20528
rect 119200 20408 120000 20528
rect 0 19728 800 19848
rect 119200 19728 120000 19848
rect 0 19048 800 19168
rect 119200 19048 120000 19168
rect 0 18368 800 18488
rect 119200 18368 120000 18488
rect 0 17688 800 17808
rect 119200 17688 120000 17808
rect 0 17008 800 17128
rect 0 16328 800 16448
rect 119200 16328 120000 16448
rect 0 15648 800 15768
rect 119200 15648 120000 15768
rect 0 14968 800 15088
rect 119200 14968 120000 15088
rect 0 14288 800 14408
rect 119200 14288 120000 14408
rect 0 13608 800 13728
rect 119200 13608 120000 13728
rect 0 12928 800 13048
rect 119200 12928 120000 13048
rect 0 12248 800 12368
rect 119200 12248 120000 12368
rect 0 11568 800 11688
rect 119200 11568 120000 11688
rect 0 10888 800 11008
rect 119200 10888 120000 11008
rect 0 10208 800 10328
rect 119200 10208 120000 10328
rect 0 9528 800 9648
rect 119200 9528 120000 9648
rect 0 8848 800 8968
rect 119200 8848 120000 8968
rect 0 8168 800 8288
rect 119200 8168 120000 8288
rect 0 7488 800 7608
rect 119200 7488 120000 7608
rect 0 6808 800 6928
rect 119200 6808 120000 6928
rect 0 6128 800 6248
rect 119200 6128 120000 6248
rect 0 5448 800 5568
rect 119200 5448 120000 5568
rect 0 4768 800 4888
rect 119200 4768 120000 4888
rect 0 4088 800 4208
rect 119200 4088 120000 4208
rect 0 3408 800 3528
rect 119200 3408 120000 3528
rect 0 2728 800 2848
rect 119200 2728 120000 2848
rect 0 2048 800 2168
rect 119200 2048 120000 2168
rect 0 1368 800 1488
rect 119200 1368 120000 1488
rect 0 688 800 808
rect 119200 688 120000 808
rect 119200 8 120000 128
<< obsm3 >>
rect 880 208688 119120 208861
rect 800 208288 119200 208688
rect 880 208008 119120 208288
rect 800 207608 119200 208008
rect 880 207328 119120 207608
rect 800 206928 119200 207328
rect 880 206648 119120 206928
rect 800 206248 119200 206648
rect 880 205968 119120 206248
rect 800 205568 119200 205968
rect 880 205288 119120 205568
rect 800 204888 119200 205288
rect 880 204608 119120 204888
rect 800 204208 119200 204608
rect 880 203928 119120 204208
rect 800 203528 119200 203928
rect 880 203248 119120 203528
rect 800 202848 119200 203248
rect 880 202568 119120 202848
rect 800 202168 119200 202568
rect 880 201888 119120 202168
rect 800 201488 119200 201888
rect 880 201208 119120 201488
rect 800 200808 119200 201208
rect 880 200528 119120 200808
rect 800 200128 119200 200528
rect 880 199848 119120 200128
rect 800 199448 119200 199848
rect 880 199168 119120 199448
rect 800 198768 119200 199168
rect 880 198488 119120 198768
rect 800 198088 119200 198488
rect 880 197808 119120 198088
rect 800 197408 119200 197808
rect 880 197128 119120 197408
rect 800 196728 119200 197128
rect 880 196448 119120 196728
rect 800 196048 119200 196448
rect 880 195768 119120 196048
rect 800 195368 119200 195768
rect 880 195088 119120 195368
rect 800 194688 119200 195088
rect 880 194408 119120 194688
rect 800 194008 119200 194408
rect 880 193728 119120 194008
rect 800 193328 119200 193728
rect 880 193048 119120 193328
rect 800 192648 119200 193048
rect 800 192368 119120 192648
rect 800 191968 119200 192368
rect 880 191688 119120 191968
rect 800 191288 119200 191688
rect 880 191008 119120 191288
rect 800 190608 119200 191008
rect 880 190328 119120 190608
rect 800 189928 119200 190328
rect 880 189648 119120 189928
rect 800 189248 119200 189648
rect 880 188968 119120 189248
rect 800 188568 119200 188968
rect 880 188288 119120 188568
rect 800 187888 119200 188288
rect 880 187608 119120 187888
rect 800 187208 119200 187608
rect 880 186928 119120 187208
rect 800 186528 119200 186928
rect 880 186248 119120 186528
rect 800 185848 119200 186248
rect 880 185568 119200 185848
rect 800 185168 119200 185568
rect 880 184888 119120 185168
rect 800 184488 119200 184888
rect 880 184208 119120 184488
rect 800 183808 119200 184208
rect 880 183528 119120 183808
rect 800 183128 119200 183528
rect 880 182848 119120 183128
rect 800 182448 119200 182848
rect 880 182168 119120 182448
rect 800 181768 119200 182168
rect 880 181488 119120 181768
rect 800 181088 119200 181488
rect 880 180808 119120 181088
rect 800 180408 119200 180808
rect 880 180128 119120 180408
rect 800 179728 119200 180128
rect 880 179448 119120 179728
rect 800 179048 119200 179448
rect 880 178768 119120 179048
rect 800 178368 119200 178768
rect 880 178088 119120 178368
rect 800 177688 119200 178088
rect 880 177408 119120 177688
rect 800 177008 119200 177408
rect 880 176728 119120 177008
rect 800 176328 119200 176728
rect 880 176048 119120 176328
rect 800 175648 119200 176048
rect 880 175368 119120 175648
rect 800 174968 119200 175368
rect 880 174688 119120 174968
rect 800 174288 119200 174688
rect 880 174008 119120 174288
rect 800 173608 119200 174008
rect 880 173328 119120 173608
rect 800 172928 119200 173328
rect 880 172648 119120 172928
rect 800 172248 119200 172648
rect 880 171968 119120 172248
rect 800 171568 119200 171968
rect 880 171288 119120 171568
rect 800 170888 119200 171288
rect 880 170608 119120 170888
rect 800 170208 119200 170608
rect 880 169928 119120 170208
rect 800 169528 119200 169928
rect 880 169248 119120 169528
rect 800 168848 119200 169248
rect 880 168568 119120 168848
rect 800 168168 119200 168568
rect 800 167888 119120 168168
rect 800 167488 119200 167888
rect 880 167208 119120 167488
rect 800 166808 119200 167208
rect 880 166528 119120 166808
rect 800 166128 119200 166528
rect 880 165848 119120 166128
rect 800 165448 119200 165848
rect 880 165168 119120 165448
rect 800 164768 119200 165168
rect 880 164488 119120 164768
rect 800 164088 119200 164488
rect 880 163808 119120 164088
rect 800 163408 119200 163808
rect 880 163128 119120 163408
rect 800 162728 119200 163128
rect 880 162448 119120 162728
rect 800 162048 119200 162448
rect 880 161768 119200 162048
rect 800 161368 119200 161768
rect 880 161088 119120 161368
rect 800 160688 119200 161088
rect 880 160408 119120 160688
rect 800 160008 119200 160408
rect 880 159728 119120 160008
rect 800 159328 119200 159728
rect 880 159048 119120 159328
rect 800 158648 119200 159048
rect 880 158368 119120 158648
rect 800 157968 119200 158368
rect 880 157688 119120 157968
rect 800 157288 119200 157688
rect 880 157008 119120 157288
rect 800 156608 119200 157008
rect 880 156328 119120 156608
rect 800 155928 119200 156328
rect 880 155648 119120 155928
rect 800 155248 119200 155648
rect 880 154968 119120 155248
rect 800 154568 119200 154968
rect 880 154288 119120 154568
rect 800 153888 119200 154288
rect 880 153608 119120 153888
rect 800 153208 119200 153608
rect 880 152928 119120 153208
rect 800 152528 119200 152928
rect 880 152248 119120 152528
rect 800 151848 119200 152248
rect 880 151568 119120 151848
rect 800 151168 119200 151568
rect 880 150888 119120 151168
rect 800 150488 119200 150888
rect 880 150208 119120 150488
rect 800 149808 119200 150208
rect 880 149528 119120 149808
rect 800 149128 119200 149528
rect 880 148848 119120 149128
rect 800 148448 119200 148848
rect 880 148168 119120 148448
rect 800 147768 119200 148168
rect 880 147488 119120 147768
rect 800 147088 119200 147488
rect 880 146808 119120 147088
rect 800 146408 119200 146808
rect 880 146128 119120 146408
rect 800 145728 119200 146128
rect 880 145448 119120 145728
rect 800 145048 119200 145448
rect 880 144768 119120 145048
rect 800 144368 119200 144768
rect 800 144088 119120 144368
rect 800 143688 119200 144088
rect 880 143408 119120 143688
rect 800 143008 119200 143408
rect 880 142728 119120 143008
rect 800 142328 119200 142728
rect 880 142048 119120 142328
rect 800 141648 119200 142048
rect 880 141368 119120 141648
rect 800 140968 119200 141368
rect 880 140688 119120 140968
rect 800 140288 119200 140688
rect 880 140008 119120 140288
rect 800 139608 119200 140008
rect 880 139328 119120 139608
rect 800 138928 119200 139328
rect 880 138648 119120 138928
rect 800 138248 119200 138648
rect 880 137968 119120 138248
rect 800 137568 119200 137968
rect 880 137288 119200 137568
rect 800 136888 119200 137288
rect 880 136608 119120 136888
rect 800 136208 119200 136608
rect 880 135928 119120 136208
rect 800 135528 119200 135928
rect 880 135248 119120 135528
rect 800 134848 119200 135248
rect 880 134568 119120 134848
rect 800 134168 119200 134568
rect 880 133888 119120 134168
rect 800 133488 119200 133888
rect 880 133208 119120 133488
rect 800 132808 119200 133208
rect 880 132528 119120 132808
rect 800 132128 119200 132528
rect 880 131848 119120 132128
rect 800 131448 119200 131848
rect 880 131168 119120 131448
rect 800 130768 119200 131168
rect 880 130488 119120 130768
rect 800 130088 119200 130488
rect 880 129808 119120 130088
rect 800 129408 119200 129808
rect 880 129128 119120 129408
rect 800 128728 119200 129128
rect 880 128448 119120 128728
rect 800 128048 119200 128448
rect 880 127768 119120 128048
rect 800 127368 119200 127768
rect 880 127088 119120 127368
rect 800 126688 119200 127088
rect 880 126408 119120 126688
rect 800 126008 119200 126408
rect 880 125728 119120 126008
rect 800 125328 119200 125728
rect 880 125048 119120 125328
rect 800 124648 119200 125048
rect 880 124368 119120 124648
rect 800 123968 119200 124368
rect 880 123688 119120 123968
rect 800 123288 119200 123688
rect 880 123008 119120 123288
rect 800 122608 119200 123008
rect 880 122328 119120 122608
rect 800 121928 119200 122328
rect 880 121648 119120 121928
rect 800 121248 119200 121648
rect 880 120968 119120 121248
rect 800 120568 119200 120968
rect 800 120288 119120 120568
rect 800 119888 119200 120288
rect 880 119608 119120 119888
rect 800 119208 119200 119608
rect 880 118928 119120 119208
rect 800 118528 119200 118928
rect 880 118248 119120 118528
rect 800 117848 119200 118248
rect 880 117568 119120 117848
rect 800 117168 119200 117568
rect 880 116888 119120 117168
rect 800 116488 119200 116888
rect 880 116208 119120 116488
rect 800 115808 119200 116208
rect 880 115528 119120 115808
rect 800 115128 119200 115528
rect 880 114848 119120 115128
rect 800 114448 119200 114848
rect 880 114168 119120 114448
rect 800 113768 119200 114168
rect 880 113488 119200 113768
rect 800 113088 119200 113488
rect 880 112808 119120 113088
rect 800 112408 119200 112808
rect 880 112128 119120 112408
rect 800 111728 119200 112128
rect 880 111448 119120 111728
rect 800 111048 119200 111448
rect 880 110768 119120 111048
rect 800 110368 119200 110768
rect 880 110088 119120 110368
rect 800 109688 119200 110088
rect 880 109408 119120 109688
rect 800 109008 119200 109408
rect 880 108728 119120 109008
rect 800 108328 119200 108728
rect 880 108048 119120 108328
rect 800 107648 119200 108048
rect 880 107368 119120 107648
rect 800 106968 119200 107368
rect 880 106688 119120 106968
rect 800 106288 119200 106688
rect 880 106008 119120 106288
rect 800 105608 119200 106008
rect 880 105328 119120 105608
rect 800 104928 119200 105328
rect 880 104648 119120 104928
rect 800 104248 119200 104648
rect 880 103968 119120 104248
rect 800 103568 119200 103968
rect 880 103288 119120 103568
rect 800 102888 119200 103288
rect 880 102608 119120 102888
rect 800 102208 119200 102608
rect 880 101928 119120 102208
rect 800 101528 119200 101928
rect 880 101248 119120 101528
rect 800 100848 119200 101248
rect 880 100568 119120 100848
rect 800 100168 119200 100568
rect 880 99888 119120 100168
rect 800 99488 119200 99888
rect 880 99208 119120 99488
rect 800 98808 119200 99208
rect 880 98528 119120 98808
rect 800 98128 119200 98528
rect 880 97848 119120 98128
rect 800 97448 119200 97848
rect 880 97168 119120 97448
rect 800 96768 119200 97168
rect 880 96488 119120 96768
rect 800 96088 119200 96488
rect 800 95808 119120 96088
rect 800 95408 119200 95808
rect 880 95128 119120 95408
rect 800 94728 119200 95128
rect 880 94448 119120 94728
rect 800 94048 119200 94448
rect 880 93768 119120 94048
rect 800 93368 119200 93768
rect 880 93088 119120 93368
rect 800 92688 119200 93088
rect 880 92408 119120 92688
rect 800 92008 119200 92408
rect 880 91728 119120 92008
rect 800 91328 119200 91728
rect 880 91048 119120 91328
rect 800 90648 119200 91048
rect 880 90368 119120 90648
rect 800 89968 119200 90368
rect 880 89688 119120 89968
rect 800 89288 119200 89688
rect 880 89008 119200 89288
rect 800 88608 119200 89008
rect 880 88328 119120 88608
rect 800 87928 119200 88328
rect 880 87648 119120 87928
rect 800 87248 119200 87648
rect 880 86968 119120 87248
rect 800 86568 119200 86968
rect 880 86288 119120 86568
rect 800 85888 119200 86288
rect 880 85608 119120 85888
rect 800 85208 119200 85608
rect 880 84928 119120 85208
rect 800 84528 119200 84928
rect 880 84248 119120 84528
rect 800 83848 119200 84248
rect 880 83568 119120 83848
rect 800 83168 119200 83568
rect 880 82888 119120 83168
rect 800 82488 119200 82888
rect 880 82208 119120 82488
rect 800 81808 119200 82208
rect 880 81528 119120 81808
rect 800 81128 119200 81528
rect 880 80848 119120 81128
rect 800 80448 119200 80848
rect 880 80168 119120 80448
rect 800 79768 119200 80168
rect 880 79488 119120 79768
rect 800 79088 119200 79488
rect 880 78808 119120 79088
rect 800 78408 119200 78808
rect 880 78128 119120 78408
rect 800 77728 119200 78128
rect 880 77448 119120 77728
rect 800 77048 119200 77448
rect 880 76768 119120 77048
rect 800 76368 119200 76768
rect 880 76088 119120 76368
rect 800 75688 119200 76088
rect 880 75408 119120 75688
rect 800 75008 119200 75408
rect 880 74728 119120 75008
rect 800 74328 119200 74728
rect 880 74048 119120 74328
rect 800 73648 119200 74048
rect 880 73368 119120 73648
rect 800 72968 119200 73368
rect 880 72688 119120 72968
rect 800 72288 119200 72688
rect 800 72008 119120 72288
rect 800 71608 119200 72008
rect 880 71328 119120 71608
rect 800 70928 119200 71328
rect 880 70648 119120 70928
rect 800 70248 119200 70648
rect 880 69968 119120 70248
rect 800 69568 119200 69968
rect 880 69288 119120 69568
rect 800 68888 119200 69288
rect 880 68608 119120 68888
rect 800 68208 119200 68608
rect 880 67928 119120 68208
rect 800 67528 119200 67928
rect 880 67248 119120 67528
rect 800 66848 119200 67248
rect 880 66568 119120 66848
rect 800 66168 119200 66568
rect 880 65888 119120 66168
rect 800 65488 119200 65888
rect 880 65208 119200 65488
rect 800 64808 119200 65208
rect 880 64528 119120 64808
rect 800 64128 119200 64528
rect 880 63848 119120 64128
rect 800 63448 119200 63848
rect 880 63168 119120 63448
rect 800 62768 119200 63168
rect 880 62488 119120 62768
rect 800 62088 119200 62488
rect 880 61808 119120 62088
rect 800 61408 119200 61808
rect 880 61128 119120 61408
rect 800 60728 119200 61128
rect 880 60448 119120 60728
rect 800 60048 119200 60448
rect 880 59768 119120 60048
rect 800 59368 119200 59768
rect 880 59088 119120 59368
rect 800 58688 119200 59088
rect 880 58408 119120 58688
rect 800 58008 119200 58408
rect 880 57728 119120 58008
rect 800 57328 119200 57728
rect 880 57048 119120 57328
rect 800 56648 119200 57048
rect 880 56368 119120 56648
rect 800 55968 119200 56368
rect 880 55688 119120 55968
rect 800 55288 119200 55688
rect 880 55008 119120 55288
rect 800 54608 119200 55008
rect 880 54328 119120 54608
rect 800 53928 119200 54328
rect 880 53648 119120 53928
rect 800 53248 119200 53648
rect 880 52968 119120 53248
rect 800 52568 119200 52968
rect 880 52288 119120 52568
rect 800 51888 119200 52288
rect 880 51608 119120 51888
rect 800 51208 119200 51608
rect 880 50928 119120 51208
rect 800 50528 119200 50928
rect 880 50248 119120 50528
rect 800 49848 119200 50248
rect 880 49568 119120 49848
rect 800 49168 119200 49568
rect 880 48888 119120 49168
rect 800 48488 119200 48888
rect 880 48208 119120 48488
rect 800 47808 119200 48208
rect 800 47528 119120 47808
rect 800 47128 119200 47528
rect 880 46848 119120 47128
rect 800 46448 119200 46848
rect 880 46168 119120 46448
rect 800 45768 119200 46168
rect 880 45488 119120 45768
rect 800 45088 119200 45488
rect 880 44808 119120 45088
rect 800 44408 119200 44808
rect 880 44128 119120 44408
rect 800 43728 119200 44128
rect 880 43448 119120 43728
rect 800 43048 119200 43448
rect 880 42768 119120 43048
rect 800 42368 119200 42768
rect 880 42088 119120 42368
rect 800 41688 119200 42088
rect 880 41408 119200 41688
rect 800 41008 119200 41408
rect 880 40728 119120 41008
rect 800 40328 119200 40728
rect 880 40048 119120 40328
rect 800 39648 119200 40048
rect 880 39368 119120 39648
rect 800 38968 119200 39368
rect 880 38688 119120 38968
rect 800 38288 119200 38688
rect 880 38008 119120 38288
rect 800 37608 119200 38008
rect 880 37328 119120 37608
rect 800 36928 119200 37328
rect 880 36648 119120 36928
rect 800 36248 119200 36648
rect 880 35968 119120 36248
rect 800 35568 119200 35968
rect 880 35288 119120 35568
rect 800 34888 119200 35288
rect 880 34608 119120 34888
rect 800 34208 119200 34608
rect 880 33928 119120 34208
rect 800 33528 119200 33928
rect 880 33248 119120 33528
rect 800 32848 119200 33248
rect 880 32568 119120 32848
rect 800 32168 119200 32568
rect 880 31888 119120 32168
rect 800 31488 119200 31888
rect 880 31208 119120 31488
rect 800 30808 119200 31208
rect 880 30528 119120 30808
rect 800 30128 119200 30528
rect 880 29848 119120 30128
rect 800 29448 119200 29848
rect 880 29168 119120 29448
rect 800 28768 119200 29168
rect 880 28488 119120 28768
rect 800 28088 119200 28488
rect 880 27808 119120 28088
rect 800 27408 119200 27808
rect 880 27128 119120 27408
rect 800 26728 119200 27128
rect 880 26448 119120 26728
rect 800 26048 119200 26448
rect 880 25768 119120 26048
rect 800 25368 119200 25768
rect 880 25088 119120 25368
rect 800 24688 119200 25088
rect 880 24408 119120 24688
rect 800 24008 119200 24408
rect 800 23728 119120 24008
rect 800 23328 119200 23728
rect 880 23048 119120 23328
rect 800 22648 119200 23048
rect 880 22368 119120 22648
rect 800 21968 119200 22368
rect 880 21688 119120 21968
rect 800 21288 119200 21688
rect 880 21008 119120 21288
rect 800 20608 119200 21008
rect 880 20328 119120 20608
rect 800 19928 119200 20328
rect 880 19648 119120 19928
rect 800 19248 119200 19648
rect 880 18968 119120 19248
rect 800 18568 119200 18968
rect 880 18288 119120 18568
rect 800 17888 119200 18288
rect 880 17608 119120 17888
rect 800 17208 119200 17608
rect 880 16928 119200 17208
rect 800 16528 119200 16928
rect 880 16248 119120 16528
rect 800 15848 119200 16248
rect 880 15568 119120 15848
rect 800 15168 119200 15568
rect 880 14888 119120 15168
rect 800 14488 119200 14888
rect 880 14208 119120 14488
rect 800 13808 119200 14208
rect 880 13528 119120 13808
rect 800 13128 119200 13528
rect 880 12848 119120 13128
rect 800 12448 119200 12848
rect 880 12168 119120 12448
rect 800 11768 119200 12168
rect 880 11488 119120 11768
rect 800 11088 119200 11488
rect 880 10808 119120 11088
rect 800 10408 119200 10808
rect 880 10128 119120 10408
rect 800 9728 119200 10128
rect 880 9448 119120 9728
rect 800 9048 119200 9448
rect 880 8768 119120 9048
rect 800 8368 119200 8768
rect 880 8088 119120 8368
rect 800 7688 119200 8088
rect 880 7408 119120 7688
rect 800 7008 119200 7408
rect 880 6728 119120 7008
rect 800 6328 119200 6728
rect 880 6048 119120 6328
rect 800 5648 119200 6048
rect 880 5368 119120 5648
rect 800 4968 119200 5368
rect 880 4688 119120 4968
rect 800 4288 119200 4688
rect 880 4008 119120 4288
rect 800 3608 119200 4008
rect 880 3328 119120 3608
rect 800 2928 119200 3328
rect 880 2648 119120 2928
rect 800 2248 119200 2648
rect 880 1968 119120 2248
rect 800 1568 119200 1968
rect 880 1288 119120 1568
rect 800 888 119200 1288
rect 880 608 119120 888
rect 800 208 119200 608
rect 800 35 119120 208
<< metal4 >>
rect 4208 2128 4528 207856
rect 19568 2128 19888 207856
rect 34928 2128 35248 207856
rect 50288 2128 50608 207856
rect 65648 2128 65968 207856
rect 81008 2128 81328 207856
rect 96368 2128 96688 207856
rect 111728 2128 112048 207856
<< obsm4 >>
rect 1715 2483 4128 207637
rect 4608 2483 19488 207637
rect 19968 2483 34848 207637
rect 35328 2483 50208 207637
rect 50688 2483 65568 207637
rect 66048 2483 76485 207637
<< labels >>
rlabel metal2 s 41878 0 41934 800 6 cpu2dmux_ack
port 1 nsew signal output
rlabel metal2 s 92754 209200 92810 210000 6 cpu2dmux_addr[0]
port 2 nsew signal input
rlabel metal3 s 119200 19048 120000 19168 6 cpu2dmux_addr[10]
port 3 nsew signal input
rlabel metal3 s 0 155728 800 155848 6 cpu2dmux_addr[11]
port 4 nsew signal input
rlabel metal3 s 119200 55088 120000 55208 6 cpu2dmux_addr[12]
port 5 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 cpu2dmux_addr[13]
port 6 nsew signal input
rlabel metal3 s 119200 88408 120000 88528 6 cpu2dmux_addr[14]
port 7 nsew signal input
rlabel metal2 s 38658 209200 38714 210000 6 cpu2dmux_addr[15]
port 8 nsew signal input
rlabel metal2 s 74078 209200 74134 210000 6 cpu2dmux_addr[16]
port 9 nsew signal input
rlabel metal2 s 81806 209200 81862 210000 6 cpu2dmux_addr[17]
port 10 nsew signal input
rlabel metal3 s 119200 43528 120000 43648 6 cpu2dmux_addr[18]
port 11 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 cpu2dmux_addr[19]
port 12 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 cpu2dmux_addr[1]
port 13 nsew signal input
rlabel metal3 s 0 145528 800 145648 6 cpu2dmux_addr[20]
port 14 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 cpu2dmux_addr[21]
port 15 nsew signal input
rlabel metal2 s 75366 209200 75422 210000 6 cpu2dmux_addr[22]
port 16 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 cpu2dmux_addr[23]
port 17 nsew signal input
rlabel metal3 s 119200 49648 120000 49768 6 cpu2dmux_addr[24]
port 18 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 cpu2dmux_addr[25]
port 19 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 cpu2dmux_addr[26]
port 20 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 cpu2dmux_addr[27]
port 21 nsew signal input
rlabel metal2 s 117226 209200 117282 210000 6 cpu2dmux_addr[28]
port 22 nsew signal input
rlabel metal2 s 662 209200 718 210000 6 cpu2dmux_addr[29]
port 23 nsew signal input
rlabel metal3 s 119200 133288 120000 133408 6 cpu2dmux_addr[2]
port 24 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 cpu2dmux_addr[30]
port 25 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 cpu2dmux_addr[31]
port 26 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 cpu2dmux_addr[3]
port 27 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 cpu2dmux_addr[4]
port 28 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 cpu2dmux_addr[5]
port 29 nsew signal input
rlabel metal3 s 119200 55768 120000 55888 6 cpu2dmux_addr[6]
port 30 nsew signal input
rlabel metal3 s 119200 161168 120000 161288 6 cpu2dmux_addr[7]
port 31 nsew signal input
rlabel metal2 s 10322 209200 10378 210000 6 cpu2dmux_addr[8]
port 32 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 cpu2dmux_addr[9]
port 33 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 cpu2dmux_bl[0]
port 34 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 cpu2dmux_bl[1]
port 35 nsew signal input
rlabel metal3 s 0 198568 800 198688 6 cpu2dmux_bl[2]
port 36 nsew signal input
rlabel metal3 s 119200 12928 120000 13048 6 cpu2dmux_bl[3]
port 37 nsew signal input
rlabel metal3 s 119200 28568 120000 28688 6 cpu2dmux_bl[4]
port 38 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 cpu2dmux_bl[5]
port 39 nsew signal input
rlabel metal3 s 119200 194488 120000 194608 6 cpu2dmux_bl[6]
port 40 nsew signal input
rlabel metal2 s 16762 209200 16818 210000 6 cpu2dmux_bl[7]
port 41 nsew signal input
rlabel metal3 s 119200 128528 120000 128648 6 cpu2dmux_bl[8]
port 42 nsew signal input
rlabel metal3 s 119200 197208 120000 197328 6 cpu2dmux_bl[9]
port 43 nsew signal input
rlabel metal3 s 119200 19728 120000 19848 6 cpu2dmux_bry
port 44 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 cpu2dmux_cyc
port 45 nsew signal input
rlabel metal3 s 119200 119688 120000 119808 6 cpu2dmux_rdata[0]
port 46 nsew signal output
rlabel metal3 s 119200 1368 120000 1488 6 cpu2dmux_rdata[10]
port 47 nsew signal output
rlabel metal3 s 119200 162528 120000 162648 6 cpu2dmux_rdata[11]
port 48 nsew signal output
rlabel metal2 s 96618 209200 96674 210000 6 cpu2dmux_rdata[12]
port 49 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 cpu2dmux_rdata[13]
port 50 nsew signal output
rlabel metal3 s 119200 182928 120000 183048 6 cpu2dmux_rdata[14]
port 51 nsew signal output
rlabel metal3 s 0 176128 800 176248 6 cpu2dmux_rdata[15]
port 52 nsew signal output
rlabel metal3 s 119200 66648 120000 66768 6 cpu2dmux_rdata[16]
port 53 nsew signal output
rlabel metal3 s 119200 167288 120000 167408 6 cpu2dmux_rdata[17]
port 54 nsew signal output
rlabel metal2 s 78586 209200 78642 210000 6 cpu2dmux_rdata[18]
port 55 nsew signal output
rlabel metal3 s 119200 148248 120000 148368 6 cpu2dmux_rdata[19]
port 56 nsew signal output
rlabel metal2 s 82450 209200 82506 210000 6 cpu2dmux_rdata[1]
port 57 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 cpu2dmux_rdata[20]
port 58 nsew signal output
rlabel metal2 s 47030 209200 47086 210000 6 cpu2dmux_rdata[21]
port 59 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 cpu2dmux_rdata[22]
port 60 nsew signal output
rlabel metal3 s 119200 59168 120000 59288 6 cpu2dmux_rdata[23]
port 61 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 cpu2dmux_rdata[24]
port 62 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 cpu2dmux_rdata[25]
port 63 nsew signal output
rlabel metal3 s 0 172048 800 172168 6 cpu2dmux_rdata[26]
port 64 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 cpu2dmux_rdata[27]
port 65 nsew signal output
rlabel metal2 s 72790 209200 72846 210000 6 cpu2dmux_rdata[28]
port 66 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 cpu2dmux_rdata[29]
port 67 nsew signal output
rlabel metal2 s 23846 209200 23902 210000 6 cpu2dmux_rdata[2]
port 68 nsew signal output
rlabel metal2 s 25778 209200 25834 210000 6 cpu2dmux_rdata[30]
port 69 nsew signal output
rlabel metal2 s 9034 209200 9090 210000 6 cpu2dmux_rdata[31]
port 70 nsew signal output
rlabel metal3 s 119200 38088 120000 38208 6 cpu2dmux_rdata[3]
port 71 nsew signal output
rlabel metal2 s 29642 209200 29698 210000 6 cpu2dmux_rdata[4]
port 72 nsew signal output
rlabel metal2 s 104990 209200 105046 210000 6 cpu2dmux_rdata[5]
port 73 nsew signal output
rlabel metal3 s 119200 206048 120000 206168 6 cpu2dmux_rdata[6]
port 74 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 cpu2dmux_rdata[7]
port 75 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 cpu2dmux_rdata[8]
port 76 nsew signal output
rlabel metal3 s 119200 117648 120000 117768 6 cpu2dmux_rdata[9]
port 77 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 cpu2dmux_sel[0]
port 78 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 cpu2dmux_sel[1]
port 79 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 cpu2dmux_sel[2]
port 80 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 cpu2dmux_sel[3]
port 81 nsew signal input
rlabel metal3 s 0 163208 800 163328 6 cpu2dmux_stb
port 82 nsew signal input
rlabel metal3 s 119200 103368 120000 103488 6 cpu2dmux_wdata[0]
port 83 nsew signal input
rlabel metal3 s 119200 9528 120000 9648 6 cpu2dmux_wdata[10]
port 84 nsew signal input
rlabel metal3 s 119200 183608 120000 183728 6 cpu2dmux_wdata[11]
port 85 nsew signal input
rlabel metal3 s 119200 76848 120000 76968 6 cpu2dmux_wdata[12]
port 86 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 cpu2dmux_wdata[13]
port 87 nsew signal input
rlabel metal3 s 0 188368 800 188488 6 cpu2dmux_wdata[14]
port 88 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 cpu2dmux_wdata[15]
port 89 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 cpu2dmux_wdata[16]
port 90 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 cpu2dmux_wdata[17]
port 91 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 cpu2dmux_wdata[18]
port 92 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 cpu2dmux_wdata[19]
port 93 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 cpu2dmux_wdata[1]
port 94 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 cpu2dmux_wdata[20]
port 95 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 cpu2dmux_wdata[21]
port 96 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 cpu2dmux_wdata[22]
port 97 nsew signal input
rlabel metal2 s 76654 209200 76710 210000 6 cpu2dmux_wdata[23]
port 98 nsew signal input
rlabel metal3 s 119200 25168 120000 25288 6 cpu2dmux_wdata[24]
port 99 nsew signal input
rlabel metal3 s 119200 202648 120000 202768 6 cpu2dmux_wdata[25]
port 100 nsew signal input
rlabel metal2 s 1950 209200 2006 210000 6 cpu2dmux_wdata[26]
port 101 nsew signal input
rlabel metal3 s 119200 142808 120000 142928 6 cpu2dmux_wdata[27]
port 102 nsew signal input
rlabel metal2 s 102414 209200 102470 210000 6 cpu2dmux_wdata[28]
port 103 nsew signal input
rlabel metal3 s 119200 86368 120000 86488 6 cpu2dmux_wdata[29]
port 104 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 cpu2dmux_wdata[2]
port 105 nsew signal input
rlabel metal2 s 86958 209200 87014 210000 6 cpu2dmux_wdata[30]
port 106 nsew signal input
rlabel metal3 s 119200 118328 120000 118448 6 cpu2dmux_wdata[31]
port 107 nsew signal input
rlabel metal3 s 119200 197888 120000 198008 6 cpu2dmux_wdata[3]
port 108 nsew signal input
rlabel metal3 s 119200 149608 120000 149728 6 cpu2dmux_wdata[4]
port 109 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 cpu2dmux_wdata[5]
port 110 nsew signal input
rlabel metal3 s 119200 170688 120000 170808 6 cpu2dmux_wdata[6]
port 111 nsew signal input
rlabel metal2 s 103702 209200 103758 210000 6 cpu2dmux_wdata[7]
port 112 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 cpu2dmux_wdata[8]
port 113 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 cpu2dmux_wdata[9]
port 114 nsew signal input
rlabel metal2 s 40590 209200 40646 210000 6 cpu2dmux_we
port 115 nsew signal input
rlabel metal3 s 119200 123088 120000 123208 6 cpu2imux_ack
port 116 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 cpu2imux_addr[0]
port 117 nsew signal input
rlabel metal3 s 119200 138048 120000 138168 6 cpu2imux_addr[10]
port 118 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 cpu2imux_addr[11]
port 119 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 cpu2imux_addr[12]
port 120 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 cpu2imux_addr[13]
port 121 nsew signal input
rlabel metal3 s 119200 133968 120000 134088 6 cpu2imux_addr[14]
port 122 nsew signal input
rlabel metal3 s 0 165248 800 165368 6 cpu2imux_addr[15]
port 123 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 cpu2imux_addr[16]
port 124 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 cpu2imux_addr[17]
port 125 nsew signal input
rlabel metal3 s 119200 42848 120000 42968 6 cpu2imux_addr[18]
port 126 nsew signal input
rlabel metal3 s 119200 75488 120000 75608 6 cpu2imux_addr[19]
port 127 nsew signal input
rlabel metal2 s 59266 209200 59322 210000 6 cpu2imux_addr[1]
port 128 nsew signal input
rlabel metal3 s 119200 104728 120000 104848 6 cpu2imux_addr[20]
port 129 nsew signal input
rlabel metal3 s 119200 52368 120000 52488 6 cpu2imux_addr[21]
port 130 nsew signal input
rlabel metal3 s 119200 46248 120000 46368 6 cpu2imux_addr[22]
port 131 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 cpu2imux_addr[23]
port 132 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 cpu2imux_addr[24]
port 133 nsew signal input
rlabel metal3 s 119200 145528 120000 145648 6 cpu2imux_addr[25]
port 134 nsew signal input
rlabel metal3 s 0 182248 800 182368 6 cpu2imux_addr[26]
port 135 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 cpu2imux_addr[27]
port 136 nsew signal input
rlabel metal3 s 119200 121048 120000 121168 6 cpu2imux_addr[28]
port 137 nsew signal input
rlabel metal2 s 25134 209200 25190 210000 6 cpu2imux_addr[29]
port 138 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 cpu2imux_addr[2]
port 139 nsew signal input
rlabel metal3 s 119200 62568 120000 62688 6 cpu2imux_addr[30]
port 140 nsew signal input
rlabel metal3 s 119200 176808 120000 176928 6 cpu2imux_addr[31]
port 141 nsew signal input
rlabel metal3 s 119200 208088 120000 208208 6 cpu2imux_addr[3]
port 142 nsew signal input
rlabel metal3 s 119200 73448 120000 73568 6 cpu2imux_addr[4]
port 143 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 cpu2imux_addr[5]
port 144 nsew signal input
rlabel metal2 s 48962 209200 49018 210000 6 cpu2imux_addr[6]
port 145 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 cpu2imux_addr[7]
port 146 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 cpu2imux_addr[8]
port 147 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 cpu2imux_addr[9]
port 148 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 cpu2imux_bl[0]
port 149 nsew signal input
rlabel metal2 s 662 0 718 800 6 cpu2imux_bl[1]
port 150 nsew signal input
rlabel metal3 s 119200 26528 120000 26648 6 cpu2imux_bl[2]
port 151 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 cpu2imux_bl[3]
port 152 nsew signal input
rlabel metal2 s 31574 209200 31630 210000 6 cpu2imux_bl[4]
port 153 nsew signal input
rlabel metal2 s 27066 209200 27122 210000 6 cpu2imux_bl[5]
port 154 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 cpu2imux_bl[6]
port 155 nsew signal input
rlabel metal3 s 119200 129888 120000 130008 6 cpu2imux_bl[7]
port 156 nsew signal input
rlabel metal2 s 63130 209200 63186 210000 6 cpu2imux_bl[8]
port 157 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 cpu2imux_bl[9]
port 158 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 cpu2imux_bry
port 159 nsew signal input
rlabel metal3 s 0 185648 800 185768 6 cpu2imux_cyc
port 160 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 cpu2imux_rdata[0]
port 161 nsew signal output
rlabel metal3 s 119200 76168 120000 76288 6 cpu2imux_rdata[10]
port 162 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 cpu2imux_rdata[11]
port 163 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 cpu2imux_rdata[12]
port 164 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 cpu2imux_rdata[13]
port 165 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 cpu2imux_rdata[14]
port 166 nsew signal output
rlabel metal3 s 119200 193128 120000 193248 6 cpu2imux_rdata[15]
port 167 nsew signal output
rlabel metal3 s 119200 169328 120000 169448 6 cpu2imux_rdata[16]
port 168 nsew signal output
rlabel metal2 s 68282 209200 68338 210000 6 cpu2imux_rdata[17]
port 169 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 cpu2imux_rdata[18]
port 170 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 cpu2imux_rdata[19]
port 171 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 cpu2imux_rdata[1]
port 172 nsew signal output
rlabel metal3 s 119200 106768 120000 106888 6 cpu2imux_rdata[20]
port 173 nsew signal output
rlabel metal3 s 119200 156408 120000 156528 6 cpu2imux_rdata[21]
port 174 nsew signal output
rlabel metal3 s 119200 188368 120000 188488 6 cpu2imux_rdata[22]
port 175 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 cpu2imux_rdata[23]
port 176 nsew signal output
rlabel metal3 s 119200 95208 120000 95328 6 cpu2imux_rdata[24]
port 177 nsew signal output
rlabel metal3 s 119200 114928 120000 115048 6 cpu2imux_rdata[25]
port 178 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 cpu2imux_rdata[26]
port 179 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 cpu2imux_rdata[27]
port 180 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 cpu2imux_rdata[28]
port 181 nsew signal output
rlabel metal3 s 119200 85688 120000 85808 6 cpu2imux_rdata[29]
port 182 nsew signal output
rlabel metal3 s 119200 69368 120000 69488 6 cpu2imux_rdata[2]
port 183 nsew signal output
rlabel metal3 s 119200 208768 120000 208888 6 cpu2imux_rdata[30]
port 184 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 cpu2imux_rdata[31]
port 185 nsew signal output
rlabel metal3 s 119200 175448 120000 175568 6 cpu2imux_rdata[3]
port 186 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 cpu2imux_rdata[4]
port 187 nsew signal output
rlabel metal2 s 110142 209200 110198 210000 6 cpu2imux_rdata[5]
port 188 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 cpu2imux_rdata[6]
port 189 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 cpu2imux_rdata[7]
port 190 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 cpu2imux_rdata[8]
port 191 nsew signal output
rlabel metal2 s 53470 209200 53526 210000 6 cpu2imux_rdata[9]
port 192 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 cpu2imux_stb
port 193 nsew signal input
rlabel metal3 s 119200 40808 120000 40928 6 cpu2imux_we
port 194 nsew signal input
rlabel metal2 s 71502 209200 71558 210000 6 dram_addr0[0]
port 195 nsew signal output
rlabel metal3 s 119200 100648 120000 100768 6 dram_addr0[1]
port 196 nsew signal output
rlabel metal3 s 119200 204688 120000 204808 6 dram_addr0[2]
port 197 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 dram_addr0[3]
port 198 nsew signal output
rlabel metal3 s 119200 2728 120000 2848 6 dram_addr0[4]
port 199 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 dram_addr0[5]
port 200 nsew signal output
rlabel metal3 s 119200 199928 120000 200048 6 dram_addr0[6]
port 201 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 dram_addr0[7]
port 202 nsew signal output
rlabel metal3 s 119200 22448 120000 22568 6 dram_clk0
port 203 nsew signal output
rlabel metal3 s 0 202648 800 202768 6 dram_csb0
port 204 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 dram_din0[0]
port 205 nsew signal output
rlabel metal2 s 15474 209200 15530 210000 6 dram_din0[10]
port 206 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 dram_din0[11]
port 207 nsew signal output
rlabel metal3 s 119200 200608 120000 200728 6 dram_din0[12]
port 208 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 dram_din0[13]
port 209 nsew signal output
rlabel metal3 s 119200 191768 120000 191888 6 dram_din0[14]
port 210 nsew signal output
rlabel metal3 s 0 161848 800 161968 6 dram_din0[15]
port 211 nsew signal output
rlabel metal3 s 119200 115608 120000 115728 6 dram_din0[16]
port 212 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 dram_din0[17]
port 213 nsew signal output
rlabel metal2 s 41234 209200 41290 210000 6 dram_din0[18]
port 214 nsew signal output
rlabel metal2 s 12254 209200 12310 210000 6 dram_din0[19]
port 215 nsew signal output
rlabel metal2 s 70858 209200 70914 210000 6 dram_din0[1]
port 216 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 dram_din0[20]
port 217 nsew signal output
rlabel metal3 s 0 180888 800 181008 6 dram_din0[21]
port 218 nsew signal output
rlabel metal3 s 119200 89768 120000 89888 6 dram_din0[22]
port 219 nsew signal output
rlabel metal3 s 119200 155048 120000 155168 6 dram_din0[23]
port 220 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 dram_din0[24]
port 221 nsew signal output
rlabel metal3 s 0 204688 800 204808 6 dram_din0[25]
port 222 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 dram_din0[26]
port 223 nsew signal output
rlabel metal3 s 0 195168 800 195288 6 dram_din0[27]
port 224 nsew signal output
rlabel metal3 s 119200 68008 120000 68128 6 dram_din0[28]
port 225 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 dram_din0[29]
port 226 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 dram_din0[2]
port 227 nsew signal output
rlabel metal3 s 0 146208 800 146328 6 dram_din0[30]
port 228 nsew signal output
rlabel metal3 s 119200 120368 120000 120488 6 dram_din0[31]
port 229 nsew signal output
rlabel metal3 s 119200 18368 120000 18488 6 dram_din0[3]
port 230 nsew signal output
rlabel metal3 s 119200 151648 120000 151768 6 dram_din0[4]
port 231 nsew signal output
rlabel metal2 s 36082 209200 36138 210000 6 dram_din0[5]
port 232 nsew signal output
rlabel metal3 s 119200 6128 120000 6248 6 dram_din0[6]
port 233 nsew signal output
rlabel metal2 s 68926 209200 68982 210000 6 dram_din0[7]
port 234 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 dram_din0[8]
port 235 nsew signal output
rlabel metal3 s 119200 27888 120000 28008 6 dram_din0[9]
port 236 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 dram_dout0[0]
port 237 nsew signal input
rlabel metal3 s 0 193128 800 193248 6 dram_dout0[10]
port 238 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 dram_dout0[11]
port 239 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 dram_dout0[12]
port 240 nsew signal input
rlabel metal2 s 42522 209200 42578 210000 6 dram_dout0[13]
port 241 nsew signal input
rlabel metal2 s 77942 209200 77998 210000 6 dram_dout0[14]
port 242 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 dram_dout0[15]
port 243 nsew signal input
rlabel metal2 s 88246 209200 88302 210000 6 dram_dout0[16]
port 244 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 dram_dout0[17]
port 245 nsew signal input
rlabel metal3 s 119200 195848 120000 195968 6 dram_dout0[18]
port 246 nsew signal input
rlabel metal3 s 119200 10208 120000 10328 6 dram_dout0[19]
port 247 nsew signal input
rlabel metal3 s 119200 35368 120000 35488 6 dram_dout0[1]
port 248 nsew signal input
rlabel metal3 s 119200 165248 120000 165368 6 dram_dout0[20]
port 249 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 dram_dout0[21]
port 250 nsew signal input
rlabel metal3 s 119200 71408 120000 71528 6 dram_dout0[22]
port 251 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 dram_dout0[23]
port 252 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 dram_dout0[24]
port 253 nsew signal input
rlabel metal3 s 0 174088 800 174208 6 dram_dout0[25]
port 254 nsew signal input
rlabel metal3 s 119200 61208 120000 61328 6 dram_dout0[26]
port 255 nsew signal input
rlabel metal3 s 119200 126488 120000 126608 6 dram_dout0[27]
port 256 nsew signal input
rlabel metal3 s 119200 203328 120000 203448 6 dram_dout0[28]
port 257 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 dram_dout0[29]
port 258 nsew signal input
rlabel metal3 s 0 161168 800 161288 6 dram_dout0[2]
port 259 nsew signal input
rlabel metal3 s 0 197888 800 198008 6 dram_dout0[30]
port 260 nsew signal input
rlabel metal3 s 119200 176128 120000 176248 6 dram_dout0[31]
port 261 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 dram_dout0[3]
port 262 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 dram_dout0[4]
port 263 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 dram_dout0[5]
port 264 nsew signal input
rlabel metal2 s 38014 209200 38070 210000 6 dram_dout0[6]
port 265 nsew signal input
rlabel metal2 s 79230 209200 79286 210000 6 dram_dout0[7]
port 266 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 dram_dout0[8]
port 267 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 dram_dout0[9]
port 268 nsew signal input
rlabel metal2 s 66350 209200 66406 210000 6 dram_web0
port 269 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 dram_wmask0[0]
port 270 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 dram_wmask0[1]
port 271 nsew signal output
rlabel metal3 s 119200 172048 120000 172168 6 dram_wmask0[2]
port 272 nsew signal output
rlabel metal3 s 119200 160488 120000 160608 6 dram_wmask0[3]
port 273 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 gpio_in[0]
port 274 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 gpio_in[10]
port 275 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 gpio_in[11]
port 276 nsew signal input
rlabel metal3 s 0 204008 800 204128 6 gpio_in[12]
port 277 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 gpio_in[13]
port 278 nsew signal input
rlabel metal3 s 119200 165928 120000 166048 6 gpio_in[14]
port 279 nsew signal input
rlabel metal2 s 110786 209200 110842 210000 6 gpio_in[15]
port 280 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 gpio_in[16]
port 281 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 gpio_in[17]
port 282 nsew signal input
rlabel metal2 s 36726 209200 36782 210000 6 gpio_in[18]
port 283 nsew signal input
rlabel metal2 s 30930 209200 30986 210000 6 gpio_in[19]
port 284 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 gpio_in[1]
port 285 nsew signal input
rlabel metal3 s 0 187688 800 187808 6 gpio_in[20]
port 286 nsew signal input
rlabel metal3 s 119200 81608 120000 81728 6 gpio_in[21]
port 287 nsew signal input
rlabel metal3 s 119200 136008 120000 136128 6 gpio_in[22]
port 288 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 gpio_in[23]
port 289 nsew signal input
rlabel metal3 s 119200 14968 120000 15088 6 gpio_in[2]
port 290 nsew signal input
rlabel metal3 s 119200 72088 120000 72208 6 gpio_in[3]
port 291 nsew signal input
rlabel metal3 s 119200 46928 120000 47048 6 gpio_in[4]
port 292 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 gpio_in[5]
port 293 nsew signal input
rlabel metal3 s 119200 140768 120000 140888 6 gpio_in[6]
port 294 nsew signal input
rlabel metal2 s 94042 209200 94098 210000 6 gpio_in[7]
port 295 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 gpio_in[8]
port 296 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 gpio_in[9]
port 297 nsew signal input
rlabel metal3 s 119200 163888 120000 164008 6 gpio_oeb[0]
port 298 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 gpio_oeb[10]
port 299 nsew signal output
rlabel metal3 s 0 179528 800 179648 6 gpio_oeb[11]
port 300 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 gpio_oeb[12]
port 301 nsew signal output
rlabel metal3 s 119200 153688 120000 153808 6 gpio_oeb[13]
port 302 nsew signal output
rlabel metal2 s 95330 209200 95386 210000 6 gpio_oeb[14]
port 303 nsew signal output
rlabel metal2 s 34150 209200 34206 210000 6 gpio_oeb[15]
port 304 nsew signal output
rlabel metal2 s 50250 209200 50306 210000 6 gpio_oeb[16]
port 305 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 gpio_oeb[17]
port 306 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 gpio_oeb[18]
port 307 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 gpio_oeb[19]
port 308 nsew signal output
rlabel metal3 s 119200 29928 120000 30048 6 gpio_oeb[1]
port 309 nsew signal output
rlabel metal3 s 119200 4768 120000 4888 6 gpio_oeb[20]
port 310 nsew signal output
rlabel metal3 s 119200 141448 120000 141568 6 gpio_oeb[21]
port 311 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 gpio_oeb[22]
port 312 nsew signal output
rlabel metal2 s 73434 209200 73490 210000 6 gpio_oeb[23]
port 313 nsew signal output
rlabel metal3 s 119200 34008 120000 34128 6 gpio_oeb[24]
port 314 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 gpio_oeb[25]
port 315 nsew signal output
rlabel metal3 s 119200 159808 120000 159928 6 gpio_oeb[26]
port 316 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 gpio_oeb[27]
port 317 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 gpio_oeb[28]
port 318 nsew signal output
rlabel metal2 s 79874 209200 79930 210000 6 gpio_oeb[29]
port 319 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 gpio_oeb[2]
port 320 nsew signal output
rlabel metal3 s 119200 173408 120000 173528 6 gpio_oeb[30]
port 321 nsew signal output
rlabel metal3 s 119200 150968 120000 151088 6 gpio_oeb[31]
port 322 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 gpio_oeb[32]
port 323 nsew signal output
rlabel metal3 s 0 178168 800 178288 6 gpio_oeb[33]
port 324 nsew signal output
rlabel metal2 s 61842 209200 61898 210000 6 gpio_oeb[34]
port 325 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 gpio_oeb[35]
port 326 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 gpio_oeb[36]
port 327 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 gpio_oeb[37]
port 328 nsew signal output
rlabel metal3 s 119200 174088 120000 174208 6 gpio_oeb[3]
port 329 nsew signal output
rlabel metal2 s 18694 209200 18750 210000 6 gpio_oeb[4]
port 330 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 gpio_oeb[5]
port 331 nsew signal output
rlabel metal2 s 60554 209200 60610 210000 6 gpio_oeb[6]
port 332 nsew signal output
rlabel metal3 s 119200 174768 120000 174888 6 gpio_oeb[7]
port 333 nsew signal output
rlabel metal3 s 119200 34688 120000 34808 6 gpio_oeb[8]
port 334 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 gpio_oeb[9]
port 335 nsew signal output
rlabel metal2 s 114650 209200 114706 210000 6 gpio_out[0]
port 336 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 gpio_out[10]
port 337 nsew signal output
rlabel metal3 s 119200 99968 120000 100088 6 gpio_out[11]
port 338 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 gpio_out[12]
port 339 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 gpio_out[13]
port 340 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 gpio_out[14]
port 341 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 gpio_out[15]
port 342 nsew signal output
rlabel metal3 s 119200 184968 120000 185088 6 gpio_out[16]
port 343 nsew signal output
rlabel metal3 s 0 189728 800 189848 6 gpio_out[17]
port 344 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 gpio_out[18]
port 345 nsew signal output
rlabel metal3 s 0 126488 800 126608 6 gpio_out[19]
port 346 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 gpio_out[1]
port 347 nsew signal output
rlabel metal3 s 119200 65968 120000 66088 6 gpio_out[20]
port 348 nsew signal output
rlabel metal3 s 0 121728 800 121848 6 gpio_out[21]
port 349 nsew signal output
rlabel metal2 s 112074 209200 112130 210000 6 gpio_out[22]
port 350 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 gpio_out[23]
port 351 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 gpio_out[2]
port 352 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 gpio_out[3]
port 353 nsew signal output
rlabel metal3 s 119200 114248 120000 114368 6 gpio_out[4]
port 354 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 gpio_out[5]
port 355 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 gpio_out[6]
port 356 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 gpio_out[7]
port 357 nsew signal output
rlabel metal3 s 0 191088 800 191208 6 gpio_out[8]
port 358 nsew signal output
rlabel metal3 s 119200 48288 120000 48408 6 gpio_out[9]
port 359 nsew signal output
rlabel metal3 s 119200 8168 120000 8288 6 iram_addr0[0]
port 360 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 iram_addr0[1]
port 361 nsew signal output
rlabel metal3 s 0 201968 800 202088 6 iram_addr0[2]
port 362 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 iram_addr0[3]
port 363 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 iram_addr0[4]
port 364 nsew signal output
rlabel metal3 s 119200 87048 120000 87168 6 iram_addr0[5]
port 365 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 iram_addr0[6]
port 366 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 iram_addr0[7]
port 367 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 iram_clk0
port 368 nsew signal output
rlabel metal3 s 119200 205368 120000 205488 6 iram_csb0_A
port 369 nsew signal output
rlabel metal3 s 119200 159128 120000 159248 6 iram_csb0_B
port 370 nsew signal output
rlabel metal3 s 0 201288 800 201408 6 iram_din0[0]
port 371 nsew signal output
rlabel metal3 s 119200 157088 120000 157208 6 iram_din0[10]
port 372 nsew signal output
rlabel metal3 s 0 148928 800 149048 6 iram_din0[11]
port 373 nsew signal output
rlabel metal2 s 58622 209200 58678 210000 6 iram_din0[12]
port 374 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 iram_din0[13]
port 375 nsew signal output
rlabel metal2 s 67638 209200 67694 210000 6 iram_din0[14]
port 376 nsew signal output
rlabel metal3 s 119200 201968 120000 202088 6 iram_din0[15]
port 377 nsew signal output
rlabel metal3 s 0 174768 800 174888 6 iram_din0[16]
port 378 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 iram_din0[17]
port 379 nsew signal output
rlabel metal3 s 119200 91128 120000 91248 6 iram_din0[18]
port 380 nsew signal output
rlabel metal3 s 119200 144168 120000 144288 6 iram_din0[19]
port 381 nsew signal output
rlabel metal3 s 119200 147568 120000 147688 6 iram_din0[1]
port 382 nsew signal output
rlabel metal2 s 20626 209200 20682 210000 6 iram_din0[20]
port 383 nsew signal output
rlabel metal2 s 63774 209200 63830 210000 6 iram_din0[21]
port 384 nsew signal output
rlabel metal3 s 119200 104048 120000 104168 6 iram_din0[22]
port 385 nsew signal output
rlabel metal2 s 19982 209200 20038 210000 6 iram_din0[23]
port 386 nsew signal output
rlabel metal2 s 48318 209200 48374 210000 6 iram_din0[24]
port 387 nsew signal output
rlabel metal2 s 8390 209200 8446 210000 6 iram_din0[25]
port 388 nsew signal output
rlabel metal3 s 119200 186328 120000 186448 6 iram_din0[26]
port 389 nsew signal output
rlabel metal3 s 119200 20408 120000 20528 6 iram_din0[27]
port 390 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 iram_din0[28]
port 391 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 iram_din0[29]
port 392 nsew signal output
rlabel metal2 s 99194 209200 99250 210000 6 iram_din0[2]
port 393 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 iram_din0[30]
port 394 nsew signal output
rlabel metal3 s 119200 57808 120000 57928 6 iram_din0[31]
port 395 nsew signal output
rlabel metal3 s 0 171368 800 171488 6 iram_din0[3]
port 396 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 iram_din0[4]
port 397 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 iram_din0[5]
port 398 nsew signal output
rlabel metal3 s 119200 33328 120000 33448 6 iram_din0[6]
port 399 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 iram_din0[7]
port 400 nsew signal output
rlabel metal2 s 115294 209200 115350 210000 6 iram_din0[8]
port 401 nsew signal output
rlabel metal2 s 45742 209200 45798 210000 6 iram_din0[9]
port 402 nsew signal output
rlabel metal3 s 119200 122408 120000 122528 6 iram_dout0_A[0]
port 403 nsew signal input
rlabel metal3 s 0 190408 800 190528 6 iram_dout0_A[10]
port 404 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 iram_dout0_A[11]
port 405 nsew signal input
rlabel metal2 s 101770 209200 101826 210000 6 iram_dout0_A[12]
port 406 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 iram_dout0_A[13]
port 407 nsew signal input
rlabel metal3 s 119200 72768 120000 72888 6 iram_dout0_A[14]
port 408 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 iram_dout0_A[15]
port 409 nsew signal input
rlabel metal3 s 119200 58488 120000 58608 6 iram_dout0_A[16]
port 410 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 iram_dout0_A[17]
port 411 nsew signal input
rlabel metal3 s 0 155048 800 155168 6 iram_dout0_A[18]
port 412 nsew signal input
rlabel metal3 s 119200 53728 120000 53848 6 iram_dout0_A[19]
port 413 nsew signal input
rlabel metal3 s 119200 17688 120000 17808 6 iram_dout0_A[1]
port 414 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 iram_dout0_A[20]
port 415 nsew signal input
rlabel metal3 s 119200 21088 120000 21208 6 iram_dout0_A[21]
port 416 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 iram_dout0_A[22]
port 417 nsew signal input
rlabel metal2 s 85026 209200 85082 210000 6 iram_dout0_A[23]
port 418 nsew signal input
rlabel metal3 s 0 170688 800 170808 6 iram_dout0_A[24]
port 419 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 iram_dout0_A[25]
port 420 nsew signal input
rlabel metal2 s 33506 209200 33562 210000 6 iram_dout0_A[26]
port 421 nsew signal input
rlabel metal2 s 17406 209200 17462 210000 6 iram_dout0_A[27]
port 422 nsew signal input
rlabel metal3 s 0 157768 800 157888 6 iram_dout0_A[28]
port 423 nsew signal input
rlabel metal2 s 90178 209200 90234 210000 6 iram_dout0_A[29]
port 424 nsew signal input
rlabel metal2 s 86314 209200 86370 210000 6 iram_dout0_A[2]
port 425 nsew signal input
rlabel metal2 s 99838 209200 99894 210000 6 iram_dout0_A[30]
port 426 nsew signal input
rlabel metal2 s 13542 209200 13598 210000 6 iram_dout0_A[31]
port 427 nsew signal input
rlabel metal2 s 50894 209200 50950 210000 6 iram_dout0_A[3]
port 428 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 iram_dout0_A[4]
port 429 nsew signal input
rlabel metal2 s 100482 209200 100538 210000 6 iram_dout0_A[5]
port 430 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 iram_dout0_A[6]
port 431 nsew signal input
rlabel metal3 s 119200 82968 120000 83088 6 iram_dout0_A[7]
port 432 nsew signal input
rlabel metal3 s 119200 129208 120000 129328 6 iram_dout0_A[8]
port 433 nsew signal input
rlabel metal3 s 119200 97248 120000 97368 6 iram_dout0_A[9]
port 434 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 iram_dout0_B[0]
port 435 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 iram_dout0_B[10]
port 436 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 iram_dout0_B[11]
port 437 nsew signal input
rlabel metal3 s 119200 31288 120000 31408 6 iram_dout0_B[12]
port 438 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 iram_dout0_B[13]
port 439 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 iram_dout0_B[14]
port 440 nsew signal input
rlabel metal2 s 7102 209200 7158 210000 6 iram_dout0_B[15]
port 441 nsew signal input
rlabel metal2 s 23202 209200 23258 210000 6 iram_dout0_B[16]
port 442 nsew signal input
rlabel metal3 s 119200 80248 120000 80368 6 iram_dout0_B[17]
port 443 nsew signal input
rlabel metal3 s 119200 63248 120000 63368 6 iram_dout0_B[18]
port 444 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 iram_dout0_B[19]
port 445 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 iram_dout0_B[1]
port 446 nsew signal input
rlabel metal3 s 0 133968 800 134088 6 iram_dout0_B[20]
port 447 nsew signal input
rlabel metal3 s 119200 51008 120000 51128 6 iram_dout0_B[21]
port 448 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 iram_dout0_B[22]
port 449 nsew signal input
rlabel metal3 s 119200 91808 120000 91928 6 iram_dout0_B[23]
port 450 nsew signal input
rlabel metal3 s 119200 138728 120000 138848 6 iram_dout0_B[24]
port 451 nsew signal input
rlabel metal3 s 119200 206728 120000 206848 6 iram_dout0_B[25]
port 452 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 iram_dout0_B[26]
port 453 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 iram_dout0_B[27]
port 454 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 iram_dout0_B[28]
port 455 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 iram_dout0_B[29]
port 456 nsew signal input
rlabel metal3 s 119200 27208 120000 27328 6 iram_dout0_B[2]
port 457 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 iram_dout0_B[30]
port 458 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 iram_dout0_B[31]
port 459 nsew signal input
rlabel metal3 s 0 166608 800 166728 6 iram_dout0_B[3]
port 460 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 iram_dout0_B[4]
port 461 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 iram_dout0_B[5]
port 462 nsew signal input
rlabel metal2 s 52182 209200 52238 210000 6 iram_dout0_B[6]
port 463 nsew signal input
rlabel metal2 s 98550 209200 98606 210000 6 iram_dout0_B[7]
port 464 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 iram_dout0_B[8]
port 465 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 iram_dout0_B[9]
port 466 nsew signal input
rlabel metal3 s 119200 192448 120000 192568 6 iram_web0
port 467 nsew signal output
rlabel metal3 s 119200 187688 120000 187808 6 iram_wmask0[0]
port 468 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 iram_wmask0[1]
port 469 nsew signal output
rlabel metal3 s 119200 190408 120000 190528 6 iram_wmask0[2]
port 470 nsew signal output
rlabel metal3 s 119200 54408 120000 54528 6 iram_wmask0[3]
port 471 nsew signal output
rlabel metal2 s 21270 209200 21326 210000 6 la_data_in[0]
port 472 nsew signal input
rlabel metal3 s 0 205368 800 205488 6 la_data_in[100]
port 473 nsew signal input
rlabel metal3 s 119200 180208 120000 180328 6 la_data_in[101]
port 474 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 la_data_in[102]
port 475 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 la_data_in[103]
port 476 nsew signal input
rlabel metal2 s 112718 209200 112774 210000 6 la_data_in[104]
port 477 nsew signal input
rlabel metal2 s 106922 209200 106978 210000 6 la_data_in[105]
port 478 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 la_data_in[106]
port 479 nsew signal input
rlabel metal2 s 69570 209200 69626 210000 6 la_data_in[107]
port 480 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[108]
port 481 nsew signal input
rlabel metal2 s 19338 209200 19394 210000 6 la_data_in[109]
port 482 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 la_data_in[10]
port 483 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 la_data_in[110]
port 484 nsew signal input
rlabel metal3 s 119200 209448 120000 209568 6 la_data_in[111]
port 485 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 la_data_in[112]
port 486 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 la_data_in[113]
port 487 nsew signal input
rlabel metal3 s 119200 92488 120000 92608 6 la_data_in[114]
port 488 nsew signal input
rlabel metal2 s 81162 209200 81218 210000 6 la_data_in[115]
port 489 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 la_data_in[116]
port 490 nsew signal input
rlabel metal3 s 119200 68688 120000 68808 6 la_data_in[117]
port 491 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[118]
port 492 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 la_data_in[119]
port 493 nsew signal input
rlabel metal3 s 119200 121728 120000 121848 6 la_data_in[11]
port 494 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_data_in[120]
port 495 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[121]
port 496 nsew signal input
rlabel metal3 s 119200 172728 120000 172848 6 la_data_in[122]
port 497 nsew signal input
rlabel metal3 s 119200 44208 120000 44328 6 la_data_in[123]
port 498 nsew signal input
rlabel metal3 s 119200 105408 120000 105528 6 la_data_in[124]
port 499 nsew signal input
rlabel metal3 s 119200 74128 120000 74248 6 la_data_in[125]
port 500 nsew signal input
rlabel metal3 s 119200 98608 120000 98728 6 la_data_in[126]
port 501 nsew signal input
rlabel metal3 s 119200 48968 120000 49088 6 la_data_in[127]
port 502 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 la_data_in[12]
port 503 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_data_in[13]
port 504 nsew signal input
rlabel metal3 s 119200 25848 120000 25968 6 la_data_in[14]
port 505 nsew signal input
rlabel metal3 s 119200 95888 120000 96008 6 la_data_in[15]
port 506 nsew signal input
rlabel metal3 s 119200 193808 120000 193928 6 la_data_in[16]
port 507 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 la_data_in[17]
port 508 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 la_data_in[18]
port 509 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_data_in[19]
port 510 nsew signal input
rlabel metal2 s 108210 209200 108266 210000 6 la_data_in[1]
port 511 nsew signal input
rlabel metal2 s 109498 209200 109554 210000 6 la_data_in[20]
port 512 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 la_data_in[21]
port 513 nsew signal input
rlabel metal2 s 41878 209200 41934 210000 6 la_data_in[22]
port 514 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 la_data_in[23]
port 515 nsew signal input
rlabel metal3 s 0 163888 800 164008 6 la_data_in[24]
port 516 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 la_data_in[25]
port 517 nsew signal input
rlabel metal3 s 119200 5448 120000 5568 6 la_data_in[26]
port 518 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 la_data_in[27]
port 519 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[28]
port 520 nsew signal input
rlabel metal3 s 119200 70048 120000 70168 6 la_data_in[29]
port 521 nsew signal input
rlabel metal3 s 119200 79568 120000 79688 6 la_data_in[2]
port 522 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[30]
port 523 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 la_data_in[31]
port 524 nsew signal input
rlabel metal3 s 119200 136688 120000 136808 6 la_data_in[32]
port 525 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 la_data_in[33]
port 526 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 la_data_in[34]
port 527 nsew signal input
rlabel metal3 s 119200 112208 120000 112328 6 la_data_in[35]
port 528 nsew signal input
rlabel metal3 s 119200 7488 120000 7608 6 la_data_in[36]
port 529 nsew signal input
rlabel metal3 s 119200 148928 120000 149048 6 la_data_in[37]
port 530 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 la_data_in[38]
port 531 nsew signal input
rlabel metal3 s 0 195848 800 195968 6 la_data_in[39]
port 532 nsew signal input
rlabel metal2 s 80518 209200 80574 210000 6 la_data_in[3]
port 533 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[40]
port 534 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 la_data_in[41]
port 535 nsew signal input
rlabel metal3 s 119200 139408 120000 139528 6 la_data_in[42]
port 536 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[43]
port 537 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[44]
port 538 nsew signal input
rlabel metal2 s 84382 209200 84438 210000 6 la_data_in[45]
port 539 nsew signal input
rlabel metal3 s 119200 119008 120000 119128 6 la_data_in[46]
port 540 nsew signal input
rlabel metal2 s 35438 209200 35494 210000 6 la_data_in[47]
port 541 nsew signal input
rlabel metal3 s 119200 134648 120000 134768 6 la_data_in[48]
port 542 nsew signal input
rlabel metal3 s 119200 56448 120000 56568 6 la_data_in[49]
port 543 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 la_data_in[4]
port 544 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 la_data_in[50]
port 545 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[51]
port 546 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 la_data_in[52]
port 547 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 la_data_in[53]
port 548 nsew signal input
rlabel metal2 s 85670 209200 85726 210000 6 la_data_in[54]
port 549 nsew signal input
rlabel metal3 s 119200 127168 120000 127288 6 la_data_in[55]
port 550 nsew signal input
rlabel metal2 s 12898 209200 12954 210000 6 la_data_in[56]
port 551 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[57]
port 552 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 la_data_in[58]
port 553 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[59]
port 554 nsew signal input
rlabel metal2 s 3882 209200 3938 210000 6 la_data_in[5]
port 555 nsew signal input
rlabel metal3 s 119200 108128 120000 108248 6 la_data_in[60]
port 556 nsew signal input
rlabel metal3 s 119200 132608 120000 132728 6 la_data_in[61]
port 557 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 la_data_in[62]
port 558 nsew signal input
rlabel metal3 s 119200 179528 120000 179648 6 la_data_in[63]
port 559 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[64]
port 560 nsew signal input
rlabel metal2 s 43810 209200 43866 210000 6 la_data_in[65]
port 561 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[66]
port 562 nsew signal input
rlabel metal3 s 119200 207408 120000 207528 6 la_data_in[67]
port 563 nsew signal input
rlabel metal2 s 6458 209200 6514 210000 6 la_data_in[68]
port 564 nsew signal input
rlabel metal2 s 30286 209200 30342 210000 6 la_data_in[69]
port 565 nsew signal input
rlabel metal2 s 28354 209200 28410 210000 6 la_data_in[6]
port 566 nsew signal input
rlabel metal3 s 0 209448 800 209568 6 la_data_in[70]
port 567 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 la_data_in[71]
port 568 nsew signal input
rlabel metal2 s 116582 209200 116638 210000 6 la_data_in[72]
port 569 nsew signal input
rlabel metal2 s 56690 209200 56746 210000 6 la_data_in[73]
port 570 nsew signal input
rlabel metal2 s 47674 209200 47730 210000 6 la_data_in[74]
port 571 nsew signal input
rlabel metal3 s 0 158448 800 158568 6 la_data_in[75]
port 572 nsew signal input
rlabel metal3 s 119200 153008 120000 153128 6 la_data_in[76]
port 573 nsew signal input
rlabel metal3 s 119200 12248 120000 12368 6 la_data_in[77]
port 574 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 la_data_in[78]
port 575 nsew signal input
rlabel metal3 s 0 173408 800 173528 6 la_data_in[79]
port 576 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[7]
port 577 nsew signal input
rlabel metal3 s 119200 127848 120000 127968 6 la_data_in[80]
port 578 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 la_data_in[81]
port 579 nsew signal input
rlabel metal2 s 54758 209200 54814 210000 6 la_data_in[82]
port 580 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 la_data_in[83]
port 581 nsew signal input
rlabel metal2 s 93398 209200 93454 210000 6 la_data_in[84]
port 582 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 la_data_in[85]
port 583 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[86]
port 584 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 la_data_in[87]
port 585 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[88]
port 586 nsew signal input
rlabel metal2 s 45098 209200 45154 210000 6 la_data_in[89]
port 587 nsew signal input
rlabel metal3 s 119200 90448 120000 90568 6 la_data_in[8]
port 588 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 la_data_in[90]
port 589 nsew signal input
rlabel metal3 s 119200 101328 120000 101448 6 la_data_in[91]
port 590 nsew signal input
rlabel metal2 s 55402 209200 55458 210000 6 la_data_in[92]
port 591 nsew signal input
rlabel metal3 s 0 199928 800 200048 6 la_data_in[93]
port 592 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[94]
port 593 nsew signal input
rlabel metal3 s 119200 146888 120000 147008 6 la_data_in[95]
port 594 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 la_data_in[96]
port 595 nsew signal input
rlabel metal2 s 10966 209200 11022 210000 6 la_data_in[97]
port 596 nsew signal input
rlabel metal3 s 119200 163208 120000 163328 6 la_data_in[98]
port 597 nsew signal input
rlabel metal2 s 92110 209200 92166 210000 6 la_data_in[99]
port 598 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 la_data_in[9]
port 599 nsew signal input
rlabel metal2 s 72146 209200 72202 210000 6 la_data_out[0]
port 600 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[100]
port 601 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[101]
port 602 nsew signal output
rlabel metal3 s 119200 182248 120000 182368 6 la_data_out[102]
port 603 nsew signal output
rlabel metal3 s 119200 16328 120000 16448 6 la_data_out[103]
port 604 nsew signal output
rlabel metal3 s 119200 157768 120000 157888 6 la_data_out[104]
port 605 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 la_data_out[105]
port 606 nsew signal output
rlabel metal2 s 103058 209200 103114 210000 6 la_data_out[106]
port 607 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 la_data_out[107]
port 608 nsew signal output
rlabel metal3 s 119200 93168 120000 93288 6 la_data_out[108]
port 609 nsew signal output
rlabel metal3 s 0 186328 800 186448 6 la_data_out[109]
port 610 nsew signal output
rlabel metal3 s 119200 42168 120000 42288 6 la_data_out[10]
port 611 nsew signal output
rlabel metal2 s 26422 209200 26478 210000 6 la_data_out[110]
port 612 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 la_data_out[111]
port 613 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 la_data_out[112]
port 614 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 la_data_out[113]
port 615 nsew signal output
rlabel metal3 s 119200 150288 120000 150408 6 la_data_out[114]
port 616 nsew signal output
rlabel metal3 s 0 154368 800 154488 6 la_data_out[115]
port 617 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[116]
port 618 nsew signal output
rlabel metal2 s 107566 209200 107622 210000 6 la_data_out[117]
port 619 nsew signal output
rlabel metal3 s 119200 94528 120000 94648 6 la_data_out[118]
port 620 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 la_data_out[119]
port 621 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 la_data_out[11]
port 622 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 la_data_out[120]
port 623 nsew signal output
rlabel metal3 s 119200 167968 120000 168088 6 la_data_out[121]
port 624 nsew signal output
rlabel metal3 s 0 200608 800 200728 6 la_data_out[122]
port 625 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 la_data_out[123]
port 626 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 la_data_out[124]
port 627 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 la_data_out[125]
port 628 nsew signal output
rlabel metal3 s 119200 178168 120000 178288 6 la_data_out[126]
port 629 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 la_data_out[127]
port 630 nsew signal output
rlabel metal3 s 119200 96568 120000 96688 6 la_data_out[12]
port 631 nsew signal output
rlabel metal3 s 119200 13608 120000 13728 6 la_data_out[13]
port 632 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 la_data_out[14]
port 633 nsew signal output
rlabel metal2 s 88890 209200 88946 210000 6 la_data_out[15]
port 634 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 la_data_out[16]
port 635 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 la_data_out[17]
port 636 nsew signal output
rlabel metal2 s 94686 209200 94742 210000 6 la_data_out[18]
port 637 nsew signal output
rlabel metal3 s 119200 110848 120000 110968 6 la_data_out[19]
port 638 nsew signal output
rlabel metal3 s 119200 50328 120000 50448 6 la_data_out[1]
port 639 nsew signal output
rlabel metal2 s 14830 209200 14886 210000 6 la_data_out[20]
port 640 nsew signal output
rlabel metal2 s 21914 209200 21970 210000 6 la_data_out[21]
port 641 nsew signal output
rlabel metal3 s 0 149608 800 149728 6 la_data_out[22]
port 642 nsew signal output
rlabel metal3 s 119200 83648 120000 83768 6 la_data_out[23]
port 643 nsew signal output
rlabel metal3 s 119200 37408 120000 37528 6 la_data_out[24]
port 644 nsew signal output
rlabel metal2 s 95974 209200 96030 210000 6 la_data_out[25]
port 645 nsew signal output
rlabel metal3 s 119200 201288 120000 201408 6 la_data_out[26]
port 646 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[27]
port 647 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 la_data_out[28]
port 648 nsew signal output
rlabel metal3 s 119200 39448 120000 39568 6 la_data_out[29]
port 649 nsew signal output
rlabel metal2 s 111430 209200 111486 210000 6 la_data_out[2]
port 650 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_out[30]
port 651 nsew signal output
rlabel metal3 s 119200 178848 120000 178968 6 la_data_out[31]
port 652 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 la_data_out[32]
port 653 nsew signal output
rlabel metal2 s 1306 209200 1362 210000 6 la_data_out[33]
port 654 nsew signal output
rlabel metal3 s 119200 125808 120000 125928 6 la_data_out[34]
port 655 nsew signal output
rlabel metal3 s 0 170008 800 170128 6 la_data_out[35]
port 656 nsew signal output
rlabel metal3 s 119200 78208 120000 78328 6 la_data_out[36]
port 657 nsew signal output
rlabel metal3 s 119200 97928 120000 98048 6 la_data_out[37]
port 658 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 la_data_out[38]
port 659 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 la_data_out[39]
port 660 nsew signal output
rlabel metal3 s 119200 187008 120000 187128 6 la_data_out[3]
port 661 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 la_data_out[40]
port 662 nsew signal output
rlabel metal3 s 119200 166608 120000 166728 6 la_data_out[41]
port 663 nsew signal output
rlabel metal2 s 39946 209200 40002 210000 6 la_data_out[42]
port 664 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 la_data_out[43]
port 665 nsew signal output
rlabel metal3 s 119200 2048 120000 2168 6 la_data_out[44]
port 666 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 la_data_out[45]
port 667 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 la_data_out[46]
port 668 nsew signal output
rlabel metal3 s 119200 63928 120000 64048 6 la_data_out[47]
port 669 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 la_data_out[48]
port 670 nsew signal output
rlabel metal2 s 5170 209200 5226 210000 6 la_data_out[49]
port 671 nsew signal output
rlabel metal3 s 119200 158448 120000 158568 6 la_data_out[4]
port 672 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[50]
port 673 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 la_data_out[51]
port 674 nsew signal output
rlabel metal3 s 0 203328 800 203448 6 la_data_out[52]
port 675 nsew signal output
rlabel metal3 s 119200 6808 120000 6928 6 la_data_out[53]
port 676 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[54]
port 677 nsew signal output
rlabel metal3 s 119200 14288 120000 14408 6 la_data_out[55]
port 678 nsew signal output
rlabel metal2 s 119158 209200 119214 210000 6 la_data_out[56]
port 679 nsew signal output
rlabel metal3 s 119200 108808 120000 108928 6 la_data_out[57]
port 680 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 la_data_out[58]
port 681 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 la_data_out[59]
port 682 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[5]
port 683 nsew signal output
rlabel metal2 s 3238 209200 3294 210000 6 la_data_out[60]
port 684 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[61]
port 685 nsew signal output
rlabel metal3 s 0 208088 800 208208 6 la_data_out[62]
port 686 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 la_data_out[63]
port 687 nsew signal output
rlabel metal3 s 0 177488 800 177608 6 la_data_out[64]
port 688 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 la_data_out[65]
port 689 nsew signal output
rlabel metal3 s 0 184288 800 184408 6 la_data_out[66]
port 690 nsew signal output
rlabel metal3 s 0 144848 800 144968 6 la_data_out[67]
port 691 nsew signal output
rlabel metal3 s 119200 123768 120000 123888 6 la_data_out[68]
port 692 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 la_data_out[69]
port 693 nsew signal output
rlabel metal3 s 119200 29248 120000 29368 6 la_data_out[6]
port 694 nsew signal output
rlabel metal3 s 0 180208 800 180328 6 la_data_out[70]
port 695 nsew signal output
rlabel metal2 s 4526 209200 4582 210000 6 la_data_out[71]
port 696 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[72]
port 697 nsew signal output
rlabel metal3 s 0 167288 800 167408 6 la_data_out[73]
port 698 nsew signal output
rlabel metal3 s 119200 4088 120000 4208 6 la_data_out[74]
port 699 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[75]
port 700 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 la_data_out[76]
port 701 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[77]
port 702 nsew signal output
rlabel metal3 s 119200 110168 120000 110288 6 la_data_out[78]
port 703 nsew signal output
rlabel metal3 s 119200 77528 120000 77648 6 la_data_out[79]
port 704 nsew signal output
rlabel metal3 s 119200 135328 120000 135448 6 la_data_out[7]
port 705 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 la_data_out[80]
port 706 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[81]
port 707 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 la_data_out[82]
port 708 nsew signal output
rlabel metal3 s 0 123088 800 123208 6 la_data_out[83]
port 709 nsew signal output
rlabel metal2 s 34794 209200 34850 210000 6 la_data_out[84]
port 710 nsew signal output
rlabel metal3 s 119200 47608 120000 47728 6 la_data_out[85]
port 711 nsew signal output
rlabel metal2 s 54114 209200 54170 210000 6 la_data_out[86]
port 712 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 la_data_out[87]
port 713 nsew signal output
rlabel metal3 s 119200 85008 120000 85128 6 la_data_out[88]
port 714 nsew signal output
rlabel metal3 s 119200 196528 120000 196648 6 la_data_out[89]
port 715 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 la_data_out[8]
port 716 nsew signal output
rlabel metal3 s 119200 8848 120000 8968 6 la_data_out[90]
port 717 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[91]
port 718 nsew signal output
rlabel metal3 s 0 156408 800 156528 6 la_data_out[92]
port 719 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 la_data_out[93]
port 720 nsew signal output
rlabel metal3 s 119200 51688 120000 51808 6 la_data_out[94]
port 721 nsew signal output
rlabel metal2 s 11610 209200 11666 210000 6 la_data_out[95]
port 722 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_data_out[96]
port 723 nsew signal output
rlabel metal2 s 52826 209200 52882 210000 6 la_data_out[97]
port 724 nsew signal output
rlabel metal3 s 119200 36728 120000 36848 6 la_data_out[98]
port 725 nsew signal output
rlabel metal3 s 119200 146208 120000 146328 6 la_data_out[99]
port 726 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 la_data_out[9]
port 727 nsew signal output
rlabel metal2 s 9678 209200 9734 210000 6 la_oenb[0]
port 728 nsew signal input
rlabel metal3 s 119200 84328 120000 84448 6 la_oenb[100]
port 729 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[101]
port 730 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 la_oenb[102]
port 731 nsew signal input
rlabel metal2 s 49606 209200 49662 210000 6 la_oenb[103]
port 732 nsew signal input
rlabel metal3 s 119200 106088 120000 106208 6 la_oenb[104]
port 733 nsew signal input
rlabel metal2 s 16118 209200 16174 210000 6 la_oenb[105]
port 734 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[106]
port 735 nsew signal input
rlabel metal3 s 119200 198568 120000 198688 6 la_oenb[107]
port 736 nsew signal input
rlabel metal3 s 119200 24488 120000 24608 6 la_oenb[108]
port 737 nsew signal input
rlabel metal2 s 44454 209200 44510 210000 6 la_oenb[109]
port 738 nsew signal input
rlabel metal3 s 119200 195168 120000 195288 6 la_oenb[10]
port 739 nsew signal input
rlabel metal3 s 0 193808 800 193928 6 la_oenb[110]
port 740 nsew signal input
rlabel metal2 s 7746 209200 7802 210000 6 la_oenb[111]
port 741 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_oenb[112]
port 742 nsew signal input
rlabel metal2 s 97906 209200 97962 210000 6 la_oenb[113]
port 743 nsew signal input
rlabel metal3 s 119200 23128 120000 23248 6 la_oenb[114]
port 744 nsew signal input
rlabel metal3 s 119200 184288 120000 184408 6 la_oenb[115]
port 745 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_oenb[116]
port 746 nsew signal input
rlabel metal3 s 0 181568 800 181688 6 la_oenb[117]
port 747 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 la_oenb[118]
port 748 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 la_oenb[119]
port 749 nsew signal input
rlabel metal2 s 64418 209200 64474 210000 6 la_oenb[11]
port 750 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 la_oenb[120]
port 751 nsew signal input
rlabel metal3 s 119200 87728 120000 87848 6 la_oenb[121]
port 752 nsew signal input
rlabel metal3 s 119200 191088 120000 191208 6 la_oenb[122]
port 753 nsew signal input
rlabel metal3 s 119200 3408 120000 3528 6 la_oenb[123]
port 754 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oenb[124]
port 755 nsew signal input
rlabel metal3 s 0 194488 800 194608 6 la_oenb[125]
port 756 nsew signal input
rlabel metal2 s 90822 209200 90878 210000 6 la_oenb[126]
port 757 nsew signal input
rlabel metal3 s 119200 142128 120000 142248 6 la_oenb[127]
port 758 nsew signal input
rlabel metal3 s 119200 171368 120000 171488 6 la_oenb[12]
port 759 nsew signal input
rlabel metal3 s 119200 38768 120000 38888 6 la_oenb[13]
port 760 nsew signal input
rlabel metal3 s 0 688 800 808 6 la_oenb[14]
port 761 nsew signal input
rlabel metal2 s 118514 209200 118570 210000 6 la_oenb[15]
port 762 nsew signal input
rlabel metal3 s 0 196528 800 196648 6 la_oenb[16]
port 763 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 la_oenb[17]
port 764 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_oenb[18]
port 765 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 la_oenb[19]
port 766 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 la_oenb[1]
port 767 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 la_oenb[20]
port 768 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[21]
port 769 nsew signal input
rlabel metal3 s 119200 102688 120000 102808 6 la_oenb[22]
port 770 nsew signal input
rlabel metal2 s 77298 209200 77354 210000 6 la_oenb[23]
port 771 nsew signal input
rlabel metal3 s 119200 154368 120000 154488 6 la_oenb[24]
port 772 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_oenb[25]
port 773 nsew signal input
rlabel metal3 s 119200 140088 120000 140208 6 la_oenb[26]
port 774 nsew signal input
rlabel metal3 s 119200 10888 120000 11008 6 la_oenb[27]
port 775 nsew signal input
rlabel metal2 s 43166 209200 43222 210000 6 la_oenb[28]
port 776 nsew signal input
rlabel metal3 s 119200 688 120000 808 6 la_oenb[29]
port 777 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 la_oenb[2]
port 778 nsew signal input
rlabel metal2 s 66994 209200 67050 210000 6 la_oenb[30]
port 779 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 la_oenb[31]
port 780 nsew signal input
rlabel metal2 s 18 209200 74 210000 6 la_oenb[32]
port 781 nsew signal input
rlabel metal2 s 70214 209200 70270 210000 6 la_oenb[33]
port 782 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 la_oenb[34]
port 783 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 la_oenb[35]
port 784 nsew signal input
rlabel metal3 s 119200 82288 120000 82408 6 la_oenb[36]
port 785 nsew signal input
rlabel metal3 s 119200 131928 120000 132048 6 la_oenb[37]
port 786 nsew signal input
rlabel metal3 s 119200 180888 120000 181008 6 la_oenb[38]
port 787 nsew signal input
rlabel metal3 s 0 184968 800 185088 6 la_oenb[39]
port 788 nsew signal input
rlabel metal3 s 119200 23808 120000 23928 6 la_oenb[3]
port 789 nsew signal input
rlabel metal2 s 106278 209200 106334 210000 6 la_oenb[40]
port 790 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 la_oenb[41]
port 791 nsew signal input
rlabel metal2 s 57334 209200 57390 210000 6 la_oenb[42]
port 792 nsew signal input
rlabel metal2 s 89534 209200 89590 210000 6 la_oenb[43]
port 793 nsew signal input
rlabel metal3 s 119200 53048 120000 53168 6 la_oenb[44]
port 794 nsew signal input
rlabel metal2 s 87602 209200 87658 210000 6 la_oenb[45]
port 795 nsew signal input
rlabel metal3 s 119200 45568 120000 45688 6 la_oenb[46]
port 796 nsew signal input
rlabel metal3 s 119200 78888 120000 79008 6 la_oenb[47]
port 797 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_oenb[48]
port 798 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[49]
port 799 nsew signal input
rlabel metal3 s 119200 57128 120000 57248 6 la_oenb[4]
port 800 nsew signal input
rlabel metal3 s 119200 124448 120000 124568 6 la_oenb[50]
port 801 nsew signal input
rlabel metal2 s 108854 209200 108910 210000 6 la_oenb[51]
port 802 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 la_oenb[52]
port 803 nsew signal input
rlabel metal3 s 0 189048 800 189168 6 la_oenb[53]
port 804 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 la_oenb[54]
port 805 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[55]
port 806 nsew signal input
rlabel metal2 s 91466 209200 91522 210000 6 la_oenb[56]
port 807 nsew signal input
rlabel metal3 s 119200 74808 120000 74928 6 la_oenb[57]
port 808 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 la_oenb[58]
port 809 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_oenb[59]
port 810 nsew signal input
rlabel metal2 s 114006 209200 114062 210000 6 la_oenb[5]
port 811 nsew signal input
rlabel metal2 s 24490 209200 24546 210000 6 la_oenb[60]
port 812 nsew signal input
rlabel metal2 s 14186 209200 14242 210000 6 la_oenb[61]
port 813 nsew signal input
rlabel metal2 s 46386 209200 46442 210000 6 la_oenb[62]
port 814 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_oenb[63]
port 815 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 la_oenb[64]
port 816 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_oenb[65]
port 817 nsew signal input
rlabel metal3 s 0 207408 800 207528 6 la_oenb[66]
port 818 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 la_oenb[67]
port 819 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 la_oenb[68]
port 820 nsew signal input
rlabel metal3 s 119200 40128 120000 40248 6 la_oenb[69]
port 821 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oenb[6]
port 822 nsew signal input
rlabel metal3 s 119200 99288 120000 99408 6 la_oenb[70]
port 823 nsew signal input
rlabel metal2 s 18050 209200 18106 210000 6 la_oenb[71]
port 824 nsew signal input
rlabel metal3 s 119200 116968 120000 117088 6 la_oenb[72]
port 825 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 la_oenb[73]
port 826 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 la_oenb[74]
port 827 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[75]
port 828 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oenb[76]
port 829 nsew signal input
rlabel metal3 s 0 208768 800 208888 6 la_oenb[77]
port 830 nsew signal input
rlabel metal3 s 119200 44888 120000 45008 6 la_oenb[78]
port 831 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_oenb[79]
port 832 nsew signal input
rlabel metal3 s 119200 32648 120000 32768 6 la_oenb[7]
port 833 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 la_oenb[80]
port 834 nsew signal input
rlabel metal2 s 104346 209200 104402 210000 6 la_oenb[81]
port 835 nsew signal input
rlabel metal3 s 119200 36048 120000 36168 6 la_oenb[82]
port 836 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 la_oenb[83]
port 837 nsew signal input
rlabel metal3 s 119200 80928 120000 81048 6 la_oenb[84]
port 838 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 la_oenb[85]
port 839 nsew signal input
rlabel metal3 s 0 187008 800 187128 6 la_oenb[86]
port 840 nsew signal input
rlabel metal3 s 119200 189728 120000 189848 6 la_oenb[87]
port 841 nsew signal input
rlabel metal3 s 119200 31968 120000 32088 6 la_oenb[88]
port 842 nsew signal input
rlabel metal2 s 22558 209200 22614 210000 6 la_oenb[89]
port 843 nsew signal input
rlabel metal3 s 119200 102008 120000 102128 6 la_oenb[8]
port 844 nsew signal input
rlabel metal3 s 0 175448 800 175568 6 la_oenb[90]
port 845 nsew signal input
rlabel metal3 s 119200 64608 120000 64728 6 la_oenb[91]
port 846 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 la_oenb[92]
port 847 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_oenb[93]
port 848 nsew signal input
rlabel metal3 s 119200 181568 120000 181688 6 la_oenb[94]
port 849 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_oenb[95]
port 850 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 la_oenb[96]
port 851 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[97]
port 852 nsew signal input
rlabel metal3 s 119200 67328 120000 67448 6 la_oenb[98]
port 853 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 la_oenb[99]
port 854 nsew signal input
rlabel metal2 s 27710 209200 27766 210000 6 la_oenb[9]
port 855 nsew signal input
rlabel metal2 s 101126 209200 101182 210000 6 user_irq[0]
port 856 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 user_irq[1]
port 857 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 user_irq[2]
port 858 nsew signal output
rlabel metal4 s 4208 2128 4528 207856 6 vccd1
port 859 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 207856 6 vccd1
port 859 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 207856 6 vccd1
port 859 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 207856 6 vccd1
port 859 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 207856 6 vssd1
port 860 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 207856 6 vssd1
port 860 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 207856 6 vssd1
port 860 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 207856 6 vssd1
port 860 nsew ground bidirectional
rlabel metal3 s 119200 109488 120000 109608 6 wb_clk_i
port 861 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 wb_rst_i
port 862 nsew signal input
rlabel metal3 s 119200 143488 120000 143608 6 wbs_ack_o
port 863 nsew signal output
rlabel metal3 s 0 206728 800 206848 6 wbs_adr_i[0]
port 864 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 wbs_adr_i[10]
port 865 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 wbs_adr_i[11]
port 866 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[12]
port 867 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 wbs_adr_i[13]
port 868 nsew signal input
rlabel metal2 s 113362 209200 113418 210000 6 wbs_adr_i[14]
port 869 nsew signal input
rlabel metal3 s 119200 204008 120000 204128 6 wbs_adr_i[15]
port 870 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 wbs_adr_i[16]
port 871 nsew signal input
rlabel metal3 s 119200 189048 120000 189168 6 wbs_adr_i[17]
port 872 nsew signal input
rlabel metal3 s 119200 131248 120000 131368 6 wbs_adr_i[18]
port 873 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 wbs_adr_i[19]
port 874 nsew signal input
rlabel metal2 s 2594 209200 2650 210000 6 wbs_adr_i[1]
port 875 nsew signal input
rlabel metal2 s 56046 209200 56102 210000 6 wbs_adr_i[20]
port 876 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 wbs_adr_i[21]
port 877 nsew signal input
rlabel metal3 s 119200 30608 120000 30728 6 wbs_adr_i[22]
port 878 nsew signal input
rlabel metal3 s 119200 111528 120000 111648 6 wbs_adr_i[23]
port 879 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 wbs_adr_i[24]
port 880 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 wbs_adr_i[25]
port 881 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[26]
port 882 nsew signal input
rlabel metal3 s 0 160488 800 160608 6 wbs_adr_i[27]
port 883 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wbs_adr_i[28]
port 884 nsew signal input
rlabel metal2 s 83094 209200 83150 210000 6 wbs_adr_i[29]
port 885 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 wbs_adr_i[2]
port 886 nsew signal input
rlabel metal2 s 39302 209200 39358 210000 6 wbs_adr_i[30]
port 887 nsew signal input
rlabel metal3 s 119200 144848 120000 144968 6 wbs_adr_i[31]
port 888 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 wbs_adr_i[3]
port 889 nsew signal input
rlabel metal2 s 37370 209200 37426 210000 6 wbs_adr_i[4]
port 890 nsew signal input
rlabel metal3 s 119200 15648 120000 15768 6 wbs_adr_i[5]
port 891 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 wbs_adr_i[6]
port 892 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[7]
port 893 nsew signal input
rlabel metal3 s 119200 61888 120000 62008 6 wbs_adr_i[8]
port 894 nsew signal input
rlabel metal3 s 119200 112888 120000 113008 6 wbs_adr_i[9]
port 895 nsew signal input
rlabel metal3 s 0 169328 800 169448 6 wbs_cyc_i
port 896 nsew signal input
rlabel metal2 s 105634 209200 105690 210000 6 wbs_dat_i[0]
port 897 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 wbs_dat_i[10]
port 898 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 wbs_dat_i[11]
port 899 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 wbs_dat_i[12]
port 900 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[13]
port 901 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[14]
port 902 nsew signal input
rlabel metal3 s 119200 155728 120000 155848 6 wbs_dat_i[15]
port 903 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 wbs_dat_i[16]
port 904 nsew signal input
rlabel metal2 s 32862 209200 32918 210000 6 wbs_dat_i[17]
port 905 nsew signal input
rlabel metal2 s 76010 209200 76066 210000 6 wbs_dat_i[18]
port 906 nsew signal input
rlabel metal3 s 0 129888 800 130008 6 wbs_dat_i[19]
port 907 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 wbs_dat_i[1]
port 908 nsew signal input
rlabel metal3 s 119200 168648 120000 168768 6 wbs_dat_i[20]
port 909 nsew signal input
rlabel metal2 s 83738 209200 83794 210000 6 wbs_dat_i[21]
port 910 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 wbs_dat_i[22]
port 911 nsew signal input
rlabel metal3 s 119200 199248 120000 199368 6 wbs_dat_i[23]
port 912 nsew signal input
rlabel metal3 s 119200 116288 120000 116408 6 wbs_dat_i[24]
port 913 nsew signal input
rlabel metal3 s 119200 8 120000 128 6 wbs_dat_i[25]
port 914 nsew signal input
rlabel metal2 s 65706 209200 65762 210000 6 wbs_dat_i[26]
port 915 nsew signal input
rlabel metal3 s 0 172728 800 172848 6 wbs_dat_i[27]
port 916 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wbs_dat_i[28]
port 917 nsew signal input
rlabel metal3 s 119200 164568 120000 164688 6 wbs_dat_i[29]
port 918 nsew signal input
rlabel metal3 s 119200 21768 120000 21888 6 wbs_dat_i[2]
port 919 nsew signal input
rlabel metal3 s 119200 107448 120000 107568 6 wbs_dat_i[30]
port 920 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 wbs_dat_i[31]
port 921 nsew signal input
rlabel metal3 s 119200 59848 120000 59968 6 wbs_dat_i[3]
port 922 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[4]
port 923 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 wbs_dat_i[5]
port 924 nsew signal input
rlabel metal3 s 119200 130568 120000 130688 6 wbs_dat_i[6]
port 925 nsew signal input
rlabel metal2 s 65062 209200 65118 210000 6 wbs_dat_i[7]
port 926 nsew signal input
rlabel metal2 s 117870 209200 117926 210000 6 wbs_dat_i[8]
port 927 nsew signal input
rlabel metal3 s 119200 60528 120000 60648 6 wbs_dat_i[9]
port 928 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[0]
port 929 nsew signal output
rlabel metal3 s 119200 152328 120000 152448 6 wbs_dat_o[10]
port 930 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[11]
port 931 nsew signal output
rlabel metal2 s 115938 209200 115994 210000 6 wbs_dat_o[12]
port 932 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 wbs_dat_o[13]
port 933 nsew signal output
rlabel metal3 s 119200 70728 120000 70848 6 wbs_dat_o[14]
port 934 nsew signal output
rlabel metal2 s 57978 209200 58034 210000 6 wbs_dat_o[15]
port 935 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 wbs_dat_o[16]
port 936 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 wbs_dat_o[17]
port 937 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 wbs_dat_o[18]
port 938 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 939 nsew signal output
rlabel metal3 s 119200 11568 120000 11688 6 wbs_dat_o[1]
port 940 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 wbs_dat_o[20]
port 941 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 wbs_dat_o[21]
port 942 nsew signal output
rlabel metal3 s 0 199248 800 199368 6 wbs_dat_o[22]
port 943 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_o[23]
port 944 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_o[24]
port 945 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[25]
port 946 nsew signal output
rlabel metal2 s 32218 209200 32274 210000 6 wbs_dat_o[26]
port 947 nsew signal output
rlabel metal3 s 0 206048 800 206168 6 wbs_dat_o[27]
port 948 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 wbs_dat_o[28]
port 949 nsew signal output
rlabel metal2 s 62486 209200 62542 210000 6 wbs_dat_o[29]
port 950 nsew signal output
rlabel metal3 s 119200 93848 120000 93968 6 wbs_dat_o[2]
port 951 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 wbs_dat_o[30]
port 952 nsew signal output
rlabel metal3 s 119200 177488 120000 177608 6 wbs_dat_o[31]
port 953 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[3]
port 954 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 wbs_dat_o[4]
port 955 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 wbs_dat_o[5]
port 956 nsew signal output
rlabel metal3 s 119200 170008 120000 170128 6 wbs_dat_o[6]
port 957 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 wbs_dat_o[7]
port 958 nsew signal output
rlabel metal2 s 61198 209200 61254 210000 6 wbs_dat_o[8]
port 959 nsew signal output
rlabel metal2 s 59910 209200 59966 210000 6 wbs_dat_o[9]
port 960 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 wbs_sel_i[0]
port 961 nsew signal input
rlabel metal3 s 0 182928 800 183048 6 wbs_sel_i[1]
port 962 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 wbs_sel_i[2]
port 963 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 wbs_sel_i[3]
port 964 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 wbs_stb_i
port 965 nsew signal input
rlabel metal3 s 119200 125128 120000 125248 6 wbs_we_i
port 966 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 210000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11671236
string GDS_FILE /root/hellochip/openlane/rvj1_caravel_soc/runs/22_09_13_01_33/results/signoff/rvj1_caravel_soc.magic.gds
string GDS_START 503236
<< end >>

