magic
tech sky130B
magscale 1 2
timestamp 1663004136
<< viali >>
rect 36645 27625 36679 27659
rect 2697 27557 2731 27591
rect 5273 27557 5307 27591
rect 7757 27557 7791 27591
rect 8493 27557 8527 27591
rect 9137 27557 9171 27591
rect 14289 27557 14323 27591
rect 14933 27557 14967 27591
rect 15577 27557 15611 27591
rect 18061 27557 18095 27591
rect 18613 27557 18647 27591
rect 20085 27557 20119 27591
rect 20637 27557 20671 27591
rect 22017 27557 22051 27591
rect 22569 27557 22603 27591
rect 24593 27557 24627 27591
rect 25329 27557 25363 27591
rect 27169 27557 27203 27591
rect 27813 27557 27847 27591
rect 29745 27557 29779 27591
rect 33517 27557 33551 27591
rect 34069 27557 34103 27591
rect 34897 27557 34931 27591
rect 35541 27557 35575 27591
rect 36093 27557 36127 27591
rect 37473 27557 37507 27591
rect 38117 27557 38151 27591
rect 38761 27557 38795 27591
rect 39865 27557 39899 27591
rect 40693 27557 40727 27591
rect 42625 27557 42659 27591
rect 43269 27557 43303 27591
rect 43821 27557 43855 27591
rect 45201 27557 45235 27591
rect 45845 27557 45879 27591
rect 46489 27557 46523 27591
rect 49065 27557 49099 27591
rect 51089 27557 51123 27591
rect 52745 27557 52779 27591
rect 56149 27557 56183 27591
rect 56793 27557 56827 27591
rect 57897 27557 57931 27591
rect 59369 27557 59403 27591
rect 60473 27557 60507 27591
rect 61485 27557 61519 27591
rect 61945 27557 61979 27591
rect 63049 27557 63083 27591
rect 65625 27557 65659 27591
rect 66177 27557 66211 27591
rect 66729 27557 66763 27591
rect 69673 27557 69707 27591
rect 71329 27557 71363 27591
rect 71881 27557 71915 27591
rect 72433 27557 72467 27591
rect 74273 27557 74307 27591
rect 74825 27557 74859 27591
rect 76849 27557 76883 27591
rect 77401 27557 77435 27591
rect 82001 27557 82035 27591
rect 83657 27557 83691 27591
rect 85313 27557 85347 27591
rect 86233 27557 86267 27591
rect 6377 27489 6411 27523
rect 11621 27489 11655 27523
rect 23121 27489 23155 27523
rect 30849 27489 30883 27523
rect 32413 27489 32447 27523
rect 87429 27489 87463 27523
rect 1409 27421 1443 27455
rect 2237 27421 2271 27455
rect 2881 27421 2915 27455
rect 3801 27421 3835 27455
rect 4721 27421 4755 27455
rect 5457 27421 5491 27455
rect 6653 27421 6687 27455
rect 7941 27421 7975 27455
rect 9321 27421 9355 27455
rect 10241 27421 10275 27455
rect 10517 27421 10551 27455
rect 11897 27421 11931 27455
rect 12817 27421 12851 27455
rect 13093 27421 13127 27455
rect 14473 27421 14507 27455
rect 15117 27421 15151 27455
rect 15761 27421 15795 27455
rect 16681 27421 16715 27455
rect 16957 27421 16991 27455
rect 18245 27421 18279 27455
rect 18797 27421 18831 27455
rect 19625 27421 19659 27455
rect 20269 27421 20303 27455
rect 20821 27421 20855 27455
rect 21373 27421 21407 27455
rect 22201 27421 22235 27455
rect 22753 27421 22787 27455
rect 23397 27421 23431 27455
rect 24777 27421 24811 27455
rect 25513 27421 25547 27455
rect 25973 27421 26007 27455
rect 27353 27421 27387 27455
rect 27997 27421 28031 27455
rect 28549 27421 28583 27455
rect 29101 27421 29135 27455
rect 29929 27421 29963 27455
rect 31125 27421 31159 27455
rect 32137 27421 32171 27455
rect 33701 27421 33735 27455
rect 34253 27421 34287 27455
rect 35081 27421 35115 27455
rect 35725 27421 35759 27455
rect 36277 27421 36311 27455
rect 36829 27421 36863 27455
rect 37657 27421 37691 27455
rect 38301 27421 38335 27455
rect 38945 27421 38979 27455
rect 40049 27421 40083 27455
rect 40877 27421 40911 27455
rect 41429 27421 41463 27455
rect 41981 27421 42015 27455
rect 42809 27421 42843 27455
rect 43453 27421 43487 27455
rect 44005 27421 44039 27455
rect 44557 27421 44591 27455
rect 45385 27421 45419 27455
rect 46029 27421 46063 27455
rect 46673 27421 46707 27455
rect 48605 27421 48639 27455
rect 49249 27421 49283 27455
rect 50537 27421 50571 27455
rect 51273 27421 51307 27455
rect 51825 27421 51859 27455
rect 52929 27421 52963 27455
rect 53573 27421 53607 27455
rect 53849 27421 53883 27455
rect 56333 27421 56367 27455
rect 56977 27421 57011 27455
rect 58081 27421 58115 27455
rect 58817 27421 58851 27455
rect 59553 27421 59587 27455
rect 60657 27421 60691 27455
rect 61301 27421 61335 27455
rect 62129 27421 62163 27455
rect 63233 27421 63267 27455
rect 63877 27421 63911 27455
rect 64153 27421 64187 27455
rect 65809 27421 65843 27455
rect 66361 27421 66395 27455
rect 66913 27421 66947 27455
rect 67465 27421 67499 27455
rect 68569 27421 68603 27455
rect 69305 27421 69339 27455
rect 69857 27421 69891 27455
rect 70961 27421 70995 27455
rect 71513 27421 71547 27455
rect 72065 27421 72099 27455
rect 72617 27421 72651 27455
rect 73721 27421 73755 27455
rect 74457 27421 74491 27455
rect 75009 27421 75043 27455
rect 76297 27421 76331 27455
rect 76481 27421 76515 27455
rect 77033 27421 77067 27455
rect 77585 27421 77619 27455
rect 78873 27421 78907 27455
rect 79425 27421 79459 27455
rect 80069 27421 80103 27455
rect 81449 27421 81483 27455
rect 82185 27421 82219 27455
rect 82553 27421 82587 27455
rect 83841 27421 83875 27455
rect 84393 27421 84427 27455
rect 85129 27421 85163 27455
rect 86417 27421 86451 27455
rect 86785 27421 86819 27455
rect 87705 27421 87739 27455
rect 1593 27285 1627 27319
rect 2053 27285 2087 27319
rect 3985 27285 4019 27319
rect 4813 27285 4847 27319
rect 9689 27285 9723 27319
rect 19441 27285 19475 27319
rect 21189 27285 21223 27319
rect 26065 27285 26099 27319
rect 28365 27285 28399 27319
rect 28917 27285 28951 27319
rect 41245 27285 41279 27319
rect 41797 27285 41831 27319
rect 44373 27285 44407 27319
rect 48421 27285 48455 27319
rect 50629 27285 50663 27319
rect 51641 27285 51675 27319
rect 58909 27285 58943 27319
rect 67281 27285 67315 27319
rect 68661 27285 68695 27319
rect 69121 27285 69155 27319
rect 70777 27285 70811 27319
rect 73813 27285 73847 27319
rect 78965 27285 78999 27319
rect 79609 27285 79643 27319
rect 80253 27285 80287 27319
rect 81541 27285 81575 27319
rect 82737 27285 82771 27319
rect 84209 27285 84243 27319
rect 86969 27285 87003 27319
rect 2605 27081 2639 27115
rect 3157 27081 3191 27115
rect 3985 27081 4019 27115
rect 7297 27081 7331 27115
rect 10425 27081 10459 27115
rect 13645 27081 13679 27115
rect 19809 27081 19843 27115
rect 20361 27081 20395 27115
rect 32965 27081 32999 27115
rect 37933 27081 37967 27115
rect 38301 27081 38335 27115
rect 40233 27081 40267 27115
rect 40693 27081 40727 27115
rect 42717 27081 42751 27115
rect 52929 27081 52963 27115
rect 53665 27081 53699 27115
rect 56149 27081 56183 27115
rect 58817 27081 58851 27115
rect 60657 27081 60691 27115
rect 64337 27081 64371 27115
rect 64889 27081 64923 27115
rect 65441 27081 65475 27115
rect 68845 27081 68879 27115
rect 70133 27081 70167 27115
rect 73353 27081 73387 27115
rect 74641 27081 74675 27115
rect 75469 27081 75503 27115
rect 79701 27081 79735 27115
rect 86325 27081 86359 27115
rect 86877 27081 86911 27115
rect 1777 27013 1811 27047
rect 6745 27013 6779 27047
rect 39313 27013 39347 27047
rect 39497 27013 39531 27047
rect 2329 26945 2363 26979
rect 2789 26945 2823 26979
rect 3341 26945 3375 26979
rect 4169 26945 4203 26979
rect 7481 26945 7515 26979
rect 10609 26945 10643 26979
rect 12357 26945 12391 26979
rect 13829 26945 13863 26979
rect 14749 26945 14783 26979
rect 17049 26945 17083 26979
rect 19533 26945 19567 26979
rect 19993 26945 20027 26979
rect 20545 26945 20579 26979
rect 24133 26945 24167 26979
rect 26341 26945 26375 26979
rect 27629 26945 27663 26979
rect 27813 26945 27847 26979
rect 28365 26945 28399 26979
rect 29193 26945 29227 26979
rect 30389 26945 30423 26979
rect 32321 26945 32355 26979
rect 33149 26945 33183 26979
rect 38117 26945 38151 26979
rect 38393 26945 38427 26979
rect 40049 26945 40083 26979
rect 40325 26945 40359 26979
rect 40877 26945 40911 26979
rect 42901 26945 42935 26979
rect 44741 26945 44775 26979
rect 49893 26945 49927 26979
rect 53113 26969 53147 27003
rect 53849 26945 53883 26979
rect 54217 26945 54251 26979
rect 56333 26945 56367 26979
rect 58449 26945 58483 26979
rect 59001 26945 59035 26979
rect 60841 26945 60875 26979
rect 64521 26945 64555 26979
rect 65073 26945 65107 26979
rect 65625 26945 65659 26979
rect 69029 26945 69063 26979
rect 70317 26945 70351 26979
rect 73537 26945 73571 26979
rect 74825 26945 74859 26979
rect 75653 26945 75687 26979
rect 77401 26945 77435 26979
rect 77585 26945 77619 26979
rect 79885 26945 79919 26979
rect 84669 26945 84703 26979
rect 85221 26945 85255 26979
rect 86509 26945 86543 26979
rect 87061 26945 87095 26979
rect 26157 26877 26191 26911
rect 27445 26877 27479 26911
rect 30665 26877 30699 26911
rect 32137 26877 32171 26911
rect 54493 26877 54527 26911
rect 77217 26877 77251 26911
rect 87429 26877 87463 26911
rect 87705 26877 87739 26911
rect 1961 26809 1995 26843
rect 6929 26809 6963 26843
rect 14565 26809 14599 26843
rect 28181 26809 28215 26843
rect 29009 26809 29043 26843
rect 39865 26809 39899 26843
rect 44925 26809 44959 26843
rect 12541 26741 12575 26775
rect 16865 26741 16899 26775
rect 23949 26741 23983 26775
rect 26525 26741 26559 26775
rect 32505 26741 32539 26775
rect 32873 26741 32907 26775
rect 49709 26741 49743 26775
rect 58265 26741 58299 26775
rect 75101 26741 75135 26775
rect 85405 26741 85439 26775
rect 2881 26537 2915 26571
rect 87429 26537 87463 26571
rect 26709 26469 26743 26503
rect 27261 26469 27295 26503
rect 40969 26469 41003 26503
rect 40601 26401 40635 26435
rect 1409 26333 1443 26367
rect 1685 26333 1719 26367
rect 3065 26333 3099 26367
rect 3985 26333 4019 26367
rect 26893 26333 26927 26367
rect 27445 26333 27479 26367
rect 29561 26333 29595 26367
rect 29745 26333 29779 26367
rect 30665 26333 30699 26367
rect 31033 26333 31067 26367
rect 31309 26333 31343 26367
rect 40785 26333 40819 26367
rect 87061 26333 87095 26367
rect 87613 26333 87647 26367
rect 87981 26333 88015 26367
rect 29929 26265 29963 26299
rect 3801 26197 3835 26231
rect 30481 26197 30515 26231
rect 86877 26197 86911 26231
rect 88165 26197 88199 26231
rect 1409 25993 1443 26027
rect 2789 25993 2823 26027
rect 44005 25993 44039 26027
rect 86785 25993 86819 26027
rect 87521 25993 87555 26027
rect 88073 25993 88107 26027
rect 27905 25925 27939 25959
rect 1593 25857 1627 25891
rect 2697 25857 2731 25891
rect 2973 25857 3007 25891
rect 27353 25857 27387 25891
rect 43821 25857 43855 25891
rect 87705 25857 87739 25891
rect 88257 25857 88291 25891
rect 2237 25789 2271 25823
rect 43637 25789 43671 25823
rect 2513 25721 2547 25755
rect 27445 25653 27479 25687
rect 87153 25653 87187 25687
rect 1409 25245 1443 25279
rect 1685 25245 1719 25279
rect 87889 25177 87923 25211
rect 87981 25109 88015 25143
rect 88257 24769 88291 24803
rect 1409 24701 1443 24735
rect 1685 24701 1719 24735
rect 88073 24565 88107 24599
rect 88257 24157 88291 24191
rect 88073 24021 88107 24055
rect 86785 23817 86819 23851
rect 1777 23681 1811 23715
rect 21833 23681 21867 23715
rect 86969 23681 87003 23715
rect 88257 23681 88291 23715
rect 1961 23545 1995 23579
rect 21925 23477 21959 23511
rect 86417 23477 86451 23511
rect 88073 23477 88107 23511
rect 73537 22593 73571 22627
rect 88073 22593 88107 22627
rect 1593 22525 1627 22559
rect 73353 22389 73387 22423
rect 88165 22389 88199 22423
rect 1593 21981 1627 22015
rect 88257 21981 88291 22015
rect 1409 21845 1443 21879
rect 87705 21845 87739 21879
rect 88073 21845 88107 21879
rect 4169 21641 4203 21675
rect 1409 21505 1443 21539
rect 3985 21505 4019 21539
rect 88257 21505 88291 21539
rect 3801 21437 3835 21471
rect 1593 21301 1627 21335
rect 87705 21301 87739 21335
rect 88073 21301 88107 21335
rect 87705 20961 87739 20995
rect 1593 20893 1627 20927
rect 87429 20893 87463 20927
rect 1409 20757 1443 20791
rect 1961 20757 1995 20791
rect 22201 20553 22235 20587
rect 22569 20485 22603 20519
rect 30297 20485 30331 20519
rect 22385 20417 22419 20451
rect 22661 20417 22695 20451
rect 30113 20417 30147 20451
rect 30389 20417 30423 20451
rect 29929 20213 29963 20247
rect 1409 19805 1443 19839
rect 1685 19805 1719 19839
rect 88257 19805 88291 19839
rect 87705 19669 87739 19703
rect 88073 19669 88107 19703
rect 26249 19397 26283 19431
rect 1777 19329 1811 19363
rect 26065 19329 26099 19363
rect 26341 19329 26375 19363
rect 56517 19329 56551 19363
rect 56701 19329 56735 19363
rect 56793 19329 56827 19363
rect 88257 19329 88291 19363
rect 56333 19261 56367 19295
rect 1961 19193 1995 19227
rect 55689 19193 55723 19227
rect 56057 19193 56091 19227
rect 25881 19125 25915 19159
rect 57161 19125 57195 19159
rect 88073 19125 88107 19159
rect 24593 18921 24627 18955
rect 56701 18921 56735 18955
rect 28089 18785 28123 18819
rect 28273 18785 28307 18819
rect 1593 18717 1627 18751
rect 1961 18717 1995 18751
rect 24777 18717 24811 18751
rect 24961 18717 24995 18751
rect 25053 18717 25087 18751
rect 36185 18717 36219 18751
rect 47777 18717 47811 18751
rect 56885 18717 56919 18751
rect 88257 18717 88291 18751
rect 57161 18649 57195 18683
rect 1409 18581 1443 18615
rect 27629 18581 27663 18615
rect 27997 18581 28031 18615
rect 36001 18581 36035 18615
rect 47593 18581 47627 18615
rect 57069 18581 57103 18615
rect 88073 18581 88107 18615
rect 26157 18377 26191 18411
rect 27997 18377 28031 18411
rect 28457 18377 28491 18411
rect 33977 18377 34011 18411
rect 36001 18377 36035 18411
rect 48053 18377 48087 18411
rect 48329 18377 48363 18411
rect 48973 18377 49007 18411
rect 49341 18377 49375 18411
rect 54953 18377 54987 18411
rect 55321 18377 55355 18411
rect 56149 18377 56183 18411
rect 67465 18377 67499 18411
rect 23857 18309 23891 18343
rect 24685 18309 24719 18343
rect 34437 18309 34471 18343
rect 36461 18309 36495 18343
rect 55781 18309 55815 18343
rect 69489 18309 69523 18343
rect 1593 18241 1627 18275
rect 24593 18241 24627 18275
rect 26065 18241 26099 18275
rect 27629 18241 27663 18275
rect 28365 18241 28399 18275
rect 29285 18241 29319 18275
rect 33609 18241 33643 18275
rect 34345 18241 34379 18275
rect 35633 18241 35667 18275
rect 36369 18241 36403 18275
rect 41889 18241 41923 18275
rect 45017 18241 45051 18275
rect 47869 18241 47903 18275
rect 48789 18241 48823 18275
rect 49065 18241 49099 18275
rect 54585 18241 54619 18275
rect 55137 18241 55171 18275
rect 55413 18241 55447 18275
rect 55965 18241 55999 18275
rect 56241 18241 56275 18275
rect 67373 18241 67407 18275
rect 69397 18241 69431 18275
rect 70501 18241 70535 18275
rect 70593 18241 70627 18275
rect 24777 18173 24811 18207
rect 26341 18173 26375 18207
rect 28641 18173 28675 18207
rect 34529 18173 34563 18207
rect 36645 18173 36679 18207
rect 47685 18173 47719 18207
rect 67557 18173 67591 18207
rect 69581 18173 69615 18207
rect 70685 18173 70719 18207
rect 48605 18105 48639 18139
rect 1409 18037 1443 18071
rect 24225 18037 24259 18071
rect 25697 18037 25731 18071
rect 27445 18037 27479 18071
rect 29101 18037 29135 18071
rect 33425 18037 33459 18071
rect 35449 18037 35483 18071
rect 41705 18037 41739 18071
rect 44833 18037 44867 18071
rect 54401 18037 54435 18071
rect 67005 18037 67039 18071
rect 69029 18037 69063 18071
rect 70133 18037 70167 18071
rect 48789 17833 48823 17867
rect 50169 17833 50203 17867
rect 24777 17765 24811 17799
rect 36093 17765 36127 17799
rect 41337 17765 41371 17799
rect 42901 17765 42935 17799
rect 44557 17765 44591 17799
rect 45477 17765 45511 17799
rect 47501 17765 47535 17799
rect 64981 17765 65015 17799
rect 67925 17765 67959 17799
rect 25329 17697 25363 17731
rect 27353 17697 27387 17731
rect 27629 17697 27663 17731
rect 28733 17697 28767 17731
rect 32137 17697 32171 17731
rect 32321 17697 32355 17731
rect 40785 17697 40819 17731
rect 40969 17697 41003 17731
rect 43269 17697 43303 17731
rect 55689 17697 55723 17731
rect 61669 17697 61703 17731
rect 68569 17697 68603 17731
rect 69949 17697 69983 17731
rect 24961 17629 24995 17663
rect 25605 17629 25639 17663
rect 33425 17629 33459 17663
rect 33609 17629 33643 17663
rect 33885 17629 33919 17663
rect 34713 17629 34747 17663
rect 36553 17629 36587 17663
rect 36809 17629 36843 17663
rect 41521 17629 41555 17663
rect 43177 17629 43211 17663
rect 44281 17629 44315 17663
rect 44373 17629 44407 17663
rect 45661 17629 45695 17663
rect 45937 17629 45971 17663
rect 46949 17629 46983 17663
rect 47225 17629 47259 17663
rect 47369 17629 47403 17663
rect 48145 17629 48179 17663
rect 48421 17629 48455 17663
rect 48973 17629 49007 17663
rect 49157 17629 49191 17663
rect 49249 17629 49283 17663
rect 50353 17629 50387 17663
rect 50629 17629 50663 17663
rect 53297 17629 53331 17663
rect 53573 17629 53607 17663
rect 54125 17629 54159 17663
rect 54401 17629 54435 17663
rect 55321 17629 55355 17663
rect 55505 17629 55539 17663
rect 56057 17629 56091 17663
rect 56241 17629 56275 17663
rect 56425 17629 56459 17663
rect 56977 17629 57011 17663
rect 58725 17629 58759 17663
rect 58863 17629 58897 17663
rect 59001 17629 59035 17663
rect 59139 17629 59173 17663
rect 60013 17629 60047 17663
rect 62405 17629 62439 17663
rect 62681 17629 62715 17663
rect 65165 17629 65199 17663
rect 65625 17629 65659 17663
rect 68109 17629 68143 17663
rect 68845 17629 68879 17663
rect 70961 17629 70995 17663
rect 26985 17561 27019 17595
rect 34980 17561 35014 17595
rect 40693 17561 40727 17595
rect 41788 17561 41822 17595
rect 47133 17561 47167 17595
rect 60841 17561 60875 17595
rect 61485 17561 61519 17595
rect 62221 17561 62255 17595
rect 65870 17561 65904 17595
rect 31677 17493 31711 17527
rect 32045 17493 32079 17527
rect 33793 17493 33827 17527
rect 37933 17493 37967 17527
rect 40325 17493 40359 17527
rect 45845 17493 45879 17527
rect 47961 17493 47995 17527
rect 48329 17493 48363 17527
rect 50537 17493 50571 17527
rect 53395 17493 53429 17527
rect 53481 17493 53515 17527
rect 53941 17493 53975 17527
rect 54309 17493 54343 17527
rect 56793 17493 56827 17527
rect 59277 17493 59311 17527
rect 59829 17493 59863 17527
rect 60933 17493 60967 17527
rect 62589 17493 62623 17527
rect 67005 17493 67039 17527
rect 70777 17493 70811 17527
rect 23213 17289 23247 17323
rect 24041 17289 24075 17323
rect 27528 17221 27562 17255
rect 32597 17221 32631 17255
rect 35716 17221 35750 17255
rect 37841 17221 37875 17255
rect 42901 17221 42935 17255
rect 53665 17221 53699 17255
rect 54392 17221 54426 17255
rect 58725 17221 58759 17255
rect 59921 17221 59955 17255
rect 63141 17221 63175 17255
rect 65165 17221 65199 17255
rect 1777 17153 1811 17187
rect 23949 17153 23983 17187
rect 24961 17153 24995 17187
rect 26249 17153 26283 17187
rect 31677 17153 31711 17187
rect 32505 17153 32539 17187
rect 33609 17153 33643 17187
rect 33793 17153 33827 17187
rect 33885 17153 33919 17187
rect 37657 17153 37691 17187
rect 38209 17153 38243 17187
rect 39589 17153 39623 17187
rect 39856 17153 39890 17187
rect 41245 17153 41279 17187
rect 41797 17153 41831 17187
rect 42809 17153 42843 17187
rect 43545 17153 43579 17187
rect 43729 17153 43763 17187
rect 43821 17153 43855 17187
rect 44833 17153 44867 17187
rect 45100 17153 45134 17187
rect 46581 17153 46615 17187
rect 46765 17153 46799 17187
rect 46949 17153 46983 17187
rect 47041 17153 47075 17187
rect 47593 17153 47627 17187
rect 47849 17153 47883 17187
rect 49709 17153 49743 17187
rect 49893 17153 49927 17187
rect 49985 17153 50019 17187
rect 50813 17153 50847 17187
rect 50997 17153 51031 17187
rect 51549 17153 51583 17187
rect 52929 17153 52963 17187
rect 53481 17153 53515 17187
rect 53757 17153 53791 17187
rect 53849 17153 53883 17187
rect 56333 17153 56367 17187
rect 57897 17153 57931 17187
rect 58081 17153 58115 17187
rect 58173 17153 58207 17187
rect 58909 17153 58943 17187
rect 59093 17153 59127 17187
rect 59185 17153 59219 17187
rect 59737 17153 59771 17187
rect 60289 17153 60323 17187
rect 60545 17153 60579 17187
rect 62129 17153 62163 17187
rect 63325 17153 63359 17187
rect 63509 17153 63543 17187
rect 63601 17153 63635 17187
rect 64521 17153 64555 17187
rect 64889 17153 64923 17187
rect 64981 17153 65015 17187
rect 66177 17153 66211 17187
rect 66913 17153 66947 17187
rect 67005 17153 67039 17187
rect 68937 17153 68971 17187
rect 69949 17153 69983 17187
rect 73813 17153 73847 17187
rect 88257 17153 88291 17187
rect 1961 17085 1995 17119
rect 24225 17085 24259 17119
rect 24685 17085 24719 17119
rect 27261 17085 27295 17119
rect 32781 17085 32815 17119
rect 35449 17085 35483 17119
rect 41613 17085 41647 17119
rect 42993 17085 43027 17119
rect 50629 17085 50663 17119
rect 54125 17085 54159 17119
rect 56149 17085 56183 17119
rect 59553 17085 59587 17119
rect 66269 17085 66303 17119
rect 66453 17085 66487 17119
rect 69673 17085 69707 17119
rect 71053 17085 71087 17119
rect 23581 17017 23615 17051
rect 32137 17017 32171 17051
rect 40969 17017 41003 17051
rect 42441 17017 42475 17051
rect 46213 17017 46247 17051
rect 48973 17017 49007 17051
rect 49525 17017 49559 17051
rect 53113 17017 53147 17051
rect 54033 17017 54067 17051
rect 55873 17017 55907 17051
rect 65809 17017 65843 17051
rect 68753 17017 68787 17051
rect 73629 17017 73663 17051
rect 88073 17017 88107 17051
rect 24777 16949 24811 16983
rect 26065 16949 26099 16983
rect 28641 16949 28675 16983
rect 31493 16949 31527 16983
rect 33425 16949 33459 16983
rect 36829 16949 36863 16983
rect 38301 16949 38335 16983
rect 41981 16949 42015 16983
rect 43545 16949 43579 16983
rect 50353 16949 50387 16983
rect 51365 16949 51399 16983
rect 55505 16949 55539 16983
rect 56517 16949 56551 16983
rect 57897 16949 57931 16983
rect 61669 16949 61703 16983
rect 62221 16949 62255 16983
rect 64337 16949 64371 16983
rect 65533 16949 65567 16983
rect 20085 16745 20119 16779
rect 21189 16745 21223 16779
rect 62313 16745 62347 16779
rect 64705 16745 64739 16779
rect 28641 16677 28675 16711
rect 40049 16677 40083 16711
rect 46581 16677 46615 16711
rect 47777 16677 47811 16711
rect 52929 16677 52963 16711
rect 57805 16677 57839 16711
rect 20913 16609 20947 16643
rect 26065 16609 26099 16643
rect 28273 16609 28307 16643
rect 33609 16609 33643 16643
rect 33701 16609 33735 16643
rect 36369 16609 36403 16643
rect 36553 16609 36587 16643
rect 50169 16609 50203 16643
rect 54309 16609 54343 16643
rect 55321 16609 55355 16643
rect 59369 16609 59403 16643
rect 65625 16609 65659 16643
rect 68385 16609 68419 16643
rect 71145 16609 71179 16643
rect 71513 16609 71547 16643
rect 1593 16541 1627 16575
rect 20269 16541 20303 16575
rect 20545 16541 20579 16575
rect 21373 16541 21407 16575
rect 21649 16541 21683 16575
rect 25697 16541 25731 16575
rect 26332 16541 26366 16575
rect 28457 16541 28491 16575
rect 30849 16541 30883 16575
rect 31217 16541 31251 16575
rect 35357 16541 35391 16575
rect 36277 16541 36311 16575
rect 38577 16541 38611 16575
rect 40233 16541 40267 16575
rect 41521 16541 41555 16575
rect 41889 16541 41923 16575
rect 43821 16541 43855 16575
rect 44097 16541 44131 16575
rect 46857 16541 46891 16575
rect 47225 16541 47259 16575
rect 47409 16541 47443 16575
rect 47598 16541 47632 16575
rect 50436 16541 50470 16575
rect 52377 16541 52411 16575
rect 52561 16541 52595 16575
rect 52750 16541 52784 16575
rect 53389 16541 53423 16575
rect 53573 16541 53607 16575
rect 53757 16541 53791 16575
rect 54493 16541 54527 16575
rect 54769 16541 54803 16575
rect 57253 16541 57287 16575
rect 58081 16541 58115 16575
rect 58633 16541 58667 16575
rect 58725 16541 58759 16575
rect 60565 16541 60599 16575
rect 61117 16541 61151 16575
rect 61393 16541 61427 16575
rect 62497 16541 62531 16575
rect 62773 16541 62807 16575
rect 63233 16541 63267 16575
rect 63877 16541 63911 16575
rect 64061 16541 64095 16575
rect 64889 16541 64923 16575
rect 65165 16541 65199 16575
rect 65881 16541 65915 16575
rect 70317 16541 70351 16575
rect 71329 16541 71363 16575
rect 88257 16541 88291 16575
rect 20453 16473 20487 16507
rect 21557 16473 21591 16507
rect 31484 16473 31518 16507
rect 33517 16473 33551 16507
rect 38025 16473 38059 16507
rect 42134 16473 42168 16507
rect 46581 16473 46615 16507
rect 47501 16473 47535 16507
rect 52653 16473 52687 16507
rect 53665 16473 53699 16507
rect 54677 16473 54711 16507
rect 55588 16473 55622 16507
rect 57805 16473 57839 16507
rect 58449 16473 58483 16507
rect 59185 16473 59219 16507
rect 59829 16473 59863 16507
rect 60013 16473 60047 16507
rect 62681 16473 62715 16507
rect 68652 16473 68686 16507
rect 1409 16405 1443 16439
rect 25513 16405 25547 16439
rect 27445 16405 27479 16439
rect 30665 16405 30699 16439
rect 32597 16405 32631 16439
rect 33149 16405 33183 16439
rect 35449 16405 35483 16439
rect 35909 16405 35943 16439
rect 38117 16405 38151 16439
rect 38669 16405 38703 16439
rect 41337 16405 41371 16439
rect 43269 16405 43303 16439
rect 43637 16405 43671 16439
rect 44005 16405 44039 16439
rect 46765 16405 46799 16439
rect 51549 16405 51583 16439
rect 53941 16405 53975 16439
rect 56701 16405 56735 16439
rect 57069 16405 57103 16439
rect 57989 16405 58023 16439
rect 58547 16405 58581 16439
rect 60657 16405 60691 16439
rect 63325 16405 63359 16439
rect 65073 16405 65107 16439
rect 67005 16405 67039 16439
rect 69765 16405 69799 16439
rect 70133 16405 70167 16439
rect 88073 16405 88107 16439
rect 2973 16201 3007 16235
rect 21833 16201 21867 16235
rect 24409 16201 24443 16235
rect 30389 16201 30423 16235
rect 31493 16201 31527 16235
rect 34713 16201 34747 16235
rect 35633 16201 35667 16235
rect 36093 16201 36127 16235
rect 43185 16201 43219 16235
rect 51641 16201 51675 16235
rect 65809 16201 65843 16235
rect 69397 16201 69431 16235
rect 71237 16201 71271 16235
rect 71973 16201 72007 16235
rect 12909 16133 12943 16167
rect 25320 16133 25354 16167
rect 33578 16133 33612 16167
rect 42809 16133 42843 16167
rect 43821 16133 43855 16167
rect 44649 16133 44683 16167
rect 46489 16133 46523 16167
rect 46581 16133 46615 16167
rect 51273 16133 51307 16167
rect 52929 16133 52963 16167
rect 57161 16133 57195 16167
rect 58909 16133 58943 16167
rect 59737 16133 59771 16167
rect 64705 16133 64739 16167
rect 65441 16133 65475 16167
rect 3157 16065 3191 16099
rect 12725 16065 12759 16099
rect 22017 16065 22051 16099
rect 22201 16065 22235 16099
rect 22293 16065 22327 16099
rect 24317 16065 24351 16099
rect 25053 16065 25087 16099
rect 27241 16065 27275 16099
rect 29009 16065 29043 16099
rect 30297 16065 30331 16099
rect 31125 16065 31159 16099
rect 31677 16065 31711 16099
rect 32689 16065 32723 16099
rect 32873 16065 32907 16099
rect 32965 16065 32999 16099
rect 33333 16065 33367 16099
rect 35265 16065 35299 16099
rect 36001 16065 36035 16099
rect 37473 16065 37507 16099
rect 37657 16065 37691 16099
rect 37749 16065 37783 16099
rect 41521 16065 41555 16099
rect 42625 16065 42659 16099
rect 42901 16065 42935 16099
rect 42998 16065 43032 16099
rect 43637 16065 43671 16099
rect 43913 16065 43947 16099
rect 44010 16065 44044 16099
rect 44833 16065 44867 16099
rect 45017 16065 45051 16099
rect 45109 16065 45143 16099
rect 45845 16065 45879 16099
rect 46305 16065 46339 16099
rect 46678 16065 46712 16099
rect 47593 16065 47627 16099
rect 47777 16065 47811 16099
rect 47869 16065 47903 16099
rect 48237 16065 48271 16099
rect 48421 16065 48455 16099
rect 48513 16065 48547 16099
rect 50077 16065 50111 16099
rect 50261 16065 50295 16099
rect 50353 16065 50387 16099
rect 51457 16065 51491 16099
rect 51733 16065 51767 16099
rect 52745 16065 52779 16099
rect 53021 16065 53055 16099
rect 53165 16065 53199 16099
rect 53849 16065 53883 16099
rect 54125 16065 54159 16099
rect 55137 16065 55171 16099
rect 55404 16065 55438 16099
rect 56977 16065 57011 16099
rect 58081 16065 58115 16099
rect 58265 16065 58299 16099
rect 58357 16065 58391 16099
rect 58725 16065 58759 16099
rect 59001 16065 59035 16099
rect 59145 16065 59179 16099
rect 59921 16065 59955 16099
rect 60105 16065 60139 16099
rect 60197 16065 60231 16099
rect 60841 16065 60875 16099
rect 62129 16065 62163 16099
rect 62313 16065 62347 16099
rect 63049 16065 63083 16099
rect 63233 16065 63267 16099
rect 63417 16065 63451 16099
rect 63969 16065 64003 16099
rect 64521 16065 64555 16099
rect 64797 16065 64831 16099
rect 64889 16065 64923 16099
rect 65625 16065 65659 16099
rect 65901 16065 65935 16099
rect 68477 16065 68511 16099
rect 69213 16065 69247 16099
rect 69489 16065 69523 16099
rect 70124 16065 70158 16099
rect 72065 16065 72099 16099
rect 73813 16065 73847 16099
rect 88257 16065 88291 16099
rect 12541 15997 12575 16031
rect 24593 15997 24627 16031
rect 26985 15997 27019 16031
rect 28825 15997 28859 16031
rect 29193 15997 29227 16031
rect 36185 15997 36219 16031
rect 61117 15997 61151 16031
rect 69857 15997 69891 16031
rect 72157 15997 72191 16031
rect 30941 15929 30975 15963
rect 47593 15929 47627 15963
rect 48237 15929 48271 15963
rect 53297 15929 53331 15963
rect 58081 15929 58115 15963
rect 68569 15929 68603 15963
rect 73629 15929 73663 15963
rect 23949 15861 23983 15895
rect 26433 15861 26467 15895
rect 28365 15861 28399 15895
rect 32505 15861 32539 15895
rect 35081 15861 35115 15895
rect 37289 15861 37323 15895
rect 41613 15861 41647 15895
rect 44189 15861 44223 15895
rect 45661 15861 45695 15895
rect 46857 15861 46891 15895
rect 49893 15861 49927 15895
rect 56517 15861 56551 15895
rect 59277 15861 59311 15895
rect 63785 15861 63819 15895
rect 65073 15861 65107 15895
rect 69213 15861 69247 15895
rect 71605 15861 71639 15895
rect 88073 15861 88107 15895
rect 27445 15657 27479 15691
rect 32413 15657 32447 15691
rect 44097 15657 44131 15691
rect 45385 15657 45419 15691
rect 47501 15657 47535 15691
rect 50169 15657 50203 15691
rect 51641 15657 51675 15691
rect 55321 15657 55355 15691
rect 60013 15657 60047 15691
rect 65625 15657 65659 15691
rect 70777 15657 70811 15691
rect 71881 15657 71915 15691
rect 47133 15589 47167 15623
rect 49433 15589 49467 15623
rect 68477 15589 68511 15623
rect 72525 15589 72559 15623
rect 27905 15521 27939 15555
rect 28089 15521 28123 15555
rect 30389 15521 30423 15555
rect 32781 15521 32815 15555
rect 36093 15521 36127 15555
rect 38393 15521 38427 15555
rect 38577 15521 38611 15555
rect 41521 15521 41555 15555
rect 45753 15521 45787 15555
rect 48329 15521 48363 15555
rect 53481 15521 53515 15555
rect 53757 15521 53791 15555
rect 58265 15521 58299 15555
rect 58633 15521 58667 15555
rect 60565 15521 60599 15555
rect 60841 15521 60875 15555
rect 62957 15521 62991 15555
rect 71237 15521 71271 15555
rect 71421 15521 71455 15555
rect 1409 15453 1443 15487
rect 20545 15453 20579 15487
rect 20821 15453 20855 15487
rect 23121 15453 23155 15487
rect 25237 15453 25271 15487
rect 25605 15453 25639 15487
rect 27813 15453 27847 15487
rect 31033 15453 31067 15487
rect 33037 15453 33071 15487
rect 35081 15453 35115 15487
rect 35265 15453 35299 15487
rect 35357 15453 35391 15487
rect 42349 15453 42383 15487
rect 42717 15453 42751 15487
rect 45109 15453 45143 15487
rect 45201 15453 45235 15487
rect 46009 15453 46043 15487
rect 47685 15453 47719 15487
rect 47961 15453 47995 15487
rect 48513 15453 48547 15487
rect 48789 15453 48823 15487
rect 49249 15453 49283 15487
rect 50445 15453 50479 15487
rect 51273 15453 51307 15487
rect 51641 15453 51675 15487
rect 51917 15453 51951 15487
rect 52285 15453 52319 15487
rect 52561 15453 52595 15487
rect 55321 15453 55355 15487
rect 55597 15453 55631 15487
rect 55965 15453 55999 15487
rect 56241 15453 56275 15487
rect 57897 15453 57931 15487
rect 58081 15453 58115 15487
rect 62037 15453 62071 15487
rect 63224 15453 63258 15487
rect 64889 15453 64923 15487
rect 65809 15453 65843 15487
rect 65993 15453 66027 15487
rect 66085 15453 66119 15487
rect 68017 15453 68051 15487
rect 68385 15453 68419 15487
rect 68937 15453 68971 15487
rect 69204 15453 69238 15487
rect 72065 15453 72099 15487
rect 72433 15453 72467 15487
rect 20729 15385 20763 15419
rect 25850 15385 25884 15419
rect 28917 15385 28951 15419
rect 30205 15385 30239 15419
rect 31278 15385 31312 15419
rect 34897 15385 34931 15419
rect 36360 15385 36394 15419
rect 38301 15385 38335 15419
rect 41337 15385 41371 15419
rect 41981 15385 42015 15419
rect 42984 15385 43018 15419
rect 47869 15385 47903 15419
rect 50169 15385 50203 15419
rect 51825 15385 51859 15419
rect 55505 15385 55539 15419
rect 57253 15385 57287 15419
rect 58878 15385 58912 15419
rect 61853 15385 61887 15419
rect 62313 15385 62347 15419
rect 88073 15385 88107 15419
rect 1593 15317 1627 15351
rect 20361 15317 20395 15351
rect 23213 15317 23247 15351
rect 25053 15317 25087 15351
rect 26985 15317 27019 15351
rect 29009 15317 29043 15351
rect 34161 15317 34195 15351
rect 37473 15317 37507 15351
rect 37933 15317 37967 15351
rect 48697 15317 48731 15351
rect 50353 15317 50387 15351
rect 51089 15317 51123 15351
rect 57345 15317 57379 15351
rect 62221 15317 62255 15351
rect 64337 15317 64371 15351
rect 64705 15317 64739 15351
rect 67833 15317 67867 15351
rect 70317 15317 70351 15351
rect 71145 15317 71179 15351
rect 88165 15317 88199 15351
rect 18613 15113 18647 15147
rect 20085 15113 20119 15147
rect 20453 15113 20487 15147
rect 22293 15113 22327 15147
rect 27445 15113 27479 15147
rect 30481 15113 30515 15147
rect 32137 15113 32171 15147
rect 32597 15113 32631 15147
rect 33241 15113 33275 15147
rect 33609 15113 33643 15147
rect 53481 15113 53515 15147
rect 63785 15113 63819 15147
rect 65717 15113 65751 15147
rect 66453 15113 66487 15147
rect 67281 15113 67315 15147
rect 69305 15113 69339 15147
rect 23949 15045 23983 15079
rect 28733 15045 28767 15079
rect 28825 15045 28859 15079
rect 32505 15045 32539 15079
rect 36001 15045 36035 15079
rect 49700 15045 49734 15079
rect 51457 15045 51491 15079
rect 52193 15045 52227 15079
rect 55045 15045 55079 15079
rect 55229 15045 55263 15079
rect 56425 15045 56459 15079
rect 62221 15045 62255 15079
rect 63417 15045 63451 15079
rect 68937 15045 68971 15079
rect 18797 14977 18831 15011
rect 18981 14977 19015 15011
rect 19073 14977 19107 15011
rect 20269 14977 20303 15011
rect 20545 14977 20579 15011
rect 20913 14977 20947 15011
rect 22109 14977 22143 15011
rect 22385 14977 22419 15011
rect 22753 14977 22787 15011
rect 23673 14977 23707 15011
rect 23765 14977 23799 15011
rect 24317 14977 24351 15011
rect 24501 14977 24535 15011
rect 25053 14977 25087 15011
rect 25309 14977 25343 15011
rect 27353 14977 27387 15011
rect 28549 14977 28583 15011
rect 29193 14977 29227 15011
rect 30389 14977 30423 15011
rect 31309 14977 31343 15011
rect 33425 14977 33459 15011
rect 33701 14977 33735 15011
rect 34069 14977 34103 15011
rect 34621 14977 34655 15011
rect 35265 14977 35299 15011
rect 35449 14977 35483 15011
rect 35541 14977 35575 15011
rect 36185 14977 36219 15011
rect 36369 14977 36403 15011
rect 36461 14977 36495 15011
rect 37545 14977 37579 15011
rect 39661 14977 39695 15011
rect 41153 14977 41187 15011
rect 41705 14977 41739 15011
rect 42441 14977 42475 15011
rect 44373 14977 44407 15011
rect 44557 14977 44591 15011
rect 44741 14977 44775 15011
rect 45293 14977 45327 15011
rect 48237 14977 48271 15011
rect 48697 14977 48731 15011
rect 51181 14977 51215 15011
rect 52009 14977 52043 15011
rect 53297 14977 53331 15011
rect 53573 14977 53607 15011
rect 54309 14977 54343 15011
rect 54493 14977 54527 15011
rect 55321 14977 55355 15011
rect 55781 14977 55815 15011
rect 56609 14977 56643 15011
rect 56793 14977 56827 15011
rect 56885 14977 56919 15011
rect 57437 14977 57471 15011
rect 59277 14977 59311 15011
rect 59461 14977 59495 15011
rect 60749 14977 60783 15011
rect 62037 14977 62071 15011
rect 62313 14977 62347 15011
rect 62405 14977 62439 15011
rect 63601 14977 63635 15011
rect 63877 14977 63911 15011
rect 64337 14977 64371 15011
rect 64604 14977 64638 15011
rect 66269 14977 66303 15011
rect 66545 14977 66579 15011
rect 67097 14977 67131 15011
rect 67373 14977 67407 15011
rect 68753 14977 68787 15011
rect 69025 14977 69059 15011
rect 69121 14977 69155 15011
rect 69673 14977 69707 15011
rect 69949 14977 69983 15011
rect 71697 14977 71731 15011
rect 21925 14909 21959 14943
rect 27537 14909 27571 14943
rect 29469 14909 29503 14943
rect 31401 14909 31435 14943
rect 31585 14909 31619 14943
rect 32781 14909 32815 14943
rect 37289 14909 37323 14943
rect 39405 14909 39439 14943
rect 41245 14909 41279 14943
rect 43085 14909 43119 14943
rect 43361 14909 43395 14943
rect 45661 14909 45695 14943
rect 45937 14909 45971 14943
rect 48881 14909 48915 14943
rect 49433 14909 49467 14943
rect 58081 14909 58115 14943
rect 58403 14909 58437 14943
rect 60473 14909 60507 14943
rect 66913 14909 66947 14943
rect 71053 14909 71087 14943
rect 41889 14841 41923 14875
rect 45109 14841 45143 14875
rect 50813 14841 50847 14875
rect 51273 14841 51307 14875
rect 53113 14841 53147 14875
rect 55045 14841 55079 14875
rect 57253 14841 57287 14875
rect 21189 14773 21223 14807
rect 21373 14773 21407 14807
rect 23029 14773 23063 14807
rect 23213 14773 23247 14807
rect 24317 14773 24351 14807
rect 26433 14773 26467 14807
rect 26985 14773 27019 14807
rect 28365 14773 28399 14807
rect 30941 14773 30975 14807
rect 34161 14773 34195 14807
rect 34713 14773 34747 14807
rect 35265 14773 35299 14807
rect 38669 14773 38703 14807
rect 40785 14773 40819 14807
rect 42625 14773 42659 14807
rect 48053 14773 48087 14807
rect 51181 14773 51215 14807
rect 54677 14773 54711 14807
rect 55873 14773 55907 14807
rect 59645 14773 59679 14807
rect 62589 14773 62623 14807
rect 66085 14773 66119 14807
rect 71881 14773 71915 14807
rect 23213 14569 23247 14603
rect 26157 14569 26191 14603
rect 37105 14569 37139 14603
rect 37749 14569 37783 14603
rect 52193 14569 52227 14603
rect 28089 14501 28123 14535
rect 33701 14501 33735 14535
rect 35817 14501 35851 14535
rect 39221 14501 39255 14535
rect 41245 14501 41279 14535
rect 44189 14501 44223 14535
rect 45569 14501 45603 14535
rect 46213 14501 46247 14535
rect 61025 14501 61059 14535
rect 70317 14501 70351 14535
rect 70777 14501 70811 14535
rect 72249 14501 72283 14535
rect 22661 14433 22695 14467
rect 30849 14433 30883 14467
rect 32045 14433 32079 14467
rect 36553 14433 36587 14467
rect 39865 14433 39899 14467
rect 41613 14433 41647 14467
rect 43269 14433 43303 14467
rect 43453 14433 43487 14467
rect 45109 14433 45143 14467
rect 48881 14433 48915 14467
rect 53849 14433 53883 14467
rect 55689 14433 55723 14467
rect 58265 14433 58299 14467
rect 58633 14433 58667 14467
rect 61485 14433 61519 14467
rect 68937 14433 68971 14467
rect 71329 14433 71363 14467
rect 1593 14365 1627 14399
rect 20545 14365 20579 14399
rect 20637 14365 20671 14399
rect 21281 14365 21315 14399
rect 21373 14365 21407 14399
rect 21557 14365 21591 14399
rect 21649 14365 21683 14399
rect 22201 14365 22235 14399
rect 22293 14365 22327 14399
rect 23121 14365 23155 14399
rect 24409 14365 24443 14399
rect 24777 14365 24811 14399
rect 25789 14365 25823 14399
rect 26341 14365 26375 14399
rect 26709 14365 26743 14399
rect 28733 14365 28767 14399
rect 28917 14365 28951 14399
rect 29009 14365 29043 14399
rect 30021 14365 30055 14399
rect 30665 14365 30699 14399
rect 31309 14365 31343 14399
rect 33701 14365 33735 14399
rect 33977 14365 34011 14399
rect 34989 14365 35023 14399
rect 35173 14365 35207 14399
rect 35725 14365 35759 14399
rect 36093 14365 36127 14399
rect 36461 14365 36495 14399
rect 37289 14365 37323 14399
rect 37933 14365 37967 14399
rect 38301 14365 38335 14399
rect 38485 14365 38519 14399
rect 39405 14365 39439 14399
rect 40121 14365 40155 14399
rect 41889 14365 41923 14399
rect 43913 14365 43947 14399
rect 44189 14365 44223 14399
rect 45017 14365 45051 14399
rect 45753 14365 45787 14399
rect 46121 14365 46155 14399
rect 47593 14365 47627 14399
rect 47777 14365 47811 14399
rect 48331 14365 48365 14399
rect 49157 14365 49191 14399
rect 50537 14365 50571 14399
rect 50721 14365 50755 14399
rect 51089 14365 51123 14399
rect 51273 14365 51307 14399
rect 52101 14365 52135 14399
rect 52653 14365 52687 14399
rect 52929 14365 52963 14399
rect 54125 14365 54159 14399
rect 55321 14365 55355 14399
rect 58081 14365 58115 14399
rect 60473 14365 60507 14399
rect 60657 14365 60691 14399
rect 60893 14365 60927 14399
rect 61669 14365 61703 14399
rect 61945 14365 61979 14399
rect 62497 14365 62531 14399
rect 62681 14365 62715 14399
rect 62773 14365 62807 14399
rect 63785 14365 63819 14399
rect 63969 14365 64003 14399
rect 64061 14365 64095 14399
rect 64429 14365 64463 14399
rect 64701 14365 64735 14399
rect 64797 14365 64831 14399
rect 66453 14365 66487 14399
rect 66720 14365 66754 14399
rect 68385 14365 68419 14399
rect 71145 14365 71179 14399
rect 71237 14365 71271 14399
rect 22569 14297 22603 14331
rect 24593 14297 24627 14331
rect 24685 14297 24719 14331
rect 26954 14297 26988 14331
rect 28549 14297 28583 14331
rect 32290 14297 32324 14331
rect 34345 14297 34379 14331
rect 35817 14297 35851 14331
rect 43177 14297 43211 14331
rect 56793 14297 56827 14331
rect 57437 14297 57471 14331
rect 57621 14297 57655 14331
rect 58878 14297 58912 14331
rect 60749 14297 60783 14331
rect 61853 14297 61887 14331
rect 64613 14297 64647 14331
rect 69204 14297 69238 14331
rect 71881 14297 71915 14331
rect 72065 14297 72099 14331
rect 88073 14297 88107 14331
rect 1409 14229 1443 14263
rect 21097 14229 21131 14263
rect 22017 14229 22051 14263
rect 23581 14229 23615 14263
rect 24961 14229 24995 14263
rect 25605 14229 25639 14263
rect 30113 14229 30147 14263
rect 31401 14229 31435 14263
rect 33425 14229 33459 14263
rect 33885 14229 33919 14263
rect 35357 14229 35391 14263
rect 36001 14229 36035 14263
rect 38669 14229 38703 14263
rect 42809 14229 42843 14263
rect 47685 14229 47719 14263
rect 48421 14229 48455 14263
rect 51181 14229 51215 14263
rect 56885 14229 56919 14263
rect 60013 14229 60047 14263
rect 62313 14229 62347 14263
rect 63601 14229 63635 14263
rect 64981 14229 65015 14263
rect 67833 14229 67867 14263
rect 68477 14229 68511 14263
rect 88165 14229 88199 14263
rect 2881 14025 2915 14059
rect 19441 14025 19475 14059
rect 21005 14025 21039 14059
rect 24777 14025 24811 14059
rect 28549 14025 28583 14059
rect 29101 14025 29135 14059
rect 34253 14025 34287 14059
rect 35650 14025 35684 14059
rect 36093 14025 36127 14059
rect 39313 14025 39347 14059
rect 40601 14025 40635 14059
rect 51181 14025 51215 14059
rect 57995 14025 58029 14059
rect 64245 14025 64279 14059
rect 65073 14025 65107 14059
rect 67557 14025 67591 14059
rect 70777 14025 70811 14059
rect 72433 14025 72467 14059
rect 73905 14025 73939 14059
rect 26157 13957 26191 13991
rect 28089 13957 28123 13991
rect 29009 13957 29043 13991
rect 31493 13957 31527 13991
rect 33517 13957 33551 13991
rect 37473 13957 37507 13991
rect 41061 13957 41095 13991
rect 46397 13957 46431 13991
rect 57437 13957 57471 13991
rect 61950 13957 61984 13991
rect 63049 13957 63083 13991
rect 63417 13957 63451 13991
rect 1593 13889 1627 13923
rect 3065 13889 3099 13923
rect 18153 13889 18187 13923
rect 18981 13889 19015 13923
rect 19809 13889 19843 13923
rect 20913 13889 20947 13923
rect 21097 13889 21131 13923
rect 23029 13889 23063 13923
rect 23213 13889 23247 13923
rect 23857 13889 23891 13923
rect 24685 13889 24719 13923
rect 25237 13889 25271 13923
rect 25329 13889 25363 13923
rect 25973 13889 26007 13923
rect 26249 13889 26283 13923
rect 26341 13889 26375 13923
rect 27353 13889 27387 13923
rect 30205 13889 30239 13923
rect 31309 13889 31343 13923
rect 32505 13889 32539 13923
rect 32689 13889 32723 13923
rect 33241 13889 33275 13923
rect 34437 13889 34471 13923
rect 34805 13889 34839 13923
rect 35081 13889 35115 13923
rect 35265 13889 35299 13923
rect 35357 13889 35391 13923
rect 35477 13889 35511 13923
rect 37289 13889 37323 13923
rect 37565 13889 37599 13923
rect 37709 13889 37743 13923
rect 38301 13889 38335 13923
rect 40233 13873 40267 13907
rect 40969 13889 41003 13923
rect 41705 13889 41739 13923
rect 42625 13889 42659 13923
rect 43821 13889 43855 13923
rect 44088 13889 44122 13923
rect 45753 13889 45787 13923
rect 46581 13889 46615 13923
rect 46949 13889 46983 13923
rect 48217 13889 48251 13923
rect 50057 13889 50091 13923
rect 51733 13889 51767 13923
rect 52929 13889 52963 13923
rect 53196 13889 53230 13923
rect 55137 13889 55171 13923
rect 57069 13889 57103 13923
rect 57253 13889 57287 13923
rect 57897 13889 57931 13923
rect 58081 13889 58115 13923
rect 58182 13889 58216 13923
rect 59093 13889 59127 13923
rect 61669 13889 61703 13923
rect 61853 13889 61887 13923
rect 62042 13889 62076 13923
rect 63233 13889 63267 13923
rect 63509 13889 63543 13923
rect 64061 13889 64095 13923
rect 64337 13889 64371 13923
rect 64797 13889 64831 13923
rect 64889 13889 64923 13923
rect 67741 13893 67775 13927
rect 68201 13879 68235 13913
rect 68385 13889 68419 13923
rect 68477 13889 68511 13923
rect 68570 13895 68604 13929
rect 69653 13889 69687 13923
rect 71329 13889 71363 13923
rect 72065 13889 72099 13923
rect 72249 13889 72283 13923
rect 72525 13889 72559 13923
rect 73721 13889 73755 13923
rect 88257 13889 88291 13923
rect 18613 13821 18647 13855
rect 20269 13821 20303 13855
rect 21373 13821 21407 13855
rect 23673 13821 23707 13855
rect 23765 13821 23799 13855
rect 24133 13821 24167 13855
rect 27445 13821 27479 13855
rect 27537 13821 27571 13855
rect 39405 13821 39439 13855
rect 39589 13821 39623 13855
rect 41153 13821 41187 13855
rect 42901 13821 42935 13855
rect 45569 13821 45603 13855
rect 45937 13821 45971 13855
rect 47961 13821 47995 13855
rect 49801 13821 49835 13855
rect 51549 13821 51583 13855
rect 51917 13821 51951 13855
rect 55321 13821 55355 13855
rect 55689 13821 55723 13855
rect 55965 13821 55999 13855
rect 58817 13821 58851 13855
rect 60473 13821 60507 13855
rect 60749 13821 60783 13855
rect 69397 13821 69431 13855
rect 71237 13821 71271 13855
rect 73537 13821 73571 13855
rect 20821 13753 20855 13787
rect 22845 13753 22879 13787
rect 23581 13753 23615 13787
rect 26525 13753 26559 13787
rect 26985 13753 27019 13787
rect 28457 13753 28491 13787
rect 30389 13753 30423 13787
rect 38577 13753 38611 13787
rect 40049 13753 40083 13787
rect 41889 13753 41923 13787
rect 49341 13753 49375 13787
rect 68845 13753 68879 13787
rect 1409 13685 1443 13719
rect 18245 13685 18279 13719
rect 19165 13685 19199 13719
rect 19901 13685 19935 13719
rect 21281 13685 21315 13719
rect 22477 13685 22511 13719
rect 22753 13685 22787 13719
rect 22937 13685 22971 13719
rect 24041 13685 24075 13719
rect 25421 13685 25455 13719
rect 25605 13685 25639 13719
rect 37841 13685 37875 13719
rect 38117 13685 38151 13719
rect 38945 13685 38979 13719
rect 45201 13685 45235 13719
rect 47041 13685 47075 13719
rect 54309 13685 54343 13719
rect 62221 13685 62255 13719
rect 63877 13685 63911 13719
rect 71697 13685 71731 13719
rect 88073 13685 88107 13719
rect 20913 13481 20947 13515
rect 22109 13481 22143 13515
rect 22937 13481 22971 13515
rect 23305 13481 23339 13515
rect 23857 13481 23891 13515
rect 25697 13481 25731 13515
rect 28733 13481 28767 13515
rect 30297 13481 30331 13515
rect 37749 13481 37783 13515
rect 38945 13481 38979 13515
rect 43637 13481 43671 13515
rect 44373 13481 44407 13515
rect 50629 13481 50663 13515
rect 52009 13481 52043 13515
rect 55321 13481 55355 13515
rect 55965 13481 55999 13515
rect 60013 13481 60047 13515
rect 61853 13481 61887 13515
rect 63601 13481 63635 13515
rect 19717 13413 19751 13447
rect 19901 13413 19935 13447
rect 21373 13413 21407 13447
rect 27905 13413 27939 13447
rect 47225 13413 47259 13447
rect 49157 13413 49191 13447
rect 52469 13413 52503 13447
rect 56701 13413 56735 13447
rect 61025 13413 61059 13447
rect 67649 13413 67683 13447
rect 68293 13413 68327 13447
rect 72157 13413 72191 13447
rect 19625 13345 19659 13379
rect 21005 13345 21039 13379
rect 22477 13345 22511 13379
rect 24593 13345 24627 13379
rect 25697 13345 25731 13379
rect 31861 13345 31895 13379
rect 34713 13345 34747 13379
rect 39865 13345 39899 13379
rect 45477 13345 45511 13379
rect 45845 13345 45879 13379
rect 49065 13345 49099 13379
rect 52929 13345 52963 13379
rect 53113 13345 53147 13379
rect 1593 13277 1627 13311
rect 15025 13277 15059 13311
rect 17969 13277 18003 13311
rect 18245 13277 18279 13311
rect 19533 13277 19567 13311
rect 19717 13277 19751 13311
rect 19993 13277 20027 13311
rect 21189 13277 21223 13311
rect 22017 13277 22051 13311
rect 22845 13277 22879 13311
rect 23765 13277 23799 13311
rect 24501 13277 24535 13311
rect 25053 13277 25087 13311
rect 25881 13277 25915 13311
rect 26525 13277 26559 13311
rect 26618 13277 26652 13311
rect 26801 13277 26835 13311
rect 26893 13277 26927 13311
rect 26990 13277 27024 13311
rect 27537 13277 27571 13311
rect 28641 13277 28675 13311
rect 29561 13277 29595 13311
rect 30113 13277 30147 13311
rect 30849 13277 30883 13311
rect 31585 13277 31619 13311
rect 32965 13277 32999 13311
rect 33517 13277 33551 13311
rect 33885 13277 33919 13311
rect 34969 13277 35003 13311
rect 39129 13277 39163 13311
rect 39313 13277 39347 13311
rect 39405 13277 39439 13311
rect 40141 13277 40175 13311
rect 41429 13277 41463 13311
rect 41613 13277 41647 13311
rect 42257 13277 42291 13311
rect 44557 13277 44591 13311
rect 47593 13277 47627 13311
rect 47869 13277 47903 13311
rect 48973 13277 49007 13311
rect 49249 13277 49283 13311
rect 49433 13277 49467 13311
rect 50261 13277 50295 13311
rect 50445 13277 50479 13311
rect 51457 13277 51491 13311
rect 51825 13277 51859 13311
rect 52837 13277 52871 13311
rect 53665 13277 53699 13311
rect 55505 13277 55539 13311
rect 55873 13277 55907 13311
rect 57069 13277 57103 13311
rect 57345 13277 57379 13311
rect 58265 13277 58299 13311
rect 59461 13277 59495 13311
rect 59829 13277 59863 13311
rect 60473 13277 60507 13311
rect 60746 13277 60780 13311
rect 60846 13277 60880 13311
rect 61485 13277 61519 13311
rect 61669 13277 61703 13311
rect 62221 13277 62255 13311
rect 63969 13277 64003 13311
rect 64797 13277 64831 13311
rect 65809 13277 65843 13311
rect 67925 13277 67959 13311
rect 68569 13277 68603 13311
rect 68937 13277 68971 13311
rect 69121 13277 69155 13311
rect 69305 13277 69339 13311
rect 69857 13277 69891 13311
rect 70041 13277 70075 13311
rect 70225 13277 70259 13311
rect 70317 13277 70351 13311
rect 70777 13277 70811 13311
rect 71044 13277 71078 13311
rect 88257 13277 88291 13311
rect 20913 13209 20947 13243
rect 25605 13209 25639 13243
rect 29653 13209 29687 13243
rect 32781 13209 32815 13243
rect 33241 13209 33275 13243
rect 36461 13209 36495 13243
rect 42502 13209 42536 13243
rect 45293 13209 45327 13243
rect 46112 13209 46146 13243
rect 48789 13209 48823 13243
rect 51641 13209 51675 13243
rect 51733 13209 51767 13243
rect 53849 13209 53883 13243
rect 54309 13209 54343 13243
rect 56517 13209 56551 13243
rect 59645 13209 59679 13243
rect 59737 13209 59771 13243
rect 60657 13209 60691 13243
rect 62488 13209 62522 13243
rect 67649 13209 67683 13243
rect 68293 13209 68327 13243
rect 69213 13209 69247 13243
rect 1409 13141 1443 13175
rect 15117 13141 15151 13175
rect 25145 13141 25179 13175
rect 26065 13141 26099 13175
rect 27169 13141 27203 13175
rect 27997 13141 28031 13175
rect 30941 13141 30975 13175
rect 33149 13141 33183 13175
rect 34069 13141 34103 13175
rect 36093 13141 36127 13175
rect 41797 13141 41831 13175
rect 54401 13141 54435 13175
rect 58495 13141 58529 13175
rect 64153 13141 64187 13175
rect 64613 13141 64647 13175
rect 65625 13141 65659 13175
rect 67833 13141 67867 13175
rect 68477 13141 68511 13175
rect 69489 13141 69523 13175
rect 88073 13141 88107 13175
rect 23489 12937 23523 12971
rect 24501 12937 24535 12971
rect 25421 12937 25455 12971
rect 26433 12937 26467 12971
rect 29101 12937 29135 12971
rect 36829 12937 36863 12971
rect 38577 12937 38611 12971
rect 42671 12937 42705 12971
rect 46397 12937 46431 12971
rect 48329 12937 48363 12971
rect 52745 12937 52779 12971
rect 59277 12937 59311 12971
rect 64889 12937 64923 12971
rect 86785 12937 86819 12971
rect 23673 12869 23707 12903
rect 24961 12869 24995 12903
rect 30205 12869 30239 12903
rect 31309 12869 31343 12903
rect 34069 12869 34103 12903
rect 34805 12869 34839 12903
rect 35817 12869 35851 12903
rect 38117 12869 38151 12903
rect 39037 12869 39071 12903
rect 40601 12869 40635 12903
rect 46673 12869 46707 12903
rect 47961 12869 47995 12903
rect 48177 12869 48211 12903
rect 49709 12869 49743 12903
rect 51730 12869 51764 12903
rect 54585 12869 54619 12903
rect 56977 12869 57011 12903
rect 59829 12869 59863 12903
rect 61577 12869 61611 12903
rect 62313 12869 62347 12903
rect 63316 12869 63350 12903
rect 66453 12869 66487 12903
rect 67189 12869 67223 12903
rect 67557 12869 67591 12903
rect 1685 12801 1719 12835
rect 18613 12801 18647 12835
rect 19809 12801 19843 12835
rect 20637 12801 20671 12835
rect 24409 12801 24443 12835
rect 25145 12801 25179 12835
rect 25237 12801 25271 12835
rect 25789 12801 25823 12835
rect 26249 12801 26283 12835
rect 26525 12801 26559 12835
rect 30113 12801 30147 12835
rect 31677 12801 31711 12835
rect 32413 12801 32447 12835
rect 32597 12801 32631 12835
rect 32689 12801 32723 12835
rect 33057 12801 33091 12835
rect 33885 12801 33919 12835
rect 34161 12801 34195 12835
rect 34529 12801 34563 12835
rect 34713 12801 34747 12835
rect 34897 12801 34931 12835
rect 35541 12801 35575 12835
rect 35725 12801 35759 12835
rect 35909 12801 35943 12835
rect 36553 12801 36587 12835
rect 36645 12801 36679 12835
rect 37749 12801 37783 12835
rect 38485 12801 38519 12835
rect 41521 12801 41555 12835
rect 41705 12801 41739 12835
rect 41797 12801 41831 12835
rect 42441 12801 42475 12835
rect 44005 12801 44039 12835
rect 44557 12801 44591 12835
rect 44741 12801 44775 12835
rect 44833 12801 44867 12835
rect 45661 12801 45695 12835
rect 46581 12801 46615 12835
rect 46765 12801 46799 12835
rect 46883 12801 46917 12835
rect 47041 12801 47075 12835
rect 48789 12801 48823 12835
rect 51457 12801 51491 12835
rect 51641 12801 51675 12835
rect 51871 12801 51905 12835
rect 52929 12801 52963 12835
rect 53113 12801 53147 12835
rect 53205 12801 53239 12835
rect 53573 12801 53607 12835
rect 53757 12801 53791 12835
rect 53849 12801 53883 12835
rect 56701 12801 56735 12835
rect 56839 12801 56873 12835
rect 57069 12801 57103 12835
rect 57897 12801 57931 12835
rect 59093 12801 59127 12835
rect 59369 12801 59403 12835
rect 61945 12801 61979 12835
rect 62129 12801 62163 12835
rect 62405 12801 62439 12835
rect 65349 12801 65383 12835
rect 66269 12801 66303 12835
rect 66545 12801 66579 12835
rect 66637 12801 66671 12835
rect 67373 12801 67407 12835
rect 67649 12801 67683 12835
rect 68753 12801 68787 12835
rect 69213 12801 69247 12835
rect 69305 12801 69339 12835
rect 69489 12801 69523 12835
rect 70124 12801 70158 12835
rect 71605 12801 71639 12835
rect 71789 12801 71823 12835
rect 72341 12801 72375 12835
rect 86969 12801 87003 12835
rect 88257 12801 88291 12835
rect 1409 12733 1443 12767
rect 19073 12733 19107 12767
rect 23581 12733 23615 12767
rect 23765 12733 23799 12767
rect 24041 12733 24075 12767
rect 27445 12733 27479 12767
rect 27813 12733 27847 12767
rect 28641 12733 28675 12767
rect 30297 12733 30331 12767
rect 33701 12733 33735 12767
rect 43821 12733 43855 12767
rect 43913 12733 43947 12767
rect 44097 12733 44131 12767
rect 45570 12733 45604 12767
rect 45753 12733 45787 12767
rect 45845 12733 45879 12767
rect 49893 12733 49927 12767
rect 49985 12733 50019 12767
rect 50261 12733 50295 12767
rect 58173 12733 58207 12767
rect 63049 12733 63083 12767
rect 65073 12733 65107 12767
rect 69857 12733 69891 12767
rect 23949 12665 23983 12699
rect 26157 12665 26191 12699
rect 28089 12665 28123 12699
rect 28917 12665 28951 12699
rect 43637 12665 43671 12699
rect 51181 12665 51215 12699
rect 57253 12665 57287 12699
rect 59093 12665 59127 12699
rect 65257 12665 65291 12699
rect 68569 12665 68603 12699
rect 71973 12665 72007 12699
rect 18889 12597 18923 12631
rect 19901 12597 19935 12631
rect 20269 12597 20303 12631
rect 20729 12597 20763 12631
rect 21097 12597 21131 12631
rect 25237 12597 25271 12631
rect 26065 12597 26099 12631
rect 28273 12597 28307 12631
rect 29745 12597 29779 12631
rect 32229 12597 32263 12631
rect 33241 12597 33275 12631
rect 35081 12597 35115 12631
rect 36093 12597 36127 12631
rect 41337 12597 41371 12631
rect 44557 12597 44591 12631
rect 45385 12597 45419 12631
rect 48145 12597 48179 12631
rect 48881 12597 48915 12631
rect 52009 12597 52043 12631
rect 53573 12597 53607 12631
rect 55873 12597 55907 12631
rect 64429 12597 64463 12631
rect 66821 12597 66855 12631
rect 71237 12597 71271 12631
rect 72433 12597 72467 12631
rect 88073 12597 88107 12631
rect 20085 12393 20119 12427
rect 25789 12393 25823 12427
rect 26249 12393 26283 12427
rect 28641 12393 28675 12427
rect 30941 12393 30975 12427
rect 31585 12393 31619 12427
rect 33885 12393 33919 12427
rect 36001 12393 36035 12427
rect 39405 12393 39439 12427
rect 42349 12393 42383 12427
rect 43913 12393 43947 12427
rect 49433 12393 49467 12427
rect 53021 12393 53055 12427
rect 54033 12393 54067 12427
rect 58357 12393 58391 12427
rect 61853 12393 61887 12427
rect 64061 12393 64095 12427
rect 64889 12393 64923 12427
rect 65717 12393 65751 12427
rect 67925 12393 67959 12427
rect 69489 12393 69523 12427
rect 70041 12393 70075 12427
rect 21005 12325 21039 12359
rect 26801 12325 26835 12359
rect 28365 12325 28399 12359
rect 28917 12325 28951 12359
rect 34805 12325 34839 12359
rect 36369 12325 36403 12359
rect 45385 12325 45419 12359
rect 46305 12325 46339 12359
rect 54769 12325 54803 12359
rect 66085 12325 66119 12359
rect 72157 12325 72191 12359
rect 72525 12325 72559 12359
rect 20821 12257 20855 12291
rect 26065 12257 26099 12291
rect 27629 12257 27663 12291
rect 27813 12257 27847 12291
rect 28457 12257 28491 12291
rect 29561 12257 29595 12291
rect 32321 12257 32355 12291
rect 33517 12257 33551 12291
rect 37473 12257 37507 12291
rect 40969 12257 41003 12291
rect 42717 12257 42751 12291
rect 46489 12257 46523 12291
rect 46673 12257 46707 12291
rect 48513 12257 48547 12291
rect 50445 12257 50479 12291
rect 57253 12257 57287 12291
rect 59185 12257 59219 12291
rect 60473 12257 60507 12291
rect 64245 12257 64279 12291
rect 64429 12257 64463 12291
rect 65901 12257 65935 12291
rect 70777 12257 70811 12291
rect 19901 12189 19935 12223
rect 21005 12189 21039 12223
rect 21097 12189 21131 12223
rect 21281 12189 21315 12223
rect 25191 12189 25225 12223
rect 25431 12189 25465 12223
rect 26157 12189 26191 12223
rect 26341 12189 26375 12223
rect 26525 12189 26559 12223
rect 28549 12189 28583 12223
rect 29101 12189 29135 12223
rect 31769 12189 31803 12223
rect 32137 12189 32171 12223
rect 33149 12189 33183 12223
rect 33333 12189 33367 12223
rect 34069 12189 34103 12223
rect 34989 12189 35023 12223
rect 35725 12189 35759 12223
rect 35817 12189 35851 12223
rect 36553 12189 36587 12223
rect 36737 12189 36771 12223
rect 36829 12189 36863 12223
rect 37197 12189 37231 12223
rect 38025 12189 38059 12223
rect 38281 12189 38315 12223
rect 40049 12189 40083 12223
rect 40233 12189 40267 12223
rect 40417 12189 40451 12223
rect 42993 12189 43027 12223
rect 44097 12189 44131 12223
rect 44373 12189 44407 12223
rect 45569 12189 45603 12223
rect 45845 12189 45879 12223
rect 46581 12189 46615 12223
rect 46765 12189 46799 12223
rect 48053 12189 48087 12223
rect 48421 12189 48455 12223
rect 48605 12189 48639 12223
rect 49709 12189 49743 12223
rect 50169 12189 50203 12223
rect 51641 12189 51675 12223
rect 53481 12189 53515 12223
rect 54309 12189 54343 12223
rect 54677 12189 54711 12223
rect 55505 12189 55539 12223
rect 57437 12189 57471 12223
rect 57713 12189 57747 12223
rect 58541 12189 58575 12223
rect 58817 12189 58851 12223
rect 59461 12189 59495 12223
rect 62313 12189 62347 12223
rect 62408 12199 62442 12233
rect 63049 12189 63083 12223
rect 63233 12189 63267 12223
rect 64521 12189 64555 12223
rect 65165 12189 65199 12223
rect 66177 12189 66211 12223
rect 66545 12189 66579 12223
rect 68753 12189 68787 12223
rect 68937 12189 68971 12223
rect 70317 12189 70351 12223
rect 72709 12189 72743 12223
rect 20913 12121 20947 12155
rect 27537 12121 27571 12155
rect 27997 12121 28031 12155
rect 29806 12121 29840 12155
rect 35265 12121 35299 12155
rect 40325 12121 40359 12155
rect 41236 12121 41270 12155
rect 49433 12121 49467 12155
rect 49617 12121 49651 12155
rect 51908 12121 51942 12155
rect 54033 12121 54067 12155
rect 55750 12121 55784 12155
rect 60740 12121 60774 12155
rect 62589 12121 62623 12155
rect 64889 12121 64923 12155
rect 66812 12121 66846 12155
rect 69305 12121 69339 12155
rect 69505 12121 69539 12155
rect 70041 12121 70075 12155
rect 70225 12121 70259 12155
rect 71044 12121 71078 12155
rect 20361 12053 20395 12087
rect 24961 12053 24995 12087
rect 25329 12053 25363 12087
rect 27169 12053 27203 12087
rect 35173 12053 35207 12087
rect 40601 12053 40635 12087
rect 44281 12053 44315 12087
rect 45753 12053 45787 12087
rect 47869 12053 47903 12087
rect 53573 12053 53607 12087
rect 54217 12053 54251 12087
rect 56885 12053 56919 12087
rect 57621 12053 57655 12087
rect 58725 12053 58759 12087
rect 65073 12053 65107 12087
rect 68845 12053 68879 12087
rect 69673 12053 69707 12087
rect 24593 11849 24627 11883
rect 25421 11849 25455 11883
rect 26433 11849 26467 11883
rect 29653 11849 29687 11883
rect 30849 11849 30883 11883
rect 35817 11849 35851 11883
rect 37473 11849 37507 11883
rect 46213 11849 46247 11883
rect 46949 11849 46983 11883
rect 47593 11849 47627 11883
rect 47961 11849 47995 11883
rect 49801 11849 49835 11883
rect 51733 11849 51767 11883
rect 52101 11849 52135 11883
rect 52745 11849 52779 11883
rect 54769 11849 54803 11883
rect 55413 11849 55447 11883
rect 55873 11849 55907 11883
rect 64613 11849 64647 11883
rect 66913 11849 66947 11883
rect 70593 11849 70627 11883
rect 71237 11849 71271 11883
rect 71605 11849 71639 11883
rect 20085 11781 20119 11815
rect 26157 11781 26191 11815
rect 29745 11781 29779 11815
rect 32505 11781 32539 11815
rect 37289 11781 37323 11815
rect 44097 11781 44131 11815
rect 45100 11781 45134 11815
rect 50598 11781 50632 11815
rect 53113 11781 53147 11815
rect 54585 11781 54619 11815
rect 56977 11781 57011 11815
rect 57437 11781 57471 11815
rect 58909 11781 58943 11815
rect 63049 11781 63083 11815
rect 64429 11781 64463 11815
rect 69458 11781 69492 11815
rect 70869 11781 70903 11815
rect 1593 11713 1627 11747
rect 18797 11713 18831 11747
rect 18981 11713 19015 11747
rect 19073 11713 19107 11747
rect 19809 11713 19843 11747
rect 19901 11713 19935 11747
rect 20729 11713 20763 11747
rect 24133 11713 24167 11747
rect 25789 11713 25823 11747
rect 25882 11713 25916 11747
rect 26065 11713 26099 11747
rect 26295 11713 26329 11747
rect 31033 11713 31067 11747
rect 31493 11713 31527 11747
rect 33600 11713 33634 11747
rect 35633 11713 35667 11747
rect 35909 11713 35943 11747
rect 36461 11713 36495 11747
rect 36553 11713 36587 11747
rect 36737 11713 36771 11747
rect 37565 11713 37599 11747
rect 39497 11713 39531 11747
rect 40049 11713 40083 11747
rect 40233 11713 40267 11747
rect 41153 11713 41187 11747
rect 43913 11713 43947 11747
rect 44189 11713 44223 11747
rect 44281 11713 44315 11747
rect 46765 11713 46799 11747
rect 47041 11713 47075 11747
rect 47777 11713 47811 11747
rect 48053 11713 48087 11747
rect 49985 11713 50019 11747
rect 50353 11713 50387 11747
rect 52277 11713 52311 11747
rect 52929 11713 52963 11747
rect 53215 11713 53249 11747
rect 53757 11713 53791 11747
rect 53941 11713 53975 11747
rect 54033 11713 54067 11747
rect 54861 11713 54895 11747
rect 55229 11713 55263 11747
rect 55505 11713 55539 11747
rect 56057 11713 56091 11747
rect 57161 11713 57195 11747
rect 57345 11713 57379 11747
rect 57897 11713 57931 11747
rect 58081 11713 58115 11747
rect 58633 11713 58667 11747
rect 58817 11713 58851 11747
rect 59053 11713 59087 11747
rect 59829 11713 59863 11747
rect 60013 11713 60047 11747
rect 60105 11713 60139 11747
rect 61108 11713 61142 11747
rect 63877 11713 63911 11747
rect 64061 11713 64095 11747
rect 64705 11713 64739 11747
rect 66177 11713 66211 11747
rect 66361 11713 66395 11747
rect 66545 11713 66579 11747
rect 67097 11713 67131 11747
rect 68385 11713 68419 11747
rect 68937 11713 68971 11747
rect 69121 11713 69155 11747
rect 69213 11713 69247 11747
rect 88257 11713 88291 11747
rect 21189 11645 21223 11679
rect 24961 11645 24995 11679
rect 26985 11645 27019 11679
rect 27261 11645 27295 11679
rect 28365 11645 28399 11679
rect 29837 11645 29871 11679
rect 33333 11645 33367 11679
rect 36277 11645 36311 11679
rect 36645 11645 36679 11679
rect 37933 11645 37967 11679
rect 39313 11645 39347 11679
rect 39405 11645 39439 11679
rect 39589 11645 39623 11679
rect 44833 11645 44867 11679
rect 54657 11645 54691 11679
rect 59645 11645 59679 11679
rect 60841 11645 60875 11679
rect 63601 11645 63635 11679
rect 68201 11645 68235 11679
rect 71697 11645 71731 11679
rect 71789 11645 71823 11679
rect 1409 11577 1443 11611
rect 19349 11577 19383 11611
rect 25329 11577 25363 11611
rect 31677 11577 31711 11611
rect 35449 11577 35483 11611
rect 37289 11577 37323 11611
rect 58265 11577 58299 11611
rect 68937 11577 68971 11611
rect 88073 11577 88107 11611
rect 18613 11509 18647 11543
rect 21005 11509 21039 11543
rect 24409 11509 24443 11543
rect 29285 11509 29319 11543
rect 32597 11509 32631 11543
rect 34713 11509 34747 11543
rect 38163 11509 38197 11543
rect 39129 11509 39163 11543
rect 40417 11509 40451 11543
rect 41383 11509 41417 11543
rect 44465 11509 44499 11543
rect 46581 11509 46615 11543
rect 53573 11509 53607 11543
rect 55229 11509 55263 11543
rect 59185 11509 59219 11543
rect 62221 11509 62255 11543
rect 64429 11509 64463 11543
rect 68569 11509 68603 11543
rect 15577 11305 15611 11339
rect 24501 11305 24535 11339
rect 24869 11305 24903 11339
rect 27629 11305 27663 11339
rect 34253 11305 34287 11339
rect 35633 11305 35667 11339
rect 38761 11305 38795 11339
rect 39865 11305 39899 11339
rect 42349 11305 42383 11339
rect 45017 11305 45051 11339
rect 45661 11305 45695 11339
rect 53481 11305 53515 11339
rect 55413 11305 55447 11339
rect 55965 11305 55999 11339
rect 59737 11305 59771 11339
rect 60473 11305 60507 11339
rect 62313 11305 62347 11339
rect 25329 11237 25363 11271
rect 32137 11237 32171 11271
rect 41705 11237 41739 11271
rect 47593 11237 47627 11271
rect 49433 11237 49467 11271
rect 50813 11237 50847 11271
rect 52561 11237 52595 11271
rect 57989 11237 58023 11271
rect 61025 11237 61059 11271
rect 67281 11237 67315 11271
rect 69213 11237 69247 11271
rect 34713 11169 34747 11203
rect 36645 11169 36679 11203
rect 38210 11169 38244 11203
rect 39129 11169 39163 11203
rect 41061 11169 41095 11203
rect 41337 11169 41371 11203
rect 51181 11169 51215 11203
rect 56609 11169 56643 11203
rect 61577 11169 61611 11203
rect 63601 11169 63635 11203
rect 63785 11169 63819 11203
rect 67833 11169 67867 11203
rect 87705 11169 87739 11203
rect 46121 11135 46155 11169
rect 1593 11101 1627 11135
rect 15301 11101 15335 11135
rect 15393 11101 15427 11135
rect 24409 11101 24443 11135
rect 25237 11101 25271 11135
rect 25789 11101 25823 11135
rect 27813 11101 27847 11135
rect 29101 11101 29135 11135
rect 29561 11101 29595 11135
rect 31769 11101 31803 11135
rect 31953 11101 31987 11135
rect 32873 11101 32907 11135
rect 34897 11101 34931 11135
rect 35817 11101 35851 11135
rect 36001 11101 36035 11135
rect 36093 11101 36127 11135
rect 36921 11101 36955 11135
rect 37999 11101 38033 11135
rect 38117 11101 38151 11135
rect 38301 11101 38335 11135
rect 38945 11101 38979 11135
rect 39037 11101 39071 11135
rect 39221 11101 39255 11135
rect 40049 11101 40083 11135
rect 40325 11101 40359 11135
rect 40969 11101 41003 11135
rect 41705 11101 41739 11135
rect 41981 11101 42015 11135
rect 42533 11101 42567 11135
rect 44281 11101 44315 11135
rect 44373 11101 44407 11135
rect 44557 11101 44591 11135
rect 45201 11101 45235 11135
rect 45845 11101 45879 11135
rect 46029 11101 46063 11135
rect 46673 11101 46707 11135
rect 46857 11101 46891 11135
rect 46949 11101 46983 11135
rect 47409 11101 47443 11135
rect 49433 11101 49467 11135
rect 49709 11101 49743 11135
rect 50537 11101 50571 11135
rect 50629 11101 50663 11135
rect 52929 11101 52963 11135
rect 53113 11101 53147 11135
rect 53297 11101 53331 11135
rect 55321 11101 55355 11135
rect 56149 11101 56183 11135
rect 58357 11101 58391 11135
rect 60657 11101 60691 11135
rect 61393 11101 61427 11135
rect 61485 11101 61519 11135
rect 62313 11101 62347 11135
rect 62589 11101 62623 11135
rect 63877 11101 63911 11135
rect 64245 11101 64279 11135
rect 64429 11101 64463 11135
rect 64705 11101 64739 11135
rect 67281 11101 67315 11135
rect 67465 11101 67499 11135
rect 87429 11101 87463 11135
rect 26034 11033 26068 11067
rect 29806 11033 29840 11067
rect 33140 11033 33174 11067
rect 41889 11033 41923 11067
rect 46489 11033 46523 11067
rect 49617 11033 49651 11067
rect 51448 11033 51482 11067
rect 53205 11033 53239 11067
rect 56876 11033 56910 11067
rect 58602 11033 58636 11067
rect 63417 11033 63451 11067
rect 68078 11033 68112 11067
rect 1409 10965 1443 10999
rect 27169 10965 27203 10999
rect 28917 10965 28951 10999
rect 30941 10965 30975 10999
rect 35081 10965 35115 10999
rect 37841 10965 37875 10999
rect 40233 10965 40267 10999
rect 62497 10965 62531 10999
rect 64613 10965 64647 10999
rect 24777 10761 24811 10795
rect 26157 10761 26191 10795
rect 29101 10761 29135 10795
rect 33057 10761 33091 10795
rect 33701 10761 33735 10795
rect 35817 10761 35851 10795
rect 39037 10761 39071 10795
rect 40877 10761 40911 10795
rect 87705 10761 87739 10795
rect 50445 10693 50479 10727
rect 51917 10693 51951 10727
rect 56241 10693 56275 10727
rect 56793 10693 56827 10727
rect 58817 10693 58851 10727
rect 59829 10693 59863 10727
rect 61577 10693 61611 10727
rect 1593 10625 1627 10659
rect 28273 10625 28307 10659
rect 29009 10625 29043 10659
rect 30001 10625 30035 10659
rect 33241 10625 33275 10659
rect 33885 10625 33919 10659
rect 34253 10625 34287 10659
rect 35725 10625 35759 10659
rect 36461 10625 36495 10659
rect 36645 10625 36679 10659
rect 40049 10625 40083 10659
rect 40325 10625 40359 10659
rect 40785 10625 40819 10659
rect 42993 10625 43027 10659
rect 43361 10625 43395 10659
rect 45017 10625 45051 10659
rect 46009 10625 46043 10659
rect 47777 10625 47811 10659
rect 48697 10625 48731 10659
rect 50813 10625 50847 10659
rect 50997 10625 51031 10659
rect 51181 10625 51215 10659
rect 52929 10625 52963 10659
rect 53481 10625 53515 10659
rect 54657 10625 54691 10659
rect 56149 10625 56183 10659
rect 56701 10625 56735 10659
rect 57437 10625 57471 10659
rect 58633 10625 58667 10659
rect 58909 10625 58943 10659
rect 62313 10625 62347 10659
rect 63233 10625 63267 10659
rect 63417 10625 63451 10659
rect 63785 10625 63819 10659
rect 64041 10625 64075 10659
rect 65533 10625 65567 10659
rect 65789 10625 65823 10659
rect 88257 10625 88291 10659
rect 24869 10557 24903 10591
rect 25053 10557 25087 10591
rect 25697 10557 25731 10591
rect 29193 10557 29227 10591
rect 29745 10557 29779 10591
rect 36553 10557 36587 10591
rect 36737 10557 36771 10591
rect 37289 10557 37323 10591
rect 37565 10557 37599 10591
rect 38393 10557 38427 10591
rect 39129 10557 39163 10591
rect 39313 10557 39347 10591
rect 40233 10557 40267 10591
rect 42717 10557 42751 10591
rect 44005 10557 44039 10591
rect 45109 10557 45143 10591
rect 45385 10557 45419 10591
rect 45753 10557 45787 10591
rect 52009 10557 52043 10591
rect 52193 10557 52227 10591
rect 54401 10557 54435 10591
rect 63325 10557 63359 10591
rect 25973 10489 26007 10523
rect 28641 10489 28675 10523
rect 42901 10489 42935 10523
rect 44373 10489 44407 10523
rect 47593 10489 47627 10523
rect 52745 10489 52779 10523
rect 57253 10489 57287 10523
rect 62129 10489 62163 10523
rect 1409 10421 1443 10455
rect 24409 10421 24443 10455
rect 28089 10421 28123 10455
rect 31125 10421 31159 10455
rect 34345 10421 34379 10455
rect 36277 10421 36311 10455
rect 38669 10421 38703 10455
rect 39865 10421 39899 10455
rect 42533 10421 42567 10455
rect 43545 10421 43579 10455
rect 44465 10421 44499 10455
rect 47133 10421 47167 10455
rect 51549 10421 51583 10455
rect 53297 10421 53331 10455
rect 55781 10421 55815 10455
rect 58449 10421 58483 10455
rect 65165 10421 65199 10455
rect 66913 10421 66947 10455
rect 88073 10421 88107 10455
rect 25053 10217 25087 10251
rect 28917 10217 28951 10251
rect 33885 10217 33919 10251
rect 39865 10217 39899 10251
rect 40785 10217 40819 10251
rect 43637 10217 43671 10251
rect 47225 10217 47259 10251
rect 49617 10217 49651 10251
rect 51365 10217 51399 10251
rect 59461 10217 59495 10251
rect 61669 10217 61703 10251
rect 62221 10217 62255 10251
rect 64889 10217 64923 10251
rect 37749 10149 37783 10183
rect 46673 10149 46707 10183
rect 47409 10149 47443 10183
rect 49065 10149 49099 10183
rect 54125 10149 54159 10183
rect 39129 10081 39163 10115
rect 50629 10081 50663 10115
rect 50721 10081 50755 10115
rect 53757 10081 53791 10115
rect 54677 10081 54711 10115
rect 55321 10081 55355 10115
rect 58081 10081 58115 10115
rect 61025 10081 61059 10115
rect 64613 10081 64647 10115
rect 1593 10013 1627 10047
rect 25237 10013 25271 10047
rect 29101 10013 29135 10047
rect 29561 10013 29595 10047
rect 32505 10013 32539 10047
rect 34897 10013 34931 10047
rect 36001 10013 36035 10047
rect 40049 10013 40083 10047
rect 40233 10013 40267 10047
rect 40325 10013 40359 10047
rect 40693 10013 40727 10047
rect 42257 10013 42291 10047
rect 45293 10013 45327 10047
rect 48973 10013 49007 10047
rect 49525 10013 49559 10047
rect 51273 10013 51307 10047
rect 52009 10013 52043 10047
rect 57805 10013 57839 10047
rect 57897 10013 57931 10047
rect 59093 10013 59127 10047
rect 59277 10013 59311 10047
rect 60013 10013 60047 10047
rect 60841 10013 60875 10047
rect 61577 10013 61611 10047
rect 62129 10013 62163 10047
rect 64521 10013 64555 10047
rect 29806 9945 29840 9979
rect 32772 9945 32806 9979
rect 36461 9945 36495 9979
rect 42524 9945 42558 9979
rect 45560 9945 45594 9979
rect 47041 9945 47075 9979
rect 54493 9945 54527 9979
rect 55566 9945 55600 9979
rect 1409 9877 1443 9911
rect 30941 9877 30975 9911
rect 34713 9877 34747 9911
rect 35817 9877 35851 9911
rect 38577 9877 38611 9911
rect 38945 9877 38979 9911
rect 39037 9877 39071 9911
rect 47241 9877 47275 9911
rect 50169 9877 50203 9911
rect 50537 9877 50571 9911
rect 54585 9877 54619 9911
rect 56701 9877 56735 9911
rect 57437 9877 57471 9911
rect 58817 9877 58851 9911
rect 59829 9877 59863 9911
rect 60473 9877 60507 9911
rect 60933 9877 60967 9911
rect 29745 9673 29779 9707
rect 36553 9673 36587 9707
rect 37657 9673 37691 9707
rect 50997 9673 51031 9707
rect 54125 9673 54159 9707
rect 54493 9673 54527 9707
rect 55413 9673 55447 9707
rect 60841 9673 60875 9707
rect 64455 9673 64489 9707
rect 68201 9673 68235 9707
rect 33517 9605 33551 9639
rect 35440 9605 35474 9639
rect 37289 9605 37323 9639
rect 45201 9605 45235 9639
rect 51457 9605 51491 9639
rect 59728 9605 59762 9639
rect 64245 9605 64279 9639
rect 30113 9537 30147 9571
rect 35173 9537 35207 9571
rect 37473 9537 37507 9571
rect 37749 9537 37783 9571
rect 38577 9537 38611 9571
rect 38844 9537 38878 9571
rect 40325 9537 40359 9571
rect 40581 9537 40615 9571
rect 42625 9537 42659 9571
rect 45109 9537 45143 9571
rect 46009 9537 46043 9571
rect 49249 9537 49283 9571
rect 49617 9537 49651 9571
rect 49873 9537 49907 9571
rect 51365 9537 51399 9571
rect 52745 9537 52779 9571
rect 53012 9537 53046 9571
rect 54677 9537 54711 9571
rect 57253 9537 57287 9571
rect 59461 9537 59495 9571
rect 68385 9537 68419 9571
rect 69029 9537 69063 9571
rect 30205 9469 30239 9503
rect 30297 9469 30331 9503
rect 33609 9469 33643 9503
rect 33793 9469 33827 9503
rect 42717 9469 42751 9503
rect 42993 9469 43027 9503
rect 45753 9469 45787 9503
rect 55505 9469 55539 9503
rect 55597 9469 55631 9503
rect 68753 9469 68787 9503
rect 33149 9401 33183 9435
rect 47133 9401 47167 9435
rect 49065 9401 49099 9435
rect 55045 9401 55079 9435
rect 57069 9401 57103 9435
rect 64613 9401 64647 9435
rect 39957 9333 39991 9367
rect 41705 9333 41739 9367
rect 64429 9333 64463 9367
rect 70133 9333 70167 9367
rect 36277 9129 36311 9163
rect 37381 9129 37415 9163
rect 38669 9129 38703 9163
rect 44097 9129 44131 9163
rect 45845 9129 45879 9163
rect 48145 9129 48179 9163
rect 51733 9129 51767 9163
rect 55321 9129 55355 9163
rect 68201 9129 68235 9163
rect 47777 9061 47811 9095
rect 36829 8993 36863 9027
rect 42717 8993 42751 9027
rect 48697 8993 48731 9027
rect 52745 8993 52779 9027
rect 68753 8993 68787 9027
rect 87705 8993 87739 9027
rect 1593 8925 1627 8959
rect 36645 8925 36679 8959
rect 37565 8925 37599 8959
rect 37749 8925 37783 8959
rect 37841 8925 37875 8959
rect 38853 8925 38887 8959
rect 42349 8925 42383 8959
rect 46029 8925 46063 8959
rect 46397 8925 46431 8959
rect 48513 8925 48547 8959
rect 50169 8925 50203 8959
rect 50445 8925 50479 8959
rect 52377 8925 52411 8959
rect 55505 8925 55539 8959
rect 68569 8925 68603 8959
rect 87429 8925 87463 8959
rect 42962 8857 42996 8891
rect 46642 8857 46676 8891
rect 48605 8857 48639 8891
rect 52990 8857 53024 8891
rect 1409 8789 1443 8823
rect 36737 8789 36771 8823
rect 42165 8789 42199 8823
rect 52193 8789 52227 8823
rect 54125 8789 54159 8823
rect 68661 8789 68695 8823
rect 38025 8585 38059 8619
rect 42809 8585 42843 8619
rect 43177 8585 43211 8619
rect 46121 8585 46155 8619
rect 46489 8585 46523 8619
rect 49525 8585 49559 8619
rect 50261 8585 50295 8619
rect 52745 8585 52779 8619
rect 53113 8585 53147 8619
rect 43269 8517 43303 8551
rect 1685 8449 1719 8483
rect 38209 8449 38243 8483
rect 41613 8449 41647 8483
rect 50445 8449 50479 8483
rect 53205 8449 53239 8483
rect 88257 8449 88291 8483
rect 1409 8381 1443 8415
rect 41429 8381 41463 8415
rect 43361 8381 43395 8415
rect 46581 8381 46615 8415
rect 46673 8381 46707 8415
rect 49617 8381 49651 8415
rect 49709 8381 49743 8415
rect 53297 8381 53331 8415
rect 49157 8313 49191 8347
rect 88073 8313 88107 8347
rect 41797 8245 41831 8279
rect 46489 8041 46523 8075
rect 41889 7837 41923 7871
rect 46673 7837 46707 7871
rect 87705 7837 87739 7871
rect 88257 7837 88291 7871
rect 41705 7701 41739 7735
rect 88073 7701 88107 7735
rect 40325 7497 40359 7531
rect 39037 7429 39071 7463
rect 1593 7361 1627 7395
rect 88073 7361 88107 7395
rect 88257 7225 88291 7259
rect 1409 7157 1443 7191
rect 26157 6749 26191 6783
rect 26433 6749 26467 6783
rect 39037 6749 39071 6783
rect 39313 6749 39347 6783
rect 56793 6749 56827 6783
rect 38853 6681 38887 6715
rect 25973 6613 26007 6647
rect 26341 6613 26375 6647
rect 39221 6613 39255 6647
rect 56609 6613 56643 6647
rect 57161 6409 57195 6443
rect 1777 6273 1811 6307
rect 55781 6273 55815 6307
rect 56057 6273 56091 6307
rect 87429 6205 87463 6239
rect 87705 6205 87739 6239
rect 2053 6069 2087 6103
rect 56977 5865 57011 5899
rect 56701 5729 56735 5763
rect 57621 5729 57655 5763
rect 1593 5661 1627 5695
rect 3065 5661 3099 5695
rect 25145 5661 25179 5695
rect 25697 5661 25731 5695
rect 57345 5661 57379 5695
rect 57437 5661 57471 5695
rect 87981 5661 88015 5695
rect 25942 5593 25976 5627
rect 1409 5525 1443 5559
rect 2881 5525 2915 5559
rect 24961 5525 24995 5559
rect 27077 5525 27111 5559
rect 88165 5525 88199 5559
rect 24225 5321 24259 5355
rect 27721 5321 27755 5355
rect 30021 5321 30055 5355
rect 24593 5253 24627 5287
rect 29929 5253 29963 5287
rect 27169 5185 27203 5219
rect 87705 5185 87739 5219
rect 88257 5185 88291 5219
rect 24685 5117 24719 5151
rect 24777 5117 24811 5151
rect 26985 5117 27019 5151
rect 27353 4981 27387 5015
rect 88073 4981 88107 5015
rect 33057 4777 33091 4811
rect 24409 4709 24443 4743
rect 25513 4709 25547 4743
rect 87705 4709 87739 4743
rect 24961 4641 24995 4675
rect 26433 4641 26467 4675
rect 55321 4641 55355 4675
rect 56057 4641 56091 4675
rect 1593 4573 1627 4607
rect 25697 4573 25731 4607
rect 26157 4573 26191 4607
rect 55505 4573 55539 4607
rect 88257 4573 88291 4607
rect 24869 4505 24903 4539
rect 32781 4505 32815 4539
rect 33609 4505 33643 4539
rect 1409 4437 1443 4471
rect 24777 4437 24811 4471
rect 27537 4437 27571 4471
rect 33701 4437 33735 4471
rect 55689 4437 55723 4471
rect 88073 4437 88107 4471
rect 49433 4233 49467 4267
rect 51641 4165 51675 4199
rect 59553 4165 59587 4199
rect 70869 4165 70903 4199
rect 1685 4097 1719 4131
rect 2145 4097 2179 4131
rect 49617 4097 49651 4131
rect 51733 4097 51767 4131
rect 71329 4097 71363 4131
rect 87153 4097 87187 4131
rect 87705 4097 87739 4131
rect 88257 4097 88291 4131
rect 51825 4029 51859 4063
rect 71145 4029 71179 4063
rect 1961 3961 1995 3995
rect 87521 3961 87555 3995
rect 2421 3893 2455 3927
rect 51273 3893 51307 3927
rect 59645 3893 59679 3927
rect 71513 3893 71547 3927
rect 86601 3893 86635 3927
rect 86969 3893 87003 3927
rect 88073 3893 88107 3927
rect 27445 3689 27479 3723
rect 30849 3689 30883 3723
rect 49065 3689 49099 3723
rect 2513 3621 2547 3655
rect 86417 3621 86451 3655
rect 88349 3621 88383 3655
rect 33977 3553 34011 3587
rect 47777 3553 47811 3587
rect 51549 3553 51583 3587
rect 1593 3485 1627 3519
rect 2145 3485 2179 3519
rect 2697 3485 2731 3519
rect 24409 3485 24443 3519
rect 24593 3485 24627 3519
rect 26065 3485 26099 3519
rect 26709 3485 26743 3519
rect 27169 3485 27203 3519
rect 27261 3485 27295 3519
rect 28457 3485 28491 3519
rect 31217 3485 31251 3519
rect 31401 3485 31435 3519
rect 33057 3485 33091 3519
rect 49249 3485 49283 3519
rect 50353 3485 50387 3519
rect 50537 3485 50571 3519
rect 86601 3485 86635 3519
rect 86877 3485 86911 3519
rect 88073 3485 88107 3519
rect 88533 3485 88567 3519
rect 33793 3417 33827 3451
rect 50721 3417 50755 3451
rect 51794 3417 51828 3451
rect 87337 3417 87371 3451
rect 1409 3349 1443 3383
rect 1961 3349 1995 3383
rect 24777 3349 24811 3383
rect 25881 3349 25915 3383
rect 26525 3349 26559 3383
rect 28273 3349 28307 3383
rect 31585 3349 31619 3383
rect 32873 3349 32907 3383
rect 33425 3349 33459 3383
rect 33885 3349 33919 3383
rect 47133 3349 47167 3383
rect 47501 3349 47535 3383
rect 47593 3349 47627 3383
rect 52929 3349 52963 3383
rect 87705 3349 87739 3383
rect 1593 3145 1627 3179
rect 3525 3145 3559 3179
rect 46949 3145 46983 3179
rect 50997 3145 51031 3179
rect 52009 3145 52043 3179
rect 71421 3145 71455 3179
rect 85957 3145 85991 3179
rect 86785 3145 86819 3179
rect 88165 3145 88199 3179
rect 88349 3145 88383 3179
rect 33977 3077 34011 3111
rect 39681 3077 39715 3111
rect 49862 3077 49896 3111
rect 61945 3077 61979 3111
rect 76757 3077 76791 3111
rect 77125 3077 77159 3111
rect 1409 3009 1443 3043
rect 2237 3009 2271 3043
rect 3157 3009 3191 3043
rect 3709 3009 3743 3043
rect 4813 3009 4847 3043
rect 4997 3009 5031 3043
rect 5181 3009 5215 3043
rect 5733 3009 5767 3043
rect 6745 3009 6779 3043
rect 7113 3009 7147 3043
rect 9413 3009 9447 3043
rect 9965 3009 9999 3043
rect 12173 3009 12207 3043
rect 13829 3009 13863 3043
rect 17049 3009 17083 3043
rect 17693 3009 17727 3043
rect 19441 3009 19475 3043
rect 19809 3009 19843 3043
rect 20269 3009 20303 3043
rect 23029 3009 23063 3043
rect 25421 3009 25455 3043
rect 25973 3009 26007 3043
rect 26341 3009 26375 3043
rect 27445 3009 27479 3043
rect 27813 3009 27847 3043
rect 28069 3009 28103 3043
rect 29837 3009 29871 3043
rect 30021 3009 30055 3043
rect 30573 3009 30607 3043
rect 31677 3009 31711 3043
rect 32321 3009 32355 3043
rect 32597 3009 32631 3043
rect 34345 3009 34379 3043
rect 34805 3009 34839 3043
rect 38669 3009 38703 3043
rect 39037 3009 39071 3043
rect 39313 3009 39347 3043
rect 39497 3009 39531 3043
rect 40233 3009 40267 3043
rect 41981 3009 42015 3043
rect 42625 3009 42659 3043
rect 47133 3009 47167 3043
rect 47593 3009 47627 3043
rect 47869 3009 47903 3043
rect 49617 3009 49651 3043
rect 51641 3009 51675 3043
rect 52193 3009 52227 3043
rect 53021 3009 53055 3043
rect 53481 3009 53515 3043
rect 53757 3009 53791 3043
rect 54125 3009 54159 3043
rect 55873 3009 55907 3043
rect 58081 3009 58115 3043
rect 58633 3009 58667 3043
rect 61577 3009 61611 3043
rect 61761 3009 61795 3043
rect 63233 3009 63267 3043
rect 63509 3009 63543 3043
rect 63877 3009 63911 3043
rect 64797 3009 64831 3043
rect 68753 3009 68787 3043
rect 71605 3009 71639 3043
rect 72157 3009 72191 3043
rect 77677 3009 77711 3043
rect 77861 3009 77895 3043
rect 78689 3009 78723 3043
rect 81541 3009 81575 3043
rect 82093 3009 82127 3043
rect 86141 3009 86175 3043
rect 86969 3009 87003 3043
rect 87521 3009 87555 3043
rect 88073 3009 88107 3043
rect 88533 3009 88567 3043
rect 26433 2941 26467 2975
rect 29653 2941 29687 2975
rect 64521 2941 64555 2975
rect 77493 2941 77527 2975
rect 9229 2873 9263 2907
rect 19257 2873 19291 2907
rect 27261 2873 27295 2907
rect 29193 2873 29227 2907
rect 34621 2873 34655 2907
rect 41797 2873 41831 2907
rect 51457 2873 51491 2907
rect 53297 2873 53331 2907
rect 63693 2873 63727 2907
rect 2053 2805 2087 2839
rect 2973 2805 3007 2839
rect 5549 2805 5583 2839
rect 6561 2805 6595 2839
rect 9781 2805 9815 2839
rect 11989 2805 12023 2839
rect 13645 2805 13679 2839
rect 16865 2805 16899 2839
rect 17509 2805 17543 2839
rect 20085 2805 20119 2839
rect 22845 2805 22879 2839
rect 25237 2805 25271 2839
rect 25789 2805 25823 2839
rect 30389 2805 30423 2839
rect 31493 2805 31527 2839
rect 38485 2805 38519 2839
rect 40049 2805 40083 2839
rect 42441 2805 42475 2839
rect 49157 2805 49191 2839
rect 53573 2805 53607 2839
rect 53941 2805 53975 2839
rect 55689 2805 55723 2839
rect 57897 2805 57931 2839
rect 58449 2805 58483 2839
rect 63049 2805 63083 2839
rect 68569 2805 68603 2839
rect 71973 2805 72007 2839
rect 78505 2805 78539 2839
rect 81909 2805 81943 2839
rect 87337 2805 87371 2839
rect 11713 2601 11747 2635
rect 27905 2601 27939 2635
rect 48697 2601 48731 2635
rect 50169 2601 50203 2635
rect 51917 2601 51951 2635
rect 55321 2601 55355 2635
rect 55873 2601 55907 2635
rect 60473 2601 60507 2635
rect 61301 2601 61335 2635
rect 69029 2601 69063 2635
rect 70777 2601 70811 2635
rect 71329 2601 71363 2635
rect 4721 2533 4755 2567
rect 24041 2533 24075 2567
rect 25237 2533 25271 2567
rect 27353 2533 27387 2567
rect 44373 2533 44407 2567
rect 45201 2533 45235 2567
rect 79057 2533 79091 2567
rect 79977 2533 80011 2567
rect 80805 2533 80839 2567
rect 81725 2533 81759 2567
rect 86877 2533 86911 2567
rect 6653 2465 6687 2499
rect 13093 2465 13127 2499
rect 19257 2465 19291 2499
rect 28549 2465 28583 2499
rect 40141 2465 40175 2499
rect 50721 2465 50755 2499
rect 75101 2465 75135 2499
rect 2329 2397 2363 2431
rect 2789 2397 2823 2431
rect 3341 2397 3375 2431
rect 4905 2397 4939 2431
rect 5457 2397 5491 2431
rect 6377 2397 6411 2431
rect 7941 2397 7975 2431
rect 8493 2397 8527 2431
rect 9321 2397 9355 2431
rect 9965 2397 9999 2431
rect 10517 2397 10551 2431
rect 11069 2397 11103 2431
rect 12173 2397 12207 2431
rect 12817 2397 12851 2431
rect 14105 2397 14139 2431
rect 14381 2397 14415 2431
rect 15301 2397 15335 2431
rect 15761 2397 15795 2431
rect 16681 2397 16715 2431
rect 16957 2397 16991 2431
rect 18245 2397 18279 2431
rect 18797 2397 18831 2431
rect 19533 2397 19567 2431
rect 20821 2397 20855 2431
rect 21373 2397 21407 2431
rect 22017 2397 22051 2431
rect 23489 2397 23523 2431
rect 23949 2397 23983 2431
rect 24225 2397 24259 2431
rect 24777 2397 24811 2431
rect 25421 2397 25455 2431
rect 26065 2397 26099 2431
rect 26525 2397 26559 2431
rect 26801 2397 26835 2431
rect 27537 2397 27571 2431
rect 29929 2397 29963 2431
rect 30481 2397 30515 2431
rect 31669 2397 31703 2431
rect 32965 2397 32999 2431
rect 33241 2397 33275 2431
rect 34897 2397 34931 2431
rect 35725 2397 35759 2431
rect 36277 2397 36311 2431
rect 36829 2397 36863 2431
rect 37657 2397 37691 2431
rect 38945 2373 38979 2407
rect 39865 2397 39899 2431
rect 41245 2397 41279 2431
rect 41981 2397 42015 2431
rect 42809 2397 42843 2431
rect 43453 2397 43487 2431
rect 44005 2397 44039 2431
rect 44557 2397 44591 2431
rect 45385 2397 45419 2431
rect 46305 2397 46339 2431
rect 46581 2397 46615 2431
rect 47777 2397 47811 2431
rect 48329 2397 48363 2431
rect 48881 2397 48915 2431
rect 49525 2397 49559 2431
rect 52101 2397 52135 2431
rect 54401 2397 54435 2431
rect 55505 2397 55539 2431
rect 56057 2397 56091 2431
rect 56609 2397 56643 2431
rect 57161 2397 57195 2431
rect 58081 2397 58115 2431
rect 58633 2397 58667 2431
rect 59185 2397 59219 2431
rect 59737 2397 59771 2431
rect 60657 2397 60691 2431
rect 61485 2397 61519 2431
rect 62129 2397 62163 2431
rect 63233 2397 63267 2431
rect 63509 2397 63543 2431
rect 65809 2397 65843 2431
rect 66361 2397 66395 2431
rect 66913 2397 66947 2431
rect 67465 2397 67499 2431
rect 68385 2397 68419 2431
rect 69213 2397 69247 2431
rect 69857 2397 69891 2431
rect 70961 2397 70995 2431
rect 71513 2397 71547 2431
rect 72249 2397 72283 2431
rect 73537 2397 73571 2431
rect 74365 2397 74399 2431
rect 76113 2397 76147 2431
rect 76757 2397 76791 2431
rect 77585 2397 77619 2431
rect 78689 2397 78723 2431
rect 79241 2397 79275 2431
rect 79517 2397 79551 2431
rect 79793 2397 79827 2431
rect 80161 2397 80195 2431
rect 80437 2397 80471 2431
rect 80621 2397 80655 2431
rect 81909 2397 81943 2431
rect 83841 2397 83875 2431
rect 84669 2397 84703 2431
rect 85129 2397 85163 2431
rect 86417 2397 86451 2431
rect 86693 2397 86727 2431
rect 87061 2397 87095 2431
rect 1593 2329 1627 2363
rect 1961 2329 1995 2363
rect 4169 2329 4203 2363
rect 11621 2329 11655 2363
rect 28365 2329 28399 2363
rect 32413 2329 32447 2363
rect 51365 2329 51399 2363
rect 53113 2329 53147 2363
rect 74917 2329 74951 2363
rect 82645 2329 82679 2363
rect 87889 2329 87923 2363
rect 2605 2261 2639 2295
rect 3157 2261 3191 2295
rect 4261 2261 4295 2295
rect 5273 2261 5307 2295
rect 7757 2261 7791 2295
rect 8309 2261 8343 2295
rect 9137 2261 9171 2295
rect 9781 2261 9815 2295
rect 10333 2261 10367 2295
rect 10885 2261 10919 2295
rect 12357 2261 12391 2295
rect 15577 2261 15611 2295
rect 18613 2261 18647 2295
rect 20637 2261 20671 2295
rect 21189 2261 21223 2295
rect 22201 2261 22235 2295
rect 23765 2261 23799 2295
rect 24593 2261 24627 2295
rect 26341 2261 26375 2295
rect 26617 2261 26651 2295
rect 28273 2261 28307 2295
rect 29745 2261 29779 2295
rect 30297 2261 30331 2295
rect 31493 2261 31527 2295
rect 32505 2261 32539 2295
rect 34713 2261 34747 2295
rect 36093 2261 36127 2295
rect 36645 2261 36679 2295
rect 37473 2261 37507 2295
rect 38761 2261 38795 2295
rect 41061 2261 41095 2295
rect 41797 2261 41831 2295
rect 42625 2261 42659 2295
rect 43269 2261 43303 2295
rect 43821 2261 43855 2295
rect 48145 2261 48179 2295
rect 49617 2261 49651 2295
rect 50537 2261 50571 2295
rect 50629 2261 50663 2295
rect 51457 2261 51491 2295
rect 53205 2261 53239 2295
rect 54217 2261 54251 2295
rect 56425 2261 56459 2295
rect 56977 2261 57011 2295
rect 57897 2261 57931 2295
rect 58449 2261 58483 2295
rect 59001 2261 59035 2295
rect 61945 2261 61979 2295
rect 65625 2261 65659 2295
rect 66177 2261 66211 2295
rect 66729 2261 66763 2295
rect 67281 2261 67315 2295
rect 68201 2261 68235 2295
rect 69673 2261 69707 2295
rect 72433 2261 72467 2295
rect 73353 2261 73387 2295
rect 75929 2261 75963 2295
rect 76573 2261 76607 2295
rect 77033 2261 77067 2295
rect 77401 2261 77435 2295
rect 79333 2261 79367 2295
rect 80253 2261 80287 2295
rect 81449 2261 81483 2295
rect 82737 2261 82771 2295
rect 83657 2261 83691 2295
rect 84209 2261 84243 2295
rect 84485 2261 84519 2295
rect 85313 2261 85347 2295
rect 86233 2261 86267 2295
rect 87981 2261 88015 2295
<< metal1 >>
rect 1104 27770 88872 27792
rect 1104 27718 11924 27770
rect 11976 27718 11988 27770
rect 12040 27718 12052 27770
rect 12104 27718 12116 27770
rect 12168 27718 12180 27770
rect 12232 27718 33872 27770
rect 33924 27718 33936 27770
rect 33988 27718 34000 27770
rect 34052 27718 34064 27770
rect 34116 27718 34128 27770
rect 34180 27718 55820 27770
rect 55872 27718 55884 27770
rect 55936 27718 55948 27770
rect 56000 27718 56012 27770
rect 56064 27718 56076 27770
rect 56128 27718 77768 27770
rect 77820 27718 77832 27770
rect 77884 27718 77896 27770
rect 77948 27718 77960 27770
rect 78012 27718 78024 27770
rect 78076 27718 88872 27770
rect 1104 27696 88872 27718
rect 25866 27616 25872 27668
rect 25924 27656 25930 27668
rect 31294 27656 31300 27668
rect 25924 27628 27936 27656
rect 25924 27616 25930 27628
rect 2682 27588 2688 27600
rect 2643 27560 2688 27588
rect 2682 27548 2688 27560
rect 2740 27548 2746 27600
rect 5258 27588 5264 27600
rect 5219 27560 5264 27588
rect 5258 27548 5264 27560
rect 5316 27548 5322 27600
rect 7742 27588 7748 27600
rect 7703 27560 7748 27588
rect 7742 27548 7748 27560
rect 7800 27548 7806 27600
rect 8478 27588 8484 27600
rect 8439 27560 8484 27588
rect 8478 27548 8484 27560
rect 8536 27548 8542 27600
rect 9122 27588 9128 27600
rect 9083 27560 9128 27588
rect 9122 27548 9128 27560
rect 9180 27548 9186 27600
rect 9214 27548 9220 27600
rect 9272 27588 9278 27600
rect 12158 27588 12164 27600
rect 9272 27560 12164 27588
rect 9272 27548 9278 27560
rect 12158 27548 12164 27560
rect 12216 27548 12222 27600
rect 14274 27588 14280 27600
rect 14235 27560 14280 27588
rect 14274 27548 14280 27560
rect 14332 27548 14338 27600
rect 14918 27588 14924 27600
rect 14879 27560 14924 27588
rect 14918 27548 14924 27560
rect 14976 27548 14982 27600
rect 15562 27588 15568 27600
rect 15523 27560 15568 27588
rect 15562 27548 15568 27560
rect 15620 27548 15626 27600
rect 18046 27588 18052 27600
rect 18007 27560 18052 27588
rect 18046 27548 18052 27560
rect 18104 27548 18110 27600
rect 18598 27588 18604 27600
rect 18559 27560 18604 27588
rect 18598 27548 18604 27560
rect 18656 27548 18662 27600
rect 19978 27548 19984 27600
rect 20036 27588 20042 27600
rect 20073 27591 20131 27597
rect 20073 27588 20085 27591
rect 20036 27560 20085 27588
rect 20036 27548 20042 27560
rect 20073 27557 20085 27560
rect 20119 27557 20131 27591
rect 20622 27588 20628 27600
rect 20583 27560 20628 27588
rect 20073 27551 20131 27557
rect 20622 27548 20628 27560
rect 20680 27548 20686 27600
rect 22002 27588 22008 27600
rect 21963 27560 22008 27588
rect 22002 27548 22008 27560
rect 22060 27548 22066 27600
rect 22554 27588 22560 27600
rect 22515 27560 22560 27588
rect 22554 27548 22560 27560
rect 22612 27548 22618 27600
rect 24578 27588 24584 27600
rect 22940 27560 23244 27588
rect 24539 27560 24584 27588
rect 5810 27480 5816 27532
rect 5868 27520 5874 27532
rect 6365 27523 6423 27529
rect 6365 27520 6377 27523
rect 5868 27492 6377 27520
rect 5868 27480 5874 27492
rect 6365 27489 6377 27492
rect 6411 27489 6423 27523
rect 11606 27520 11612 27532
rect 6365 27483 6423 27489
rect 6472 27492 11468 27520
rect 11567 27492 11612 27520
rect 1302 27412 1308 27464
rect 1360 27452 1366 27464
rect 1397 27455 1455 27461
rect 1397 27452 1409 27455
rect 1360 27424 1409 27452
rect 1360 27412 1366 27424
rect 1397 27421 1409 27424
rect 1443 27421 1455 27455
rect 2222 27452 2228 27464
rect 2183 27424 2228 27452
rect 1397 27415 1455 27421
rect 2222 27412 2228 27424
rect 2280 27412 2286 27464
rect 2869 27455 2927 27461
rect 2869 27421 2881 27455
rect 2915 27452 2927 27455
rect 3142 27452 3148 27464
rect 2915 27424 3148 27452
rect 2915 27421 2927 27424
rect 2869 27415 2927 27421
rect 3142 27412 3148 27424
rect 3200 27412 3206 27464
rect 3234 27412 3240 27464
rect 3292 27452 3298 27464
rect 3789 27455 3847 27461
rect 3789 27452 3801 27455
rect 3292 27424 3801 27452
rect 3292 27412 3298 27424
rect 3789 27421 3801 27424
rect 3835 27421 3847 27455
rect 4706 27452 4712 27464
rect 4667 27424 4712 27452
rect 3789 27415 3847 27421
rect 4706 27412 4712 27424
rect 4764 27412 4770 27464
rect 5445 27455 5503 27461
rect 5445 27421 5457 27455
rect 5491 27452 5503 27455
rect 6472 27452 6500 27492
rect 6638 27452 6644 27464
rect 5491 27424 6500 27452
rect 6599 27424 6644 27452
rect 5491 27421 5503 27424
rect 5445 27415 5503 27421
rect 6638 27412 6644 27424
rect 6696 27412 6702 27464
rect 7929 27455 7987 27461
rect 7929 27421 7941 27455
rect 7975 27452 7987 27455
rect 9214 27452 9220 27464
rect 7975 27424 9220 27452
rect 7975 27421 7987 27424
rect 7929 27415 7987 27421
rect 9214 27412 9220 27424
rect 9272 27412 9278 27464
rect 9309 27455 9367 27461
rect 9309 27421 9321 27455
rect 9355 27452 9367 27455
rect 9674 27452 9680 27464
rect 9355 27424 9680 27452
rect 9355 27421 9367 27424
rect 9309 27415 9367 27421
rect 9674 27412 9680 27424
rect 9732 27412 9738 27464
rect 10229 27455 10287 27461
rect 10229 27421 10241 27455
rect 10275 27421 10287 27455
rect 10502 27452 10508 27464
rect 10463 27424 10508 27452
rect 10229 27415 10287 27421
rect 10244 27384 10272 27415
rect 10502 27412 10508 27424
rect 10560 27412 10566 27464
rect 11440 27452 11468 27492
rect 11606 27480 11612 27492
rect 11664 27480 11670 27532
rect 22940 27520 22968 27560
rect 23106 27520 23112 27532
rect 11716 27492 22968 27520
rect 23067 27492 23112 27520
rect 11716 27452 11744 27492
rect 23106 27480 23112 27492
rect 23164 27480 23170 27532
rect 23216 27520 23244 27560
rect 24578 27548 24584 27560
rect 24636 27548 24642 27600
rect 25317 27591 25375 27597
rect 25317 27557 25329 27591
rect 25363 27588 25375 27591
rect 26418 27588 26424 27600
rect 25363 27560 26424 27588
rect 25363 27557 25375 27560
rect 25317 27551 25375 27557
rect 26418 27548 26424 27560
rect 26476 27548 26482 27600
rect 27154 27588 27160 27600
rect 27115 27560 27160 27588
rect 27154 27548 27160 27560
rect 27212 27548 27218 27600
rect 27798 27588 27804 27600
rect 27759 27560 27804 27588
rect 27798 27548 27804 27560
rect 27856 27548 27862 27600
rect 27908 27588 27936 27628
rect 28966 27628 31300 27656
rect 28966 27588 28994 27628
rect 31294 27616 31300 27628
rect 31352 27616 31358 27668
rect 36538 27616 36544 27668
rect 36596 27656 36602 27668
rect 36633 27659 36691 27665
rect 36633 27656 36645 27659
rect 36596 27628 36645 27656
rect 36596 27616 36602 27628
rect 36633 27625 36645 27628
rect 36679 27625 36691 27659
rect 52270 27656 52276 27668
rect 36633 27619 36691 27625
rect 37936 27628 39988 27656
rect 29730 27588 29736 27600
rect 27908 27560 28994 27588
rect 29691 27560 29736 27588
rect 29730 27548 29736 27560
rect 29788 27548 29794 27600
rect 33502 27588 33508 27600
rect 33463 27560 33508 27588
rect 33502 27548 33508 27560
rect 33560 27548 33566 27600
rect 34057 27591 34115 27597
rect 34057 27557 34069 27591
rect 34103 27588 34115 27591
rect 34238 27588 34244 27600
rect 34103 27560 34244 27588
rect 34103 27557 34115 27560
rect 34057 27551 34115 27557
rect 34238 27548 34244 27560
rect 34296 27548 34302 27600
rect 34882 27588 34888 27600
rect 34843 27560 34888 27588
rect 34882 27548 34888 27560
rect 34940 27548 34946 27600
rect 35526 27588 35532 27600
rect 35487 27560 35532 27588
rect 35526 27548 35532 27560
rect 35584 27548 35590 27600
rect 36078 27588 36084 27600
rect 36039 27560 36084 27588
rect 36078 27548 36084 27560
rect 36136 27548 36142 27600
rect 36170 27548 36176 27600
rect 36228 27588 36234 27600
rect 37274 27588 37280 27600
rect 36228 27560 37280 27588
rect 36228 27548 36234 27560
rect 37274 27548 37280 27560
rect 37332 27548 37338 27600
rect 37458 27588 37464 27600
rect 37419 27560 37464 27588
rect 37458 27548 37464 27560
rect 37516 27548 37522 27600
rect 37550 27548 37556 27600
rect 37608 27588 37614 27600
rect 37936 27588 37964 27628
rect 38102 27588 38108 27600
rect 37608 27560 37964 27588
rect 38063 27560 38108 27588
rect 37608 27548 37614 27560
rect 38102 27548 38108 27560
rect 38160 27548 38166 27600
rect 38746 27588 38752 27600
rect 38707 27560 38752 27588
rect 38746 27548 38752 27560
rect 38804 27548 38810 27600
rect 39298 27548 39304 27600
rect 39356 27588 39362 27600
rect 39853 27591 39911 27597
rect 39853 27588 39865 27591
rect 39356 27560 39865 27588
rect 39356 27548 39362 27560
rect 39853 27557 39865 27560
rect 39899 27557 39911 27591
rect 39960 27588 39988 27628
rect 40512 27628 41552 27656
rect 40512 27588 40540 27628
rect 40678 27588 40684 27600
rect 39960 27560 40540 27588
rect 40639 27560 40684 27588
rect 39853 27551 39911 27557
rect 40678 27548 40684 27560
rect 40736 27548 40742 27600
rect 41524 27588 41552 27628
rect 42444 27628 43944 27656
rect 42444 27588 42472 27628
rect 42610 27588 42616 27600
rect 41248 27560 41414 27588
rect 41524 27560 42472 27588
rect 42571 27560 42616 27588
rect 29362 27520 29368 27532
rect 23216 27492 29368 27520
rect 29362 27480 29368 27492
rect 29420 27480 29426 27532
rect 30834 27520 30840 27532
rect 30795 27492 30840 27520
rect 30834 27480 30840 27492
rect 30892 27480 30898 27532
rect 31570 27480 31576 27532
rect 31628 27520 31634 27532
rect 32401 27523 32459 27529
rect 32401 27520 32413 27523
rect 31628 27492 32413 27520
rect 31628 27480 31634 27492
rect 32401 27489 32413 27492
rect 32447 27489 32459 27523
rect 32401 27483 32459 27489
rect 32674 27480 32680 27532
rect 32732 27520 32738 27532
rect 41248 27520 41276 27560
rect 32732 27492 39896 27520
rect 32732 27480 32738 27492
rect 39868 27464 39896 27492
rect 40052 27492 41276 27520
rect 41386 27520 41414 27560
rect 42610 27548 42616 27560
rect 42668 27548 42674 27600
rect 43254 27588 43260 27600
rect 43215 27560 43260 27588
rect 43254 27548 43260 27560
rect 43312 27548 43318 27600
rect 43806 27588 43812 27600
rect 43767 27560 43812 27588
rect 43806 27548 43812 27560
rect 43864 27548 43870 27600
rect 43916 27588 43944 27628
rect 45020 27628 46612 27656
rect 45020 27588 45048 27628
rect 45186 27588 45192 27600
rect 43916 27560 45048 27588
rect 45147 27560 45192 27588
rect 45186 27548 45192 27560
rect 45244 27548 45250 27600
rect 45830 27588 45836 27600
rect 45791 27560 45836 27588
rect 45830 27548 45836 27560
rect 45888 27548 45894 27600
rect 46474 27588 46480 27600
rect 46435 27560 46480 27588
rect 46474 27548 46480 27560
rect 46532 27548 46538 27600
rect 46584 27588 46612 27628
rect 48286 27628 52276 27656
rect 48286 27588 48314 27628
rect 52270 27616 52276 27628
rect 52328 27616 52334 27668
rect 52380 27628 52868 27656
rect 49050 27588 49056 27600
rect 46584 27560 48314 27588
rect 49011 27560 49056 27588
rect 49050 27548 49056 27560
rect 49108 27548 49114 27600
rect 51074 27548 51080 27600
rect 51132 27588 51138 27600
rect 51132 27560 51177 27588
rect 51132 27548 51138 27560
rect 51258 27548 51264 27600
rect 51316 27588 51322 27600
rect 52380 27588 52408 27628
rect 51316 27560 52408 27588
rect 51316 27548 51322 27560
rect 52454 27548 52460 27600
rect 52512 27588 52518 27600
rect 52733 27591 52791 27597
rect 52733 27588 52745 27591
rect 52512 27560 52745 27588
rect 52512 27548 52518 27560
rect 52733 27557 52745 27560
rect 52779 27557 52791 27591
rect 52840 27588 52868 27628
rect 55674 27588 55680 27600
rect 52840 27560 55680 27588
rect 52733 27551 52791 27557
rect 55674 27548 55680 27560
rect 55732 27548 55738 27600
rect 56137 27591 56195 27597
rect 56137 27557 56149 27591
rect 56183 27588 56195 27591
rect 56226 27588 56232 27600
rect 56183 27560 56232 27588
rect 56183 27557 56195 27560
rect 56137 27551 56195 27557
rect 56226 27548 56232 27560
rect 56284 27548 56290 27600
rect 56778 27588 56784 27600
rect 56739 27560 56784 27588
rect 56778 27548 56784 27560
rect 56836 27548 56842 27600
rect 57330 27548 57336 27600
rect 57388 27588 57394 27600
rect 57885 27591 57943 27597
rect 57885 27588 57897 27591
rect 57388 27560 57897 27588
rect 57388 27548 57394 27560
rect 57885 27557 57897 27560
rect 57931 27557 57943 27591
rect 59354 27588 59360 27600
rect 59315 27560 59360 27588
rect 57885 27551 57943 27557
rect 59354 27548 59360 27560
rect 59412 27548 59418 27600
rect 59906 27548 59912 27600
rect 59964 27588 59970 27600
rect 60461 27591 60519 27597
rect 60461 27588 60473 27591
rect 59964 27560 60473 27588
rect 59964 27548 59970 27560
rect 60461 27557 60473 27560
rect 60507 27557 60519 27591
rect 60461 27551 60519 27557
rect 60550 27548 60556 27600
rect 60608 27588 60614 27600
rect 61473 27591 61531 27597
rect 61473 27588 61485 27591
rect 60608 27560 61485 27588
rect 60608 27548 60614 27560
rect 61473 27557 61485 27560
rect 61519 27557 61531 27591
rect 61930 27588 61936 27600
rect 61891 27560 61936 27588
rect 61473 27551 61531 27557
rect 61930 27548 61936 27560
rect 61988 27548 61994 27600
rect 62482 27548 62488 27600
rect 62540 27588 62546 27600
rect 63037 27591 63095 27597
rect 63037 27588 63049 27591
rect 62540 27560 63049 27588
rect 62540 27548 62546 27560
rect 63037 27557 63049 27560
rect 63083 27557 63095 27591
rect 63037 27551 63095 27557
rect 65058 27548 65064 27600
rect 65116 27588 65122 27600
rect 65613 27591 65671 27597
rect 65613 27588 65625 27591
rect 65116 27560 65625 27588
rect 65116 27548 65122 27560
rect 65613 27557 65625 27560
rect 65659 27557 65671 27591
rect 65613 27551 65671 27557
rect 65702 27548 65708 27600
rect 65760 27588 65766 27600
rect 66165 27591 66223 27597
rect 66165 27588 66177 27591
rect 65760 27560 66177 27588
rect 65760 27548 65766 27560
rect 66165 27557 66177 27560
rect 66211 27557 66223 27591
rect 66165 27551 66223 27557
rect 66346 27548 66352 27600
rect 66404 27588 66410 27600
rect 66717 27591 66775 27597
rect 66717 27588 66729 27591
rect 66404 27560 66729 27588
rect 66404 27548 66410 27560
rect 66717 27557 66729 27560
rect 66763 27557 66775 27591
rect 66717 27551 66775 27557
rect 69014 27548 69020 27600
rect 69072 27588 69078 27600
rect 69661 27591 69719 27597
rect 69661 27588 69673 27591
rect 69072 27560 69673 27588
rect 69072 27548 69078 27560
rect 69661 27557 69673 27560
rect 69707 27557 69719 27591
rect 69661 27551 69719 27557
rect 70394 27548 70400 27600
rect 70452 27588 70458 27600
rect 71317 27591 71375 27597
rect 71317 27588 71329 27591
rect 70452 27560 71329 27588
rect 70452 27548 70458 27560
rect 71317 27557 71329 27560
rect 71363 27557 71375 27591
rect 71317 27551 71375 27557
rect 71498 27548 71504 27600
rect 71556 27588 71562 27600
rect 71869 27591 71927 27597
rect 71869 27588 71881 27591
rect 71556 27560 71881 27588
rect 71556 27548 71562 27560
rect 71869 27557 71881 27560
rect 71915 27557 71927 27591
rect 72418 27588 72424 27600
rect 72379 27560 72424 27588
rect 71869 27551 71927 27557
rect 72418 27548 72424 27560
rect 72476 27548 72482 27600
rect 74258 27588 74264 27600
rect 74219 27560 74264 27588
rect 74258 27548 74264 27560
rect 74316 27548 74322 27600
rect 74810 27588 74816 27600
rect 74771 27560 74816 27588
rect 74810 27548 74816 27560
rect 74868 27548 74874 27600
rect 76834 27588 76840 27600
rect 76795 27560 76840 27588
rect 76834 27548 76840 27560
rect 76892 27548 76898 27600
rect 77386 27588 77392 27600
rect 77347 27560 77392 27588
rect 77386 27548 77392 27560
rect 77444 27548 77450 27600
rect 81986 27588 81992 27600
rect 81947 27560 81992 27588
rect 81986 27548 81992 27560
rect 82044 27548 82050 27600
rect 83090 27548 83096 27600
rect 83148 27588 83154 27600
rect 83645 27591 83703 27597
rect 83645 27588 83657 27591
rect 83148 27560 83657 27588
rect 83148 27548 83154 27560
rect 83645 27557 83657 27560
rect 83691 27557 83703 27591
rect 83645 27551 83703 27557
rect 83734 27548 83740 27600
rect 83792 27588 83798 27600
rect 85301 27591 85359 27597
rect 85301 27588 85313 27591
rect 83792 27560 85313 27588
rect 83792 27548 83798 27560
rect 85301 27557 85313 27560
rect 85347 27557 85359 27591
rect 85301 27551 85359 27557
rect 85666 27548 85672 27600
rect 85724 27588 85730 27600
rect 86221 27591 86279 27597
rect 86221 27588 86233 27591
rect 85724 27560 86233 27588
rect 85724 27548 85730 27560
rect 86221 27557 86233 27560
rect 86267 27557 86279 27591
rect 89530 27588 89536 27600
rect 86221 27551 86279 27557
rect 86788 27560 89536 27588
rect 41386 27492 42104 27520
rect 11440 27424 11744 27452
rect 11885 27455 11943 27461
rect 11885 27421 11897 27455
rect 11931 27452 11943 27455
rect 12250 27452 12256 27464
rect 11931 27424 12256 27452
rect 11931 27421 11943 27424
rect 11885 27415 11943 27421
rect 12250 27412 12256 27424
rect 12308 27412 12314 27464
rect 12802 27452 12808 27464
rect 12763 27424 12808 27452
rect 12802 27412 12808 27424
rect 12860 27412 12866 27464
rect 13078 27452 13084 27464
rect 13039 27424 13084 27452
rect 13078 27412 13084 27424
rect 13136 27412 13142 27464
rect 14458 27452 14464 27464
rect 14419 27424 14464 27452
rect 14458 27412 14464 27424
rect 14516 27412 14522 27464
rect 15102 27452 15108 27464
rect 15063 27424 15108 27452
rect 15102 27412 15108 27424
rect 15160 27412 15166 27464
rect 15746 27452 15752 27464
rect 15707 27424 15752 27452
rect 15746 27412 15752 27424
rect 15804 27412 15810 27464
rect 16574 27412 16580 27464
rect 16632 27452 16638 27464
rect 16669 27455 16727 27461
rect 16669 27452 16681 27455
rect 16632 27424 16681 27452
rect 16632 27412 16638 27424
rect 16669 27421 16681 27424
rect 16715 27421 16727 27455
rect 16669 27415 16727 27421
rect 16945 27455 17003 27461
rect 16945 27421 16957 27455
rect 16991 27452 17003 27455
rect 18046 27452 18052 27464
rect 16991 27424 18052 27452
rect 16991 27421 17003 27424
rect 16945 27415 17003 27421
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 18230 27452 18236 27464
rect 18191 27424 18236 27452
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 18782 27452 18788 27464
rect 18743 27424 18788 27452
rect 18782 27412 18788 27424
rect 18840 27412 18846 27464
rect 19610 27452 19616 27464
rect 19571 27424 19616 27452
rect 19610 27412 19616 27424
rect 19668 27412 19674 27464
rect 20254 27452 20260 27464
rect 20215 27424 20260 27452
rect 20254 27412 20260 27424
rect 20312 27412 20318 27464
rect 20346 27412 20352 27464
rect 20404 27452 20410 27464
rect 20809 27455 20867 27461
rect 20809 27452 20821 27455
rect 20404 27424 20821 27452
rect 20404 27412 20410 27424
rect 20809 27421 20821 27424
rect 20855 27421 20867 27455
rect 21358 27452 21364 27464
rect 21319 27424 21364 27452
rect 20809 27415 20867 27421
rect 21358 27412 21364 27424
rect 21416 27412 21422 27464
rect 22186 27452 22192 27464
rect 22147 27424 22192 27452
rect 22186 27412 22192 27424
rect 22244 27412 22250 27464
rect 22741 27455 22799 27461
rect 22480 27424 22692 27452
rect 10962 27384 10968 27396
rect 1596 27356 10180 27384
rect 10244 27356 10968 27384
rect 1596 27325 1624 27356
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27285 1639 27319
rect 1581 27279 1639 27285
rect 1670 27276 1676 27328
rect 1728 27316 1734 27328
rect 2041 27319 2099 27325
rect 2041 27316 2053 27319
rect 1728 27288 2053 27316
rect 1728 27276 1734 27288
rect 2041 27285 2053 27288
rect 2087 27285 2099 27319
rect 2041 27279 2099 27285
rect 3973 27319 4031 27325
rect 3973 27285 3985 27319
rect 4019 27316 4031 27319
rect 4062 27316 4068 27328
rect 4019 27288 4068 27316
rect 4019 27285 4031 27288
rect 3973 27279 4031 27285
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 4798 27316 4804 27328
rect 4759 27288 4804 27316
rect 4798 27276 4804 27288
rect 4856 27276 4862 27328
rect 9674 27316 9680 27328
rect 9635 27288 9680 27316
rect 9674 27276 9680 27288
rect 9732 27276 9738 27328
rect 10152 27316 10180 27356
rect 10962 27344 10968 27356
rect 11020 27344 11026 27396
rect 12158 27344 12164 27396
rect 12216 27384 12222 27396
rect 17126 27384 17132 27396
rect 12216 27356 17132 27384
rect 12216 27344 12222 27356
rect 17126 27344 17132 27356
rect 17184 27344 17190 27396
rect 20438 27384 20444 27396
rect 17236 27356 20444 27384
rect 17236 27316 17264 27356
rect 20438 27344 20444 27356
rect 20496 27344 20502 27396
rect 22480 27384 22508 27424
rect 21192 27356 22508 27384
rect 22664 27384 22692 27424
rect 22741 27421 22753 27455
rect 22787 27452 22799 27455
rect 22830 27452 22836 27464
rect 22787 27424 22836 27452
rect 22787 27421 22799 27424
rect 22741 27415 22799 27421
rect 22830 27412 22836 27424
rect 22888 27412 22894 27464
rect 23382 27452 23388 27464
rect 23343 27424 23388 27452
rect 23382 27412 23388 27424
rect 23440 27412 23446 27464
rect 24578 27412 24584 27464
rect 24636 27452 24642 27464
rect 24765 27455 24823 27461
rect 24765 27452 24777 27455
rect 24636 27424 24777 27452
rect 24636 27412 24642 27424
rect 24765 27421 24777 27424
rect 24811 27421 24823 27455
rect 24765 27415 24823 27421
rect 25501 27455 25559 27461
rect 25501 27421 25513 27455
rect 25547 27421 25559 27455
rect 25958 27452 25964 27464
rect 25919 27424 25964 27452
rect 25501 27415 25559 27421
rect 25406 27384 25412 27396
rect 22664 27356 25412 27384
rect 10152 27288 17264 27316
rect 19429 27319 19487 27325
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 19794 27316 19800 27328
rect 19475 27288 19800 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 19794 27276 19800 27288
rect 19852 27276 19858 27328
rect 21192 27325 21220 27356
rect 25406 27344 25412 27356
rect 25464 27344 25470 27396
rect 25516 27384 25544 27415
rect 25958 27412 25964 27424
rect 26016 27412 26022 27464
rect 26694 27412 26700 27464
rect 26752 27452 26758 27464
rect 27341 27455 27399 27461
rect 27341 27452 27353 27455
rect 26752 27424 27353 27452
rect 26752 27412 26758 27424
rect 27341 27421 27353 27424
rect 27387 27421 27399 27455
rect 27341 27415 27399 27421
rect 27985 27455 28043 27461
rect 27985 27421 27997 27455
rect 28031 27452 28043 27455
rect 28166 27452 28172 27464
rect 28031 27424 28172 27452
rect 28031 27421 28043 27424
rect 27985 27415 28043 27421
rect 28166 27412 28172 27424
rect 28224 27412 28230 27464
rect 28350 27412 28356 27464
rect 28408 27452 28414 27464
rect 28537 27455 28595 27461
rect 28537 27452 28549 27455
rect 28408 27424 28549 27452
rect 28408 27412 28414 27424
rect 28537 27421 28549 27424
rect 28583 27421 28595 27455
rect 29086 27452 29092 27464
rect 29047 27424 29092 27452
rect 28537 27415 28595 27421
rect 29086 27412 29092 27424
rect 29144 27412 29150 27464
rect 29914 27452 29920 27464
rect 29875 27424 29920 27452
rect 29914 27412 29920 27424
rect 29972 27412 29978 27464
rect 31110 27452 31116 27464
rect 31071 27424 31116 27452
rect 31110 27412 31116 27424
rect 31168 27412 31174 27464
rect 31846 27412 31852 27464
rect 31904 27452 31910 27464
rect 32125 27455 32183 27461
rect 32125 27452 32137 27455
rect 31904 27424 32137 27452
rect 31904 27412 31910 27424
rect 32125 27421 32137 27424
rect 32171 27421 32183 27455
rect 33686 27452 33692 27464
rect 33647 27424 33692 27452
rect 32125 27415 32183 27421
rect 33686 27412 33692 27424
rect 33744 27412 33750 27464
rect 34238 27452 34244 27464
rect 34199 27424 34244 27452
rect 34238 27412 34244 27424
rect 34296 27412 34302 27464
rect 35066 27452 35072 27464
rect 35027 27424 35072 27452
rect 35066 27412 35072 27424
rect 35124 27412 35130 27464
rect 35710 27452 35716 27464
rect 35671 27424 35716 27452
rect 35710 27412 35716 27424
rect 35768 27412 35774 27464
rect 36265 27455 36323 27461
rect 36265 27421 36277 27455
rect 36311 27421 36323 27455
rect 36814 27452 36820 27464
rect 36775 27424 36820 27452
rect 36265 27415 36323 27421
rect 27246 27384 27252 27396
rect 25516 27356 27252 27384
rect 27246 27344 27252 27356
rect 27304 27344 27310 27396
rect 27356 27356 29040 27384
rect 21177 27319 21235 27325
rect 21177 27285 21189 27319
rect 21223 27285 21235 27319
rect 21177 27279 21235 27285
rect 21266 27276 21272 27328
rect 21324 27316 21330 27328
rect 25866 27316 25872 27328
rect 21324 27288 25872 27316
rect 21324 27276 21330 27288
rect 25866 27276 25872 27288
rect 25924 27276 25930 27328
rect 26050 27316 26056 27328
rect 26011 27288 26056 27316
rect 26050 27276 26056 27288
rect 26108 27276 26114 27328
rect 26234 27276 26240 27328
rect 26292 27316 26298 27328
rect 27356 27316 27384 27356
rect 26292 27288 27384 27316
rect 26292 27276 26298 27288
rect 28074 27276 28080 27328
rect 28132 27316 28138 27328
rect 28353 27319 28411 27325
rect 28353 27316 28365 27319
rect 28132 27288 28365 27316
rect 28132 27276 28138 27288
rect 28353 27285 28365 27288
rect 28399 27285 28411 27319
rect 28353 27279 28411 27285
rect 28534 27276 28540 27328
rect 28592 27316 28598 27328
rect 28905 27319 28963 27325
rect 28905 27316 28917 27319
rect 28592 27288 28917 27316
rect 28592 27276 28598 27288
rect 28905 27285 28917 27288
rect 28951 27285 28963 27319
rect 29012 27316 29040 27356
rect 31938 27344 31944 27396
rect 31996 27384 32002 27396
rect 36170 27384 36176 27396
rect 31996 27356 36176 27384
rect 31996 27344 32002 27356
rect 36170 27344 36176 27356
rect 36228 27344 36234 27396
rect 36280 27384 36308 27415
rect 36814 27412 36820 27424
rect 36872 27412 36878 27464
rect 37274 27412 37280 27464
rect 37332 27452 37338 27464
rect 37645 27455 37703 27461
rect 37645 27452 37657 27455
rect 37332 27424 37657 27452
rect 37332 27412 37338 27424
rect 37645 27421 37657 27424
rect 37691 27452 37703 27455
rect 37826 27452 37832 27464
rect 37691 27424 37832 27452
rect 37691 27421 37703 27424
rect 37645 27415 37703 27421
rect 37826 27412 37832 27424
rect 37884 27412 37890 27464
rect 37918 27412 37924 27464
rect 37976 27452 37982 27464
rect 38289 27455 38347 27461
rect 38289 27452 38301 27455
rect 37976 27424 38301 27452
rect 37976 27412 37982 27424
rect 38289 27421 38301 27424
rect 38335 27421 38347 27455
rect 38289 27415 38347 27421
rect 38933 27455 38991 27461
rect 38933 27421 38945 27455
rect 38979 27452 38991 27455
rect 39114 27452 39120 27464
rect 38979 27424 39120 27452
rect 38979 27421 38991 27424
rect 38933 27415 38991 27421
rect 39114 27412 39120 27424
rect 39172 27412 39178 27464
rect 39850 27412 39856 27464
rect 39908 27412 39914 27464
rect 40052 27461 40080 27492
rect 40037 27455 40095 27461
rect 40037 27421 40049 27455
rect 40083 27421 40095 27455
rect 40037 27415 40095 27421
rect 40678 27412 40684 27464
rect 40736 27452 40742 27464
rect 40865 27455 40923 27461
rect 40865 27452 40877 27455
rect 40736 27424 40877 27452
rect 40736 27412 40742 27424
rect 40865 27421 40877 27424
rect 40911 27421 40923 27455
rect 40865 27415 40923 27421
rect 41417 27455 41475 27461
rect 41417 27421 41429 27455
rect 41463 27452 41475 27455
rect 41598 27452 41604 27464
rect 41463 27424 41604 27452
rect 41463 27421 41475 27424
rect 41417 27415 41475 27421
rect 41598 27412 41604 27424
rect 41656 27412 41662 27464
rect 41966 27452 41972 27464
rect 41927 27424 41972 27452
rect 41966 27412 41972 27424
rect 42024 27412 42030 27464
rect 42076 27452 42104 27492
rect 42518 27480 42524 27532
rect 42576 27520 42582 27532
rect 86126 27520 86132 27532
rect 42576 27492 86132 27520
rect 42576 27480 42582 27492
rect 86126 27480 86132 27492
rect 86184 27480 86190 27532
rect 42702 27452 42708 27464
rect 42076 27424 42708 27452
rect 42702 27412 42708 27424
rect 42760 27412 42766 27464
rect 42794 27412 42800 27464
rect 42852 27452 42858 27464
rect 43438 27452 43444 27464
rect 42852 27424 42897 27452
rect 43399 27424 43444 27452
rect 42852 27412 42858 27424
rect 43438 27412 43444 27424
rect 43496 27412 43502 27464
rect 43990 27452 43996 27464
rect 43951 27424 43996 27452
rect 43990 27412 43996 27424
rect 44048 27412 44054 27464
rect 44542 27452 44548 27464
rect 44503 27424 44548 27452
rect 44542 27412 44548 27424
rect 44600 27412 44606 27464
rect 45370 27452 45376 27464
rect 45331 27424 45376 27452
rect 45370 27412 45376 27424
rect 45428 27412 45434 27464
rect 45462 27412 45468 27464
rect 45520 27452 45526 27464
rect 46017 27455 46075 27461
rect 46017 27452 46029 27455
rect 45520 27424 46029 27452
rect 45520 27412 45526 27424
rect 46017 27421 46029 27424
rect 46063 27421 46075 27455
rect 46658 27452 46664 27464
rect 46619 27424 46664 27452
rect 46017 27415 46075 27421
rect 46658 27412 46664 27424
rect 46716 27412 46722 27464
rect 48590 27452 48596 27464
rect 48551 27424 48596 27452
rect 48590 27412 48596 27424
rect 48648 27412 48654 27464
rect 49050 27412 49056 27464
rect 49108 27452 49114 27464
rect 49237 27455 49295 27461
rect 49237 27452 49249 27455
rect 49108 27424 49249 27452
rect 49108 27412 49114 27424
rect 49237 27421 49249 27424
rect 49283 27421 49295 27455
rect 50522 27452 50528 27464
rect 50483 27424 50528 27452
rect 49237 27415 49295 27421
rect 50522 27412 50528 27424
rect 50580 27412 50586 27464
rect 51261 27455 51319 27461
rect 51261 27421 51273 27455
rect 51307 27421 51319 27455
rect 51810 27452 51816 27464
rect 51771 27424 51816 27452
rect 51261 27415 51319 27421
rect 42610 27384 42616 27396
rect 36280 27356 42616 27384
rect 42610 27344 42616 27356
rect 42668 27344 42674 27396
rect 46750 27344 46756 27396
rect 46808 27384 46814 27396
rect 51166 27384 51172 27396
rect 46808 27356 51172 27384
rect 46808 27344 46814 27356
rect 51166 27344 51172 27356
rect 51224 27344 51230 27396
rect 51276 27384 51304 27415
rect 51810 27412 51816 27424
rect 51868 27412 51874 27464
rect 52914 27452 52920 27464
rect 52875 27424 52920 27452
rect 52914 27412 52920 27424
rect 52972 27412 52978 27464
rect 53558 27452 53564 27464
rect 53519 27424 53564 27452
rect 53558 27412 53564 27424
rect 53616 27412 53622 27464
rect 53837 27455 53895 27461
rect 53837 27421 53849 27455
rect 53883 27452 53895 27455
rect 54018 27452 54024 27464
rect 53883 27424 54024 27452
rect 53883 27421 53895 27424
rect 53837 27415 53895 27421
rect 54018 27412 54024 27424
rect 54076 27412 54082 27464
rect 56321 27455 56379 27461
rect 56321 27421 56333 27455
rect 56367 27421 56379 27455
rect 56321 27415 56379 27421
rect 56965 27455 57023 27461
rect 56965 27421 56977 27455
rect 57011 27421 57023 27455
rect 56965 27415 57023 27421
rect 51718 27384 51724 27396
rect 51276 27356 51724 27384
rect 51718 27344 51724 27356
rect 51776 27344 51782 27396
rect 52730 27344 52736 27396
rect 52788 27384 52794 27396
rect 56336 27384 56364 27415
rect 52788 27356 56364 27384
rect 52788 27344 52794 27356
rect 56980 27328 57008 27415
rect 57054 27412 57060 27464
rect 57112 27452 57118 27464
rect 58069 27455 58127 27461
rect 58069 27452 58081 27455
rect 57112 27424 58081 27452
rect 57112 27412 57118 27424
rect 58069 27421 58081 27424
rect 58115 27421 58127 27455
rect 58802 27452 58808 27464
rect 58763 27424 58808 27452
rect 58069 27415 58127 27421
rect 58802 27412 58808 27424
rect 58860 27412 58866 27464
rect 59541 27455 59599 27461
rect 59541 27421 59553 27455
rect 59587 27421 59599 27455
rect 59541 27415 59599 27421
rect 58618 27344 58624 27396
rect 58676 27384 58682 27396
rect 59556 27384 59584 27415
rect 59630 27412 59636 27464
rect 59688 27452 59694 27464
rect 60645 27455 60703 27461
rect 60645 27452 60657 27455
rect 59688 27424 60657 27452
rect 59688 27412 59694 27424
rect 60645 27421 60657 27424
rect 60691 27421 60703 27455
rect 61286 27452 61292 27464
rect 61247 27424 61292 27452
rect 60645 27415 60703 27421
rect 61286 27412 61292 27424
rect 61344 27412 61350 27464
rect 61378 27412 61384 27464
rect 61436 27452 61442 27464
rect 62117 27455 62175 27461
rect 62117 27452 62129 27455
rect 61436 27424 62129 27452
rect 61436 27412 61442 27424
rect 62117 27421 62129 27424
rect 62163 27421 62175 27455
rect 62117 27415 62175 27421
rect 63221 27455 63279 27461
rect 63221 27421 63233 27455
rect 63267 27421 63279 27455
rect 63862 27452 63868 27464
rect 63823 27424 63868 27452
rect 63221 27415 63279 27421
rect 58676 27356 59584 27384
rect 58676 27344 58682 27356
rect 59998 27344 60004 27396
rect 60056 27384 60062 27396
rect 60056 27356 61516 27384
rect 60056 27344 60062 27356
rect 41046 27316 41052 27328
rect 29012 27288 41052 27316
rect 28905 27279 28963 27285
rect 41046 27276 41052 27288
rect 41104 27276 41110 27328
rect 41230 27316 41236 27328
rect 41191 27288 41236 27316
rect 41230 27276 41236 27288
rect 41288 27276 41294 27328
rect 41785 27319 41843 27325
rect 41785 27285 41797 27319
rect 41831 27316 41843 27319
rect 42886 27316 42892 27328
rect 41831 27288 42892 27316
rect 41831 27285 41843 27288
rect 41785 27279 41843 27285
rect 42886 27276 42892 27288
rect 42944 27276 42950 27328
rect 43530 27276 43536 27328
rect 43588 27316 43594 27328
rect 44361 27319 44419 27325
rect 44361 27316 44373 27319
rect 43588 27288 44373 27316
rect 43588 27276 43594 27288
rect 44361 27285 44373 27288
rect 44407 27285 44419 27319
rect 44361 27279 44419 27285
rect 48314 27276 48320 27328
rect 48372 27316 48378 27328
rect 48409 27319 48467 27325
rect 48409 27316 48421 27319
rect 48372 27288 48421 27316
rect 48372 27276 48378 27288
rect 48409 27285 48421 27288
rect 48455 27285 48467 27319
rect 48409 27279 48467 27285
rect 50430 27276 50436 27328
rect 50488 27316 50494 27328
rect 50617 27319 50675 27325
rect 50617 27316 50629 27319
rect 50488 27288 50629 27316
rect 50488 27276 50494 27288
rect 50617 27285 50629 27288
rect 50663 27285 50675 27319
rect 50617 27279 50675 27285
rect 51629 27319 51687 27325
rect 51629 27285 51641 27319
rect 51675 27316 51687 27319
rect 52086 27316 52092 27328
rect 51675 27288 52092 27316
rect 51675 27285 51687 27288
rect 51629 27279 51687 27285
rect 52086 27276 52092 27288
rect 52144 27276 52150 27328
rect 52270 27276 52276 27328
rect 52328 27316 52334 27328
rect 53190 27316 53196 27328
rect 52328 27288 53196 27316
rect 52328 27276 52334 27288
rect 53190 27276 53196 27288
rect 53248 27276 53254 27328
rect 54294 27276 54300 27328
rect 54352 27316 54358 27328
rect 56962 27316 56968 27328
rect 54352 27288 56968 27316
rect 54352 27276 54358 27288
rect 56962 27276 56968 27288
rect 57020 27276 57026 27328
rect 58710 27276 58716 27328
rect 58768 27316 58774 27328
rect 58897 27319 58955 27325
rect 58897 27316 58909 27319
rect 58768 27288 58909 27316
rect 58768 27276 58774 27288
rect 58897 27285 58909 27288
rect 58943 27285 58955 27319
rect 58897 27279 58955 27285
rect 59262 27276 59268 27328
rect 59320 27316 59326 27328
rect 60550 27316 60556 27328
rect 59320 27288 60556 27316
rect 59320 27276 59326 27288
rect 60550 27276 60556 27288
rect 60608 27276 60614 27328
rect 61488 27316 61516 27356
rect 61562 27344 61568 27396
rect 61620 27384 61626 27396
rect 63236 27384 63264 27415
rect 63862 27412 63868 27424
rect 63920 27412 63926 27464
rect 64141 27455 64199 27461
rect 64141 27421 64153 27455
rect 64187 27421 64199 27455
rect 64141 27415 64199 27421
rect 61620 27356 63264 27384
rect 61620 27344 61626 27356
rect 64156 27316 64184 27415
rect 64414 27412 64420 27464
rect 64472 27452 64478 27464
rect 65797 27455 65855 27461
rect 65797 27452 65809 27455
rect 64472 27424 65809 27452
rect 64472 27412 64478 27424
rect 65797 27421 65809 27424
rect 65843 27421 65855 27455
rect 65797 27415 65855 27421
rect 66254 27412 66260 27464
rect 66312 27452 66318 27464
rect 66349 27455 66407 27461
rect 66349 27452 66361 27455
rect 66312 27424 66361 27452
rect 66312 27412 66318 27424
rect 66349 27421 66361 27424
rect 66395 27421 66407 27455
rect 66349 27415 66407 27421
rect 66438 27412 66444 27464
rect 66496 27452 66502 27464
rect 66901 27455 66959 27461
rect 66901 27452 66913 27455
rect 66496 27424 66913 27452
rect 66496 27412 66502 27424
rect 66901 27421 66913 27424
rect 66947 27421 66959 27455
rect 66901 27415 66959 27421
rect 66990 27412 66996 27464
rect 67048 27452 67054 27464
rect 67453 27455 67511 27461
rect 67453 27452 67465 27455
rect 67048 27424 67465 27452
rect 67048 27412 67054 27424
rect 67453 27421 67465 27424
rect 67499 27421 67511 27455
rect 67453 27415 67511 27421
rect 67634 27412 67640 27464
rect 67692 27452 67698 27464
rect 68557 27455 68615 27461
rect 68557 27452 68569 27455
rect 67692 27424 68569 27452
rect 67692 27412 67698 27424
rect 68557 27421 68569 27424
rect 68603 27421 68615 27455
rect 68557 27415 68615 27421
rect 68646 27412 68652 27464
rect 68704 27452 68710 27464
rect 69293 27455 69351 27461
rect 69293 27452 69305 27455
rect 68704 27424 69305 27452
rect 68704 27412 68710 27424
rect 69293 27421 69305 27424
rect 69339 27421 69351 27455
rect 69293 27415 69351 27421
rect 69382 27412 69388 27464
rect 69440 27452 69446 27464
rect 69845 27455 69903 27461
rect 69845 27452 69857 27455
rect 69440 27424 69857 27452
rect 69440 27412 69446 27424
rect 69845 27421 69857 27424
rect 69891 27421 69903 27455
rect 69845 27415 69903 27421
rect 70854 27412 70860 27464
rect 70912 27452 70918 27464
rect 70949 27455 71007 27461
rect 70949 27452 70961 27455
rect 70912 27424 70961 27452
rect 70912 27412 70918 27424
rect 70949 27421 70961 27424
rect 70995 27421 71007 27455
rect 71498 27452 71504 27464
rect 71459 27424 71504 27452
rect 70949 27415 71007 27421
rect 71498 27412 71504 27424
rect 71556 27412 71562 27464
rect 72050 27452 72056 27464
rect 72011 27424 72056 27452
rect 72050 27412 72056 27424
rect 72108 27412 72114 27464
rect 72605 27455 72663 27461
rect 72605 27421 72617 27455
rect 72651 27421 72663 27455
rect 73706 27452 73712 27464
rect 73667 27424 73712 27452
rect 72605 27415 72663 27421
rect 68186 27344 68192 27396
rect 68244 27384 68250 27396
rect 68244 27356 69152 27384
rect 68244 27344 68250 27356
rect 61488 27288 64184 27316
rect 67269 27319 67327 27325
rect 67269 27285 67281 27319
rect 67315 27316 67327 27319
rect 67450 27316 67456 27328
rect 67315 27288 67456 27316
rect 67315 27285 67327 27288
rect 67269 27279 67327 27285
rect 67450 27276 67456 27288
rect 67508 27276 67514 27328
rect 68646 27316 68652 27328
rect 68607 27288 68652 27316
rect 68646 27276 68652 27288
rect 68704 27276 68710 27328
rect 69124 27325 69152 27356
rect 69474 27344 69480 27396
rect 69532 27384 69538 27396
rect 72620 27384 72648 27415
rect 73706 27412 73712 27424
rect 73764 27412 73770 27464
rect 74442 27452 74448 27464
rect 74403 27424 74448 27452
rect 74442 27412 74448 27424
rect 74500 27412 74506 27464
rect 74997 27455 75055 27461
rect 74997 27421 75009 27455
rect 75043 27421 75055 27455
rect 76282 27452 76288 27464
rect 76243 27424 76288 27452
rect 74997 27415 75055 27421
rect 75012 27384 75040 27415
rect 76282 27412 76288 27424
rect 76340 27412 76346 27464
rect 76374 27412 76380 27464
rect 76432 27452 76438 27464
rect 76469 27455 76527 27461
rect 76469 27452 76481 27455
rect 76432 27424 76481 27452
rect 76432 27412 76438 27424
rect 76469 27421 76481 27424
rect 76515 27421 76527 27455
rect 76469 27415 76527 27421
rect 77021 27455 77079 27461
rect 77021 27421 77033 27455
rect 77067 27421 77079 27455
rect 77021 27415 77079 27421
rect 77573 27455 77631 27461
rect 77573 27421 77585 27455
rect 77619 27421 77631 27455
rect 77573 27415 77631 27421
rect 69532 27356 72648 27384
rect 72712 27356 75040 27384
rect 69532 27344 69538 27356
rect 69109 27319 69167 27325
rect 69109 27285 69121 27319
rect 69155 27285 69167 27319
rect 69109 27279 69167 27285
rect 69842 27276 69848 27328
rect 69900 27316 69906 27328
rect 70765 27319 70823 27325
rect 70765 27316 70777 27319
rect 69900 27288 70777 27316
rect 69900 27276 69906 27288
rect 70765 27285 70777 27288
rect 70811 27285 70823 27319
rect 70765 27279 70823 27285
rect 72510 27276 72516 27328
rect 72568 27316 72574 27328
rect 72712 27316 72740 27356
rect 75086 27344 75092 27396
rect 75144 27384 75150 27396
rect 77036 27384 77064 27415
rect 75144 27356 77064 27384
rect 75144 27344 75150 27356
rect 73798 27316 73804 27328
rect 72568 27288 72740 27316
rect 73759 27288 73804 27316
rect 72568 27276 72574 27288
rect 73798 27276 73804 27288
rect 73856 27276 73862 27328
rect 75178 27276 75184 27328
rect 75236 27316 75242 27328
rect 77588 27316 77616 27415
rect 78306 27412 78312 27464
rect 78364 27452 78370 27464
rect 78861 27455 78919 27461
rect 78861 27452 78873 27455
rect 78364 27424 78873 27452
rect 78364 27412 78370 27424
rect 78861 27421 78873 27424
rect 78907 27421 78919 27455
rect 79410 27452 79416 27464
rect 79371 27424 79416 27452
rect 78861 27415 78919 27421
rect 79410 27412 79416 27424
rect 79468 27412 79474 27464
rect 80054 27452 80060 27464
rect 80015 27424 80060 27452
rect 80054 27412 80060 27424
rect 80112 27412 80118 27464
rect 81434 27452 81440 27464
rect 81395 27424 81440 27452
rect 81434 27412 81440 27424
rect 81492 27412 81498 27464
rect 82170 27452 82176 27464
rect 82131 27424 82176 27452
rect 82170 27412 82176 27424
rect 82228 27412 82234 27464
rect 82538 27452 82544 27464
rect 82499 27424 82544 27452
rect 82538 27412 82544 27424
rect 82596 27412 82602 27464
rect 83826 27452 83832 27464
rect 83787 27424 83832 27452
rect 83826 27412 83832 27424
rect 83884 27412 83890 27464
rect 84194 27412 84200 27464
rect 84252 27452 84258 27464
rect 84381 27455 84439 27461
rect 84381 27452 84393 27455
rect 84252 27424 84393 27452
rect 84252 27412 84258 27424
rect 84381 27421 84393 27424
rect 84427 27421 84439 27455
rect 85114 27452 85120 27464
rect 85075 27424 85120 27452
rect 84381 27415 84439 27421
rect 85114 27412 85120 27424
rect 85172 27412 85178 27464
rect 86402 27452 86408 27464
rect 86363 27424 86408 27452
rect 86402 27412 86408 27424
rect 86460 27412 86466 27464
rect 86788 27461 86816 27560
rect 89530 27548 89536 27560
rect 89588 27548 89594 27600
rect 87417 27523 87475 27529
rect 87417 27489 87429 27523
rect 87463 27520 87475 27523
rect 87598 27520 87604 27532
rect 87463 27492 87604 27520
rect 87463 27489 87475 27492
rect 87417 27483 87475 27489
rect 87598 27480 87604 27492
rect 87656 27480 87662 27532
rect 86773 27455 86831 27461
rect 86773 27421 86785 27455
rect 86819 27421 86831 27455
rect 86773 27415 86831 27421
rect 87693 27455 87751 27461
rect 87693 27421 87705 27455
rect 87739 27452 87751 27455
rect 87782 27452 87788 27464
rect 87739 27424 87788 27452
rect 87739 27421 87751 27424
rect 87693 27415 87751 27421
rect 87782 27412 87788 27424
rect 87840 27412 87846 27464
rect 78122 27344 78128 27396
rect 78180 27384 78186 27396
rect 78180 27356 84240 27384
rect 78180 27344 78186 27356
rect 78950 27316 78956 27328
rect 75236 27288 77616 27316
rect 78911 27288 78956 27316
rect 75236 27276 75242 27288
rect 78950 27276 78956 27288
rect 79008 27276 79014 27328
rect 79594 27316 79600 27328
rect 79555 27288 79600 27316
rect 79594 27276 79600 27288
rect 79652 27276 79658 27328
rect 80238 27316 80244 27328
rect 80199 27288 80244 27316
rect 80238 27276 80244 27288
rect 80296 27276 80302 27328
rect 81526 27316 81532 27328
rect 81487 27288 81532 27316
rect 81526 27276 81532 27288
rect 81584 27276 81590 27328
rect 82722 27316 82728 27328
rect 82683 27288 82728 27316
rect 82722 27276 82728 27288
rect 82780 27276 82786 27328
rect 84212 27325 84240 27356
rect 84197 27319 84255 27325
rect 84197 27285 84209 27319
rect 84243 27285 84255 27319
rect 84197 27279 84255 27285
rect 86957 27319 87015 27325
rect 86957 27285 86969 27319
rect 87003 27316 87015 27319
rect 87874 27316 87880 27328
rect 87003 27288 87880 27316
rect 87003 27285 87015 27288
rect 86957 27279 87015 27285
rect 87874 27276 87880 27288
rect 87932 27276 87938 27328
rect 1104 27226 88872 27248
rect 1104 27174 22898 27226
rect 22950 27174 22962 27226
rect 23014 27174 23026 27226
rect 23078 27174 23090 27226
rect 23142 27174 23154 27226
rect 23206 27174 44846 27226
rect 44898 27174 44910 27226
rect 44962 27174 44974 27226
rect 45026 27174 45038 27226
rect 45090 27174 45102 27226
rect 45154 27174 66794 27226
rect 66846 27174 66858 27226
rect 66910 27174 66922 27226
rect 66974 27174 66986 27226
rect 67038 27174 67050 27226
rect 67102 27174 88872 27226
rect 1104 27152 88872 27174
rect 14 27072 20 27124
rect 72 27112 78 27124
rect 2593 27115 2651 27121
rect 2593 27112 2605 27115
rect 72 27084 2605 27112
rect 72 27072 78 27084
rect 2593 27081 2605 27084
rect 2639 27081 2651 27115
rect 2593 27075 2651 27081
rect 3050 27072 3056 27124
rect 3108 27112 3114 27124
rect 3145 27115 3203 27121
rect 3145 27112 3157 27115
rect 3108 27084 3157 27112
rect 3108 27072 3114 27084
rect 3145 27081 3157 27084
rect 3191 27081 3203 27115
rect 3970 27112 3976 27124
rect 3931 27084 3976 27112
rect 3145 27075 3203 27081
rect 3970 27072 3976 27084
rect 4028 27072 4034 27124
rect 7282 27112 7288 27124
rect 7243 27084 7288 27112
rect 7282 27072 7288 27084
rect 7340 27072 7346 27124
rect 10410 27112 10416 27124
rect 10371 27084 10416 27112
rect 10410 27072 10416 27084
rect 10468 27072 10474 27124
rect 13630 27112 13636 27124
rect 13591 27084 13636 27112
rect 13630 27072 13636 27084
rect 13688 27072 13694 27124
rect 18782 27072 18788 27124
rect 18840 27112 18846 27124
rect 19797 27115 19855 27121
rect 19797 27112 19809 27115
rect 18840 27084 19809 27112
rect 18840 27072 18846 27084
rect 19797 27081 19809 27084
rect 19843 27081 19855 27115
rect 20346 27112 20352 27124
rect 20307 27084 20352 27112
rect 19797 27075 19855 27081
rect 20346 27072 20352 27084
rect 20404 27072 20410 27124
rect 20438 27072 20444 27124
rect 20496 27112 20502 27124
rect 32950 27112 32956 27124
rect 20496 27084 32812 27112
rect 32911 27084 32956 27112
rect 20496 27072 20502 27084
rect 1762 27044 1768 27056
rect 1723 27016 1768 27044
rect 1762 27004 1768 27016
rect 1820 27004 1826 27056
rect 6730 27044 6736 27056
rect 6691 27016 6736 27044
rect 6730 27004 6736 27016
rect 6788 27004 6794 27056
rect 10502 27004 10508 27056
rect 10560 27044 10566 27056
rect 13538 27044 13544 27056
rect 10560 27016 13544 27044
rect 10560 27004 10566 27016
rect 13538 27004 13544 27016
rect 13596 27004 13602 27056
rect 15654 27044 15660 27056
rect 13740 27016 15660 27044
rect 2317 26979 2375 26985
rect 2317 26945 2329 26979
rect 2363 26976 2375 26979
rect 2777 26979 2835 26985
rect 2777 26976 2789 26979
rect 2363 26948 2789 26976
rect 2363 26945 2375 26948
rect 2317 26939 2375 26945
rect 2777 26945 2789 26948
rect 2823 26976 2835 26979
rect 2866 26976 2872 26988
rect 2823 26948 2872 26976
rect 2823 26945 2835 26948
rect 2777 26939 2835 26945
rect 2866 26936 2872 26948
rect 2924 26936 2930 26988
rect 3329 26979 3387 26985
rect 3329 26945 3341 26979
rect 3375 26945 3387 26979
rect 4154 26976 4160 26988
rect 4115 26948 4160 26976
rect 3329 26939 3387 26945
rect 3344 26908 3372 26939
rect 4154 26936 4160 26948
rect 4212 26936 4218 26988
rect 7466 26976 7472 26988
rect 7427 26948 7472 26976
rect 7466 26936 7472 26948
rect 7524 26936 7530 26988
rect 10594 26976 10600 26988
rect 10555 26948 10600 26976
rect 10594 26936 10600 26948
rect 10652 26936 10658 26988
rect 12342 26976 12348 26988
rect 12303 26948 12348 26976
rect 12342 26936 12348 26948
rect 12400 26936 12406 26988
rect 13740 26908 13768 27016
rect 15654 27004 15660 27016
rect 15712 27004 15718 27056
rect 15746 27004 15752 27056
rect 15804 27044 15810 27056
rect 32674 27044 32680 27056
rect 15804 27016 32680 27044
rect 15804 27004 15810 27016
rect 32674 27004 32680 27016
rect 32732 27004 32738 27056
rect 32784 27044 32812 27084
rect 32950 27072 32956 27084
rect 33008 27072 33014 27124
rect 33042 27072 33048 27124
rect 33100 27112 33106 27124
rect 37550 27112 37556 27124
rect 33100 27084 37556 27112
rect 33100 27072 33106 27084
rect 37550 27072 37556 27084
rect 37608 27072 37614 27124
rect 37918 27112 37924 27124
rect 37879 27084 37924 27112
rect 37918 27072 37924 27084
rect 37976 27072 37982 27124
rect 38010 27072 38016 27124
rect 38068 27112 38074 27124
rect 38289 27115 38347 27121
rect 38289 27112 38301 27115
rect 38068 27084 38301 27112
rect 38068 27072 38074 27084
rect 38289 27081 38301 27084
rect 38335 27112 38347 27115
rect 40221 27115 40279 27121
rect 40221 27112 40233 27115
rect 38335 27084 40233 27112
rect 38335 27081 38347 27084
rect 38289 27075 38347 27081
rect 40221 27081 40233 27084
rect 40267 27081 40279 27115
rect 40678 27112 40684 27124
rect 40639 27084 40684 27112
rect 40221 27075 40279 27081
rect 40678 27072 40684 27084
rect 40736 27072 40742 27124
rect 42518 27112 42524 27124
rect 41386 27084 42524 27112
rect 35526 27044 35532 27056
rect 32784 27016 35532 27044
rect 35526 27004 35532 27016
rect 35584 27004 35590 27056
rect 38120 27016 38516 27044
rect 38120 26988 38148 27016
rect 13817 26979 13875 26985
rect 13817 26945 13829 26979
rect 13863 26976 13875 26979
rect 14734 26976 14740 26988
rect 13863 26948 14596 26976
rect 14695 26948 14740 26976
rect 13863 26945 13875 26948
rect 13817 26939 13875 26945
rect 3344 26880 13768 26908
rect 1949 26843 2007 26849
rect 1949 26809 1961 26843
rect 1995 26840 2007 26843
rect 2038 26840 2044 26852
rect 1995 26812 2044 26840
rect 1995 26809 2007 26812
rect 1949 26803 2007 26809
rect 2038 26800 2044 26812
rect 2096 26800 2102 26852
rect 6914 26800 6920 26852
rect 6972 26840 6978 26852
rect 6972 26812 7017 26840
rect 6972 26800 6978 26812
rect 9674 26800 9680 26852
rect 9732 26840 9738 26852
rect 14568 26849 14596 26948
rect 14734 26936 14740 26948
rect 14792 26936 14798 26988
rect 17034 26976 17040 26988
rect 16995 26948 17040 26976
rect 17034 26936 17040 26948
rect 17092 26936 17098 26988
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 19426 26976 19432 26988
rect 18104 26948 19432 26976
rect 18104 26936 18110 26948
rect 19426 26936 19432 26948
rect 19484 26936 19490 26988
rect 19521 26979 19579 26985
rect 19521 26945 19533 26979
rect 19567 26976 19579 26979
rect 19978 26976 19984 26988
rect 19567 26948 19984 26976
rect 19567 26945 19579 26948
rect 19521 26939 19579 26945
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 20438 26936 20444 26988
rect 20496 26976 20502 26988
rect 20533 26979 20591 26985
rect 20533 26976 20545 26979
rect 20496 26948 20545 26976
rect 20496 26936 20502 26948
rect 20533 26945 20545 26948
rect 20579 26945 20591 26979
rect 20533 26939 20591 26945
rect 22186 26936 22192 26988
rect 22244 26976 22250 26988
rect 23934 26976 23940 26988
rect 22244 26948 23940 26976
rect 22244 26936 22250 26948
rect 23934 26936 23940 26948
rect 23992 26936 23998 26988
rect 24118 26976 24124 26988
rect 24079 26948 24124 26976
rect 24118 26936 24124 26948
rect 24176 26936 24182 26988
rect 26234 26976 26240 26988
rect 26068 26948 26240 26976
rect 26068 26908 26096 26948
rect 26234 26936 26240 26948
rect 26292 26936 26298 26988
rect 26329 26979 26387 26985
rect 26329 26945 26341 26979
rect 26375 26976 26387 26979
rect 26510 26976 26516 26988
rect 26375 26948 26516 26976
rect 26375 26945 26387 26948
rect 26329 26939 26387 26945
rect 26510 26936 26516 26948
rect 26568 26976 26574 26988
rect 27522 26976 27528 26988
rect 26568 26948 27528 26976
rect 26568 26936 26574 26948
rect 27522 26936 27528 26948
rect 27580 26936 27586 26988
rect 27617 26979 27675 26985
rect 27617 26945 27629 26979
rect 27663 26976 27675 26979
rect 27706 26976 27712 26988
rect 27663 26948 27712 26976
rect 27663 26945 27675 26948
rect 27617 26939 27675 26945
rect 27706 26936 27712 26948
rect 27764 26936 27770 26988
rect 27801 26979 27859 26985
rect 27801 26945 27813 26979
rect 27847 26976 27859 26979
rect 28353 26979 28411 26985
rect 28353 26976 28365 26979
rect 27847 26948 28365 26976
rect 27847 26945 27859 26948
rect 27801 26939 27859 26945
rect 28353 26945 28365 26948
rect 28399 26945 28411 26979
rect 28353 26939 28411 26945
rect 28718 26936 28724 26988
rect 28776 26976 28782 26988
rect 29181 26979 29239 26985
rect 29181 26976 29193 26979
rect 28776 26948 29193 26976
rect 28776 26936 28782 26948
rect 29181 26945 29193 26948
rect 29227 26945 29239 26979
rect 30374 26976 30380 26988
rect 30335 26948 30380 26976
rect 29181 26939 29239 26945
rect 30374 26936 30380 26948
rect 30432 26936 30438 26988
rect 32309 26979 32367 26985
rect 32309 26976 32321 26979
rect 30576 26948 30788 26976
rect 14660 26880 26096 26908
rect 26145 26911 26203 26917
rect 14553 26843 14611 26849
rect 9732 26812 14504 26840
rect 9732 26800 9738 26812
rect 12526 26772 12532 26784
rect 12487 26744 12532 26772
rect 12526 26732 12532 26744
rect 12584 26732 12590 26784
rect 14476 26772 14504 26812
rect 14553 26809 14565 26843
rect 14599 26809 14611 26843
rect 14553 26803 14611 26809
rect 14660 26772 14688 26880
rect 26145 26877 26157 26911
rect 26191 26908 26203 26911
rect 27433 26911 27491 26917
rect 27433 26908 27445 26911
rect 26191 26880 27445 26908
rect 26191 26877 26203 26880
rect 26145 26871 26203 26877
rect 27433 26877 27445 26880
rect 27479 26908 27491 26911
rect 28258 26908 28264 26920
rect 27479 26880 28264 26908
rect 27479 26877 27491 26880
rect 27433 26871 27491 26877
rect 28258 26868 28264 26880
rect 28316 26868 28322 26920
rect 28810 26868 28816 26920
rect 28868 26908 28874 26920
rect 30576 26908 30604 26948
rect 28868 26880 30604 26908
rect 30653 26911 30711 26917
rect 28868 26868 28874 26880
rect 30653 26877 30665 26911
rect 30699 26877 30711 26911
rect 30760 26908 30788 26948
rect 32048 26948 32321 26976
rect 32048 26908 32076 26948
rect 32309 26945 32321 26948
rect 32355 26976 32367 26979
rect 32858 26976 32864 26988
rect 32355 26948 32864 26976
rect 32355 26945 32367 26948
rect 32309 26939 32367 26945
rect 32858 26936 32864 26948
rect 32916 26936 32922 26988
rect 33137 26979 33195 26985
rect 33137 26945 33149 26979
rect 33183 26976 33195 26979
rect 33226 26976 33232 26988
rect 33183 26948 33232 26976
rect 33183 26945 33195 26948
rect 33137 26939 33195 26945
rect 33226 26936 33232 26948
rect 33284 26936 33290 26988
rect 35250 26936 35256 26988
rect 35308 26976 35314 26988
rect 38010 26976 38016 26988
rect 35308 26948 38016 26976
rect 35308 26936 35314 26948
rect 38010 26936 38016 26948
rect 38068 26936 38074 26988
rect 38102 26936 38108 26988
rect 38160 26976 38166 26988
rect 38381 26979 38439 26985
rect 38381 26976 38393 26979
rect 38160 26948 38205 26976
rect 38304 26948 38393 26976
rect 38160 26936 38166 26948
rect 38304 26920 38332 26948
rect 38381 26945 38393 26948
rect 38427 26945 38439 26979
rect 38488 26976 38516 27016
rect 38562 27004 38568 27056
rect 38620 27044 38626 27056
rect 39301 27047 39359 27053
rect 39301 27044 39313 27047
rect 38620 27016 39313 27044
rect 38620 27004 38626 27016
rect 39301 27013 39313 27016
rect 39347 27013 39359 27047
rect 39301 27007 39359 27013
rect 39485 27047 39543 27053
rect 39485 27013 39497 27047
rect 39531 27044 39543 27047
rect 41386 27044 41414 27084
rect 42518 27072 42524 27084
rect 42576 27072 42582 27124
rect 42705 27115 42763 27121
rect 42705 27081 42717 27115
rect 42751 27112 42763 27115
rect 43438 27112 43444 27124
rect 42751 27084 43444 27112
rect 42751 27081 42763 27084
rect 42705 27075 42763 27081
rect 43438 27072 43444 27084
rect 43496 27072 43502 27124
rect 45278 27072 45284 27124
rect 45336 27112 45342 27124
rect 50798 27112 50804 27124
rect 45336 27084 50804 27112
rect 45336 27072 45342 27084
rect 50798 27072 50804 27084
rect 50856 27072 50862 27124
rect 52730 27112 52736 27124
rect 51046 27084 52736 27112
rect 51046 27044 51074 27084
rect 52730 27072 52736 27084
rect 52788 27072 52794 27124
rect 52822 27072 52828 27124
rect 52880 27112 52886 27124
rect 52917 27115 52975 27121
rect 52917 27112 52929 27115
rect 52880 27084 52929 27112
rect 52880 27072 52886 27084
rect 52917 27081 52929 27084
rect 52963 27081 52975 27115
rect 53653 27115 53711 27121
rect 53653 27112 53665 27115
rect 52917 27075 52975 27081
rect 53116 27084 53665 27112
rect 39531 27016 41414 27044
rect 41524 27016 51074 27044
rect 39531 27013 39543 27016
rect 39485 27007 39543 27013
rect 40037 26979 40095 26985
rect 40037 26976 40049 26979
rect 38488 26948 40049 26976
rect 38381 26939 38439 26945
rect 40037 26945 40049 26948
rect 40083 26945 40095 26979
rect 40037 26939 40095 26945
rect 40313 26979 40371 26985
rect 40313 26945 40325 26979
rect 40359 26976 40371 26979
rect 40770 26976 40776 26988
rect 40359 26948 40776 26976
rect 40359 26945 40371 26948
rect 40313 26939 40371 26945
rect 40770 26936 40776 26948
rect 40828 26936 40834 26988
rect 40865 26979 40923 26985
rect 40865 26945 40877 26979
rect 40911 26976 40923 26979
rect 40954 26976 40960 26988
rect 40911 26948 40960 26976
rect 40911 26945 40923 26948
rect 40865 26939 40923 26945
rect 40954 26936 40960 26948
rect 41012 26936 41018 26988
rect 41046 26936 41052 26988
rect 41104 26976 41110 26988
rect 41414 26980 41420 26988
rect 41386 26976 41420 26980
rect 41104 26948 41420 26976
rect 41104 26936 41110 26948
rect 41414 26936 41420 26948
rect 41472 26936 41478 26988
rect 30760 26880 32076 26908
rect 32125 26911 32183 26917
rect 30653 26871 30711 26877
rect 32125 26877 32137 26911
rect 32171 26908 32183 26911
rect 33410 26908 33416 26920
rect 32171 26880 33416 26908
rect 32171 26877 32183 26880
rect 32125 26871 32183 26877
rect 15654 26800 15660 26852
rect 15712 26840 15718 26852
rect 21266 26840 21272 26852
rect 15712 26812 21272 26840
rect 15712 26800 15718 26812
rect 21266 26800 21272 26812
rect 21324 26800 21330 26852
rect 28166 26840 28172 26852
rect 22066 26812 28028 26840
rect 28127 26812 28172 26840
rect 16850 26772 16856 26784
rect 14476 26744 14688 26772
rect 16811 26744 16856 26772
rect 16850 26732 16856 26744
rect 16908 26732 16914 26784
rect 17126 26732 17132 26784
rect 17184 26772 17190 26784
rect 22066 26772 22094 26812
rect 23934 26772 23940 26784
rect 17184 26744 22094 26772
rect 23895 26744 23940 26772
rect 17184 26732 17190 26744
rect 23934 26732 23940 26744
rect 23992 26732 23998 26784
rect 24026 26732 24032 26784
rect 24084 26772 24090 26784
rect 26418 26772 26424 26784
rect 24084 26744 26424 26772
rect 24084 26732 24090 26744
rect 26418 26732 26424 26744
rect 26476 26732 26482 26784
rect 26513 26775 26571 26781
rect 26513 26741 26525 26775
rect 26559 26772 26571 26775
rect 27430 26772 27436 26784
rect 26559 26744 27436 26772
rect 26559 26741 26571 26744
rect 26513 26735 26571 26741
rect 27430 26732 27436 26744
rect 27488 26732 27494 26784
rect 28000 26772 28028 26812
rect 28166 26800 28172 26812
rect 28224 26800 28230 26852
rect 28997 26843 29055 26849
rect 28997 26809 29009 26843
rect 29043 26840 29055 26843
rect 29914 26840 29920 26852
rect 29043 26812 29920 26840
rect 29043 26809 29055 26812
rect 28997 26803 29055 26809
rect 29914 26800 29920 26812
rect 29972 26800 29978 26852
rect 30006 26800 30012 26852
rect 30064 26840 30070 26852
rect 30668 26840 30696 26871
rect 33410 26868 33416 26880
rect 33468 26868 33474 26920
rect 33980 26880 38240 26908
rect 30064 26812 30696 26840
rect 30064 26800 30070 26812
rect 30742 26800 30748 26852
rect 30800 26840 30806 26852
rect 33980 26840 34008 26880
rect 30800 26812 34008 26840
rect 38212 26840 38240 26880
rect 38286 26868 38292 26920
rect 38344 26868 38350 26920
rect 41524 26908 41552 27016
rect 53116 27009 53144 27084
rect 53653 27081 53665 27084
rect 53699 27081 53711 27115
rect 53653 27075 53711 27081
rect 56137 27115 56195 27121
rect 56137 27081 56149 27115
rect 56183 27112 56195 27115
rect 57054 27112 57060 27124
rect 56183 27084 57060 27112
rect 56183 27081 56195 27084
rect 56137 27075 56195 27081
rect 57054 27072 57060 27084
rect 57112 27072 57118 27124
rect 57974 27072 57980 27124
rect 58032 27112 58038 27124
rect 58805 27115 58863 27121
rect 58805 27112 58817 27115
rect 58032 27084 58817 27112
rect 58032 27072 58038 27084
rect 58805 27081 58817 27084
rect 58851 27081 58863 27115
rect 60642 27112 60648 27124
rect 60603 27084 60648 27112
rect 58805 27075 58863 27081
rect 60642 27072 60648 27084
rect 60700 27072 60706 27124
rect 64325 27115 64383 27121
rect 64325 27081 64337 27115
rect 64371 27081 64383 27115
rect 64325 27075 64383 27081
rect 53101 27003 53159 27009
rect 53190 27004 53196 27056
rect 53248 27044 53254 27056
rect 64340 27044 64368 27075
rect 64874 27072 64880 27124
rect 64932 27112 64938 27124
rect 65429 27115 65487 27121
rect 64932 27084 64977 27112
rect 64932 27072 64938 27084
rect 65429 27081 65441 27115
rect 65475 27112 65487 27115
rect 66438 27112 66444 27124
rect 65475 27084 66444 27112
rect 65475 27081 65487 27084
rect 65429 27075 65487 27081
rect 66438 27072 66444 27084
rect 66496 27072 66502 27124
rect 68833 27115 68891 27121
rect 68833 27081 68845 27115
rect 68879 27112 68891 27115
rect 69382 27112 69388 27124
rect 68879 27084 69388 27112
rect 68879 27081 68891 27084
rect 68833 27075 68891 27081
rect 69382 27072 69388 27084
rect 69440 27072 69446 27124
rect 70121 27115 70179 27121
rect 70121 27081 70133 27115
rect 70167 27112 70179 27115
rect 71498 27112 71504 27124
rect 70167 27084 71504 27112
rect 70167 27081 70179 27084
rect 70121 27075 70179 27081
rect 71498 27072 71504 27084
rect 71556 27072 71562 27124
rect 73154 27072 73160 27124
rect 73212 27112 73218 27124
rect 73341 27115 73399 27121
rect 73341 27112 73353 27115
rect 73212 27084 73353 27112
rect 73212 27072 73218 27084
rect 73341 27081 73353 27084
rect 73387 27081 73399 27115
rect 73341 27075 73399 27081
rect 74629 27115 74687 27121
rect 74629 27081 74641 27115
rect 74675 27112 74687 27115
rect 75086 27112 75092 27124
rect 74675 27084 75092 27112
rect 74675 27081 74687 27084
rect 74629 27075 74687 27081
rect 75086 27072 75092 27084
rect 75144 27072 75150 27124
rect 75454 27112 75460 27124
rect 75415 27084 75460 27112
rect 75454 27072 75460 27084
rect 75512 27072 75518 27124
rect 79689 27115 79747 27121
rect 79689 27081 79701 27115
rect 79735 27112 79747 27115
rect 83826 27112 83832 27124
rect 79735 27084 83832 27112
rect 79735 27081 79747 27084
rect 79689 27075 79747 27081
rect 83826 27072 83832 27084
rect 83884 27072 83890 27124
rect 86310 27112 86316 27124
rect 86271 27084 86316 27112
rect 86310 27072 86316 27084
rect 86368 27072 86374 27124
rect 86865 27115 86923 27121
rect 86865 27081 86877 27115
rect 86911 27112 86923 27115
rect 86954 27112 86960 27124
rect 86911 27084 86960 27112
rect 86911 27081 86923 27084
rect 86865 27075 86923 27081
rect 86954 27072 86960 27084
rect 87012 27072 87018 27124
rect 53248 27016 60872 27044
rect 64340 27016 64874 27044
rect 53248 27004 53254 27016
rect 41690 26936 41696 26988
rect 41748 26976 41754 26988
rect 42889 26979 42947 26985
rect 42889 26976 42901 26979
rect 41748 26948 42901 26976
rect 41748 26936 41754 26948
rect 42889 26945 42901 26948
rect 42935 26976 42947 26979
rect 44174 26976 44180 26988
rect 42935 26948 44180 26976
rect 42935 26945 42947 26948
rect 42889 26939 42947 26945
rect 44174 26936 44180 26948
rect 44232 26936 44238 26988
rect 44726 26976 44732 26988
rect 44687 26948 44732 26976
rect 44726 26936 44732 26948
rect 44784 26936 44790 26988
rect 44818 26936 44824 26988
rect 44876 26976 44882 26988
rect 48774 26976 48780 26988
rect 44876 26948 48780 26976
rect 44876 26936 44882 26948
rect 48774 26936 48780 26948
rect 48832 26936 48838 26988
rect 49694 26936 49700 26988
rect 49752 26976 49758 26988
rect 49881 26979 49939 26985
rect 49881 26976 49893 26979
rect 49752 26948 49893 26976
rect 49752 26936 49758 26948
rect 49881 26945 49893 26948
rect 49927 26945 49939 26979
rect 53101 26969 53113 27003
rect 53147 26969 53159 27003
rect 53101 26963 53159 26969
rect 53837 26979 53895 26985
rect 49881 26939 49939 26945
rect 53837 26945 53849 26979
rect 53883 26976 53895 26979
rect 53926 26976 53932 26988
rect 53883 26948 53932 26976
rect 53883 26945 53895 26948
rect 53837 26939 53895 26945
rect 53926 26936 53932 26948
rect 53984 26936 53990 26988
rect 54202 26976 54208 26988
rect 54163 26948 54208 26976
rect 54202 26936 54208 26948
rect 54260 26936 54266 26988
rect 55490 26936 55496 26988
rect 55548 26976 55554 26988
rect 56321 26979 56379 26985
rect 56321 26976 56333 26979
rect 55548 26948 56333 26976
rect 55548 26936 55554 26948
rect 56321 26945 56333 26948
rect 56367 26945 56379 26979
rect 58434 26976 58440 26988
rect 58395 26948 58440 26976
rect 56321 26939 56379 26945
rect 58434 26936 58440 26948
rect 58492 26936 58498 26988
rect 58986 26976 58992 26988
rect 58947 26948 58992 26976
rect 58986 26936 58992 26948
rect 59044 26936 59050 26988
rect 60844 26985 60872 27016
rect 60829 26979 60887 26985
rect 60829 26945 60841 26979
rect 60875 26945 60887 26979
rect 64506 26976 64512 26988
rect 64467 26948 64512 26976
rect 60829 26939 60887 26945
rect 64506 26936 64512 26948
rect 64564 26936 64570 26988
rect 64846 26976 64874 27016
rect 68462 27004 68468 27056
rect 68520 27044 68526 27056
rect 81526 27044 81532 27056
rect 68520 27016 81532 27044
rect 68520 27004 68526 27016
rect 81526 27004 81532 27016
rect 81584 27004 81590 27056
rect 65061 26979 65119 26985
rect 65061 26976 65073 26979
rect 64846 26948 65073 26976
rect 65061 26945 65073 26948
rect 65107 26945 65119 26979
rect 65610 26976 65616 26988
rect 65571 26948 65616 26976
rect 65061 26939 65119 26945
rect 65610 26936 65616 26948
rect 65668 26936 65674 26988
rect 69017 26979 69075 26985
rect 69017 26945 69029 26979
rect 69063 26976 69075 26979
rect 70118 26976 70124 26988
rect 69063 26948 70124 26976
rect 69063 26945 69075 26948
rect 69017 26939 69075 26945
rect 70118 26936 70124 26948
rect 70176 26976 70182 26988
rect 70305 26979 70363 26985
rect 70305 26976 70317 26979
rect 70176 26948 70317 26976
rect 70176 26936 70182 26948
rect 70305 26945 70317 26948
rect 70351 26945 70363 26979
rect 73522 26976 73528 26988
rect 73483 26948 73528 26976
rect 70305 26939 70363 26945
rect 73522 26936 73528 26948
rect 73580 26936 73586 26988
rect 73890 26936 73896 26988
rect 73948 26976 73954 26988
rect 74813 26979 74871 26985
rect 74813 26976 74825 26979
rect 73948 26948 74825 26976
rect 73948 26936 73954 26948
rect 74813 26945 74825 26948
rect 74859 26945 74871 26979
rect 75638 26976 75644 26988
rect 75599 26948 75644 26976
rect 74813 26939 74871 26945
rect 75638 26936 75644 26948
rect 75696 26936 75702 26988
rect 77389 26979 77447 26985
rect 77389 26976 77401 26979
rect 75932 26948 77401 26976
rect 38488 26880 41552 26908
rect 38488 26840 38516 26880
rect 41782 26868 41788 26920
rect 41840 26908 41846 26920
rect 54294 26908 54300 26920
rect 41840 26880 54300 26908
rect 41840 26868 41846 26880
rect 54294 26868 54300 26880
rect 54352 26868 54358 26920
rect 54478 26908 54484 26920
rect 54439 26880 54484 26908
rect 54478 26868 54484 26880
rect 54536 26868 54542 26920
rect 56962 26868 56968 26920
rect 57020 26908 57026 26920
rect 69198 26908 69204 26920
rect 57020 26880 69204 26908
rect 57020 26868 57026 26880
rect 69198 26868 69204 26880
rect 69256 26908 69262 26920
rect 75932 26908 75960 26948
rect 77389 26945 77401 26948
rect 77435 26945 77447 26979
rect 77389 26939 77447 26945
rect 77573 26979 77631 26985
rect 77573 26945 77585 26979
rect 77619 26976 77631 26979
rect 79873 26979 79931 26985
rect 79873 26976 79885 26979
rect 77619 26948 79885 26976
rect 77619 26945 77631 26948
rect 77573 26939 77631 26945
rect 79873 26945 79885 26948
rect 79919 26945 79931 26979
rect 79873 26939 79931 26945
rect 84378 26936 84384 26988
rect 84436 26976 84442 26988
rect 84657 26979 84715 26985
rect 84657 26976 84669 26979
rect 84436 26948 84669 26976
rect 84436 26936 84442 26948
rect 84657 26945 84669 26948
rect 84703 26945 84715 26979
rect 84657 26939 84715 26945
rect 85114 26936 85120 26988
rect 85172 26976 85178 26988
rect 85209 26979 85267 26985
rect 85209 26976 85221 26979
rect 85172 26948 85221 26976
rect 85172 26936 85178 26948
rect 85209 26945 85221 26948
rect 85255 26945 85267 26979
rect 85209 26939 85267 26945
rect 86497 26979 86555 26985
rect 86497 26945 86509 26979
rect 86543 26945 86555 26979
rect 86497 26939 86555 26945
rect 87049 26979 87107 26985
rect 87049 26945 87061 26979
rect 87095 26976 87107 26979
rect 87230 26976 87236 26988
rect 87095 26948 87236 26976
rect 87095 26945 87107 26948
rect 87049 26939 87107 26945
rect 69256 26880 75960 26908
rect 69256 26868 69262 26880
rect 76742 26868 76748 26920
rect 76800 26908 76806 26920
rect 77205 26911 77263 26917
rect 77205 26908 77217 26911
rect 76800 26880 77217 26908
rect 76800 26868 76806 26880
rect 77205 26877 77217 26880
rect 77251 26877 77263 26911
rect 77205 26871 77263 26877
rect 38212 26812 38516 26840
rect 39853 26843 39911 26849
rect 30800 26800 30806 26812
rect 39853 26809 39865 26843
rect 39899 26840 39911 26843
rect 44818 26840 44824 26852
rect 39899 26812 44824 26840
rect 39899 26809 39911 26812
rect 39853 26803 39911 26809
rect 44818 26800 44824 26812
rect 44876 26800 44882 26852
rect 44913 26843 44971 26849
rect 44913 26809 44925 26843
rect 44959 26840 44971 26843
rect 86512 26840 86540 26939
rect 87230 26936 87236 26948
rect 87288 26936 87294 26988
rect 87414 26908 87420 26920
rect 87375 26880 87420 26908
rect 87414 26868 87420 26880
rect 87472 26868 87478 26920
rect 87693 26911 87751 26917
rect 87693 26877 87705 26911
rect 87739 26877 87751 26911
rect 87693 26871 87751 26877
rect 44959 26812 53144 26840
rect 44959 26809 44971 26812
rect 44913 26803 44971 26809
rect 30466 26772 30472 26784
rect 28000 26744 30472 26772
rect 30466 26732 30472 26744
rect 30524 26732 30530 26784
rect 30650 26732 30656 26784
rect 30708 26772 30714 26784
rect 32493 26775 32551 26781
rect 32493 26772 32505 26775
rect 30708 26744 32505 26772
rect 30708 26732 30714 26744
rect 32493 26741 32505 26744
rect 32539 26741 32551 26775
rect 32858 26772 32864 26784
rect 32771 26744 32864 26772
rect 32493 26735 32551 26741
rect 32858 26732 32864 26744
rect 32916 26772 32922 26784
rect 41046 26772 41052 26784
rect 32916 26744 41052 26772
rect 32916 26732 32922 26744
rect 41046 26732 41052 26744
rect 41104 26732 41110 26784
rect 41414 26732 41420 26784
rect 41472 26772 41478 26784
rect 42610 26772 42616 26784
rect 41472 26744 42616 26772
rect 41472 26732 41478 26744
rect 42610 26732 42616 26744
rect 42668 26732 42674 26784
rect 42702 26732 42708 26784
rect 42760 26772 42766 26784
rect 49326 26772 49332 26784
rect 42760 26744 49332 26772
rect 42760 26732 42766 26744
rect 49326 26732 49332 26744
rect 49384 26732 49390 26784
rect 49697 26775 49755 26781
rect 49697 26741 49709 26775
rect 49743 26772 49755 26775
rect 50338 26772 50344 26784
rect 49743 26744 50344 26772
rect 49743 26741 49755 26744
rect 49697 26735 49755 26741
rect 50338 26732 50344 26744
rect 50396 26732 50402 26784
rect 53116 26772 53144 26812
rect 57946 26812 86540 26840
rect 57946 26772 57974 26812
rect 86586 26800 86592 26852
rect 86644 26840 86650 26852
rect 87708 26840 87736 26871
rect 86644 26812 87736 26840
rect 86644 26800 86650 26812
rect 53116 26744 57974 26772
rect 58253 26775 58311 26781
rect 58253 26741 58265 26775
rect 58299 26772 58311 26775
rect 59630 26772 59636 26784
rect 58299 26744 59636 26772
rect 58299 26741 58311 26744
rect 58253 26735 58311 26741
rect 59630 26732 59636 26744
rect 59688 26732 59694 26784
rect 68554 26732 68560 26784
rect 68612 26772 68618 26784
rect 75089 26775 75147 26781
rect 75089 26772 75101 26775
rect 68612 26744 75101 26772
rect 68612 26732 68618 26744
rect 75089 26741 75101 26744
rect 75135 26772 75147 26775
rect 75638 26772 75644 26784
rect 75135 26744 75644 26772
rect 75135 26741 75147 26744
rect 75089 26735 75147 26741
rect 75638 26732 75644 26744
rect 75696 26732 75702 26784
rect 85390 26772 85396 26784
rect 85351 26744 85396 26772
rect 85390 26732 85396 26744
rect 85448 26732 85454 26784
rect 1104 26682 88872 26704
rect 1104 26630 11924 26682
rect 11976 26630 11988 26682
rect 12040 26630 12052 26682
rect 12104 26630 12116 26682
rect 12168 26630 12180 26682
rect 12232 26630 33872 26682
rect 33924 26630 33936 26682
rect 33988 26630 34000 26682
rect 34052 26630 34064 26682
rect 34116 26630 34128 26682
rect 34180 26630 55820 26682
rect 55872 26630 55884 26682
rect 55936 26630 55948 26682
rect 56000 26630 56012 26682
rect 56064 26630 56076 26682
rect 56128 26630 77768 26682
rect 77820 26630 77832 26682
rect 77884 26630 77896 26682
rect 77948 26630 77960 26682
rect 78012 26630 78024 26682
rect 78076 26630 88872 26682
rect 1104 26608 88872 26630
rect 2222 26528 2228 26580
rect 2280 26568 2286 26580
rect 2869 26571 2927 26577
rect 2869 26568 2881 26571
rect 2280 26540 2881 26568
rect 2280 26528 2286 26540
rect 2869 26537 2881 26540
rect 2915 26537 2927 26571
rect 2869 26531 2927 26537
rect 12526 26528 12532 26580
rect 12584 26568 12590 26580
rect 42702 26568 42708 26580
rect 12584 26540 42708 26568
rect 12584 26528 12590 26540
rect 42702 26528 42708 26540
rect 42760 26528 42766 26580
rect 42794 26528 42800 26580
rect 42852 26568 42858 26580
rect 54754 26568 54760 26580
rect 42852 26540 54760 26568
rect 42852 26528 42858 26540
rect 54754 26528 54760 26540
rect 54812 26528 54818 26580
rect 55674 26528 55680 26580
rect 55732 26568 55738 26580
rect 65058 26568 65064 26580
rect 55732 26540 65064 26568
rect 55732 26528 55738 26540
rect 65058 26528 65064 26540
rect 65116 26568 65122 26580
rect 65610 26568 65616 26580
rect 65116 26540 65616 26568
rect 65116 26528 65122 26540
rect 65610 26528 65616 26540
rect 65668 26528 65674 26580
rect 87417 26571 87475 26577
rect 87417 26537 87429 26571
rect 87463 26568 87475 26571
rect 88242 26568 88248 26580
rect 87463 26540 88248 26568
rect 87463 26537 87475 26540
rect 87417 26531 87475 26537
rect 88242 26528 88248 26540
rect 88300 26528 88306 26580
rect 14458 26460 14464 26512
rect 14516 26500 14522 26512
rect 20070 26500 20076 26512
rect 14516 26472 20076 26500
rect 14516 26460 14522 26472
rect 20070 26460 20076 26472
rect 20128 26460 20134 26512
rect 20438 26460 20444 26512
rect 20496 26500 20502 26512
rect 26694 26500 26700 26512
rect 20496 26472 26556 26500
rect 26655 26472 26700 26500
rect 20496 26460 20502 26472
rect 18230 26392 18236 26444
rect 18288 26432 18294 26444
rect 22002 26432 22008 26444
rect 18288 26404 22008 26432
rect 18288 26392 18294 26404
rect 22002 26392 22008 26404
rect 22060 26392 22066 26444
rect 26528 26432 26556 26472
rect 26694 26460 26700 26472
rect 26752 26460 26758 26512
rect 27246 26500 27252 26512
rect 27207 26472 27252 26500
rect 27246 26460 27252 26472
rect 27304 26460 27310 26512
rect 31754 26500 31760 26512
rect 27356 26472 31760 26500
rect 27356 26432 27384 26472
rect 31754 26460 31760 26472
rect 31812 26460 31818 26512
rect 35342 26460 35348 26512
rect 35400 26500 35406 26512
rect 38286 26500 38292 26512
rect 35400 26472 38292 26500
rect 35400 26460 35406 26472
rect 38286 26460 38292 26472
rect 38344 26500 38350 26512
rect 40678 26500 40684 26512
rect 38344 26472 40684 26500
rect 38344 26460 38350 26472
rect 40678 26460 40684 26472
rect 40736 26460 40742 26512
rect 40954 26500 40960 26512
rect 40915 26472 40960 26500
rect 40954 26460 40960 26472
rect 41012 26460 41018 26512
rect 41046 26460 41052 26512
rect 41104 26500 41110 26512
rect 68554 26500 68560 26512
rect 41104 26472 68560 26500
rect 41104 26460 41110 26472
rect 68554 26460 68560 26472
rect 68612 26460 68618 26512
rect 26528 26404 27384 26432
rect 1394 26364 1400 26376
rect 1355 26336 1400 26364
rect 1394 26324 1400 26336
rect 1452 26324 1458 26376
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26364 1731 26367
rect 1854 26364 1860 26376
rect 1719 26336 1860 26364
rect 1719 26333 1731 26336
rect 1673 26327 1731 26333
rect 1854 26324 1860 26336
rect 1912 26324 1918 26376
rect 3050 26364 3056 26376
rect 3011 26336 3056 26364
rect 3050 26324 3056 26336
rect 3108 26324 3114 26376
rect 3970 26364 3976 26376
rect 3931 26336 3976 26364
rect 3970 26324 3976 26336
rect 4028 26324 4034 26376
rect 16850 26324 16856 26376
rect 16908 26364 16914 26376
rect 25958 26364 25964 26376
rect 16908 26336 25964 26364
rect 16908 26324 16914 26336
rect 25958 26324 25964 26336
rect 26016 26324 26022 26376
rect 26804 26364 26832 26404
rect 27706 26392 27712 26444
rect 27764 26432 27770 26444
rect 27764 26404 29868 26432
rect 27764 26392 27770 26404
rect 26881 26367 26939 26373
rect 26881 26364 26893 26367
rect 26804 26336 26893 26364
rect 26881 26333 26893 26336
rect 26927 26333 26939 26367
rect 27430 26364 27436 26376
rect 27391 26336 27436 26364
rect 26881 26327 26939 26333
rect 27430 26324 27436 26336
rect 27488 26324 27494 26376
rect 27798 26324 27804 26376
rect 27856 26364 27862 26376
rect 29178 26364 29184 26376
rect 27856 26336 29184 26364
rect 27856 26324 27862 26336
rect 29178 26324 29184 26336
rect 29236 26324 29242 26376
rect 29454 26324 29460 26376
rect 29512 26364 29518 26376
rect 29549 26367 29607 26373
rect 29549 26364 29561 26367
rect 29512 26336 29561 26364
rect 29512 26324 29518 26336
rect 29549 26333 29561 26336
rect 29595 26333 29607 26367
rect 29549 26327 29607 26333
rect 29638 26324 29644 26376
rect 29696 26364 29702 26376
rect 29733 26367 29791 26373
rect 29733 26364 29745 26367
rect 29696 26336 29745 26364
rect 29696 26324 29702 26336
rect 29733 26333 29745 26336
rect 29779 26333 29791 26367
rect 29840 26364 29868 26404
rect 35526 26392 35532 26444
rect 35584 26432 35590 26444
rect 39390 26432 39396 26444
rect 35584 26404 39396 26432
rect 35584 26392 35590 26404
rect 39390 26392 39396 26404
rect 39448 26392 39454 26444
rect 40589 26435 40647 26441
rect 40589 26401 40601 26435
rect 40635 26432 40647 26435
rect 43254 26432 43260 26444
rect 40635 26404 43260 26432
rect 40635 26401 40647 26404
rect 40589 26395 40647 26401
rect 43254 26392 43260 26404
rect 43312 26392 43318 26444
rect 44818 26392 44824 26444
rect 44876 26432 44882 26444
rect 58986 26432 58992 26444
rect 44876 26404 58992 26432
rect 44876 26392 44882 26404
rect 58986 26392 58992 26404
rect 59044 26392 59050 26444
rect 68922 26392 68928 26444
rect 68980 26432 68986 26444
rect 82722 26432 82728 26444
rect 68980 26404 82728 26432
rect 68980 26392 68986 26404
rect 82722 26392 82728 26404
rect 82780 26392 82786 26444
rect 85390 26392 85396 26444
rect 85448 26432 85454 26444
rect 85448 26404 87644 26432
rect 85448 26392 85454 26404
rect 30374 26364 30380 26376
rect 29840 26336 30380 26364
rect 29733 26327 29791 26333
rect 30374 26324 30380 26336
rect 30432 26324 30438 26376
rect 30650 26364 30656 26376
rect 30611 26336 30656 26364
rect 30650 26324 30656 26336
rect 30708 26324 30714 26376
rect 31018 26364 31024 26376
rect 30979 26336 31024 26364
rect 31018 26324 31024 26336
rect 31076 26324 31082 26376
rect 31294 26364 31300 26376
rect 31255 26336 31300 26364
rect 31294 26324 31300 26336
rect 31352 26324 31358 26376
rect 38194 26324 38200 26376
rect 38252 26364 38258 26376
rect 40678 26364 40684 26376
rect 38252 26336 40684 26364
rect 38252 26324 38258 26336
rect 40678 26324 40684 26336
rect 40736 26324 40742 26376
rect 40773 26367 40831 26373
rect 40773 26333 40785 26367
rect 40819 26364 40831 26367
rect 40862 26364 40868 26376
rect 40819 26336 40868 26364
rect 40819 26333 40831 26336
rect 40773 26327 40831 26333
rect 40862 26324 40868 26336
rect 40920 26324 40926 26376
rect 42610 26324 42616 26376
rect 42668 26364 42674 26376
rect 45278 26364 45284 26376
rect 42668 26336 45284 26364
rect 42668 26324 42674 26336
rect 45278 26324 45284 26336
rect 45336 26324 45342 26376
rect 45370 26324 45376 26376
rect 45428 26364 45434 26376
rect 55582 26364 55588 26376
rect 45428 26336 55588 26364
rect 45428 26324 45434 26336
rect 55582 26324 55588 26336
rect 55640 26324 55646 26376
rect 70118 26324 70124 26376
rect 70176 26364 70182 26376
rect 85114 26364 85120 26376
rect 70176 26336 85120 26364
rect 70176 26324 70182 26336
rect 85114 26324 85120 26336
rect 85172 26324 85178 26376
rect 87046 26364 87052 26376
rect 87007 26336 87052 26364
rect 87046 26324 87052 26336
rect 87104 26324 87110 26376
rect 87616 26373 87644 26404
rect 87601 26367 87659 26373
rect 87601 26333 87613 26367
rect 87647 26333 87659 26367
rect 87966 26364 87972 26376
rect 87927 26336 87972 26364
rect 87601 26327 87659 26333
rect 87966 26324 87972 26336
rect 88024 26324 88030 26376
rect 13538 26256 13544 26308
rect 13596 26296 13602 26308
rect 20346 26296 20352 26308
rect 13596 26268 20352 26296
rect 13596 26256 13602 26268
rect 20346 26256 20352 26268
rect 20404 26256 20410 26308
rect 23382 26296 23388 26308
rect 20456 26268 23388 26296
rect 3786 26228 3792 26240
rect 3747 26200 3792 26228
rect 3786 26188 3792 26200
rect 3844 26188 3850 26240
rect 19426 26188 19432 26240
rect 19484 26228 19490 26240
rect 20456 26228 20484 26268
rect 23382 26256 23388 26268
rect 23440 26256 23446 26308
rect 23934 26256 23940 26308
rect 23992 26296 23998 26308
rect 26694 26296 26700 26308
rect 23992 26268 26700 26296
rect 23992 26256 23998 26268
rect 26694 26256 26700 26268
rect 26752 26256 26758 26308
rect 29917 26299 29975 26305
rect 29917 26265 29929 26299
rect 29963 26296 29975 26299
rect 58434 26296 58440 26308
rect 29963 26268 31984 26296
rect 29963 26265 29975 26268
rect 29917 26259 29975 26265
rect 19484 26200 20484 26228
rect 19484 26188 19490 26200
rect 25498 26188 25504 26240
rect 25556 26228 25562 26240
rect 30006 26228 30012 26240
rect 25556 26200 30012 26228
rect 25556 26188 25562 26200
rect 30006 26188 30012 26200
rect 30064 26188 30070 26240
rect 30466 26228 30472 26240
rect 30427 26200 30472 26228
rect 30466 26188 30472 26200
rect 30524 26188 30530 26240
rect 31956 26228 31984 26268
rect 38626 26268 58440 26296
rect 38626 26228 38654 26268
rect 58434 26256 58440 26268
rect 58492 26256 58498 26308
rect 88886 26296 88892 26308
rect 86880 26268 87460 26296
rect 31956 26200 38654 26228
rect 40862 26188 40868 26240
rect 40920 26228 40926 26240
rect 42058 26228 42064 26240
rect 40920 26200 42064 26228
rect 40920 26188 40926 26200
rect 42058 26188 42064 26200
rect 42116 26228 42122 26240
rect 46658 26228 46664 26240
rect 42116 26200 46664 26228
rect 42116 26188 42122 26200
rect 46658 26188 46664 26200
rect 46716 26188 46722 26240
rect 86880 26237 86908 26268
rect 86865 26231 86923 26237
rect 86865 26197 86877 26231
rect 86911 26228 86923 26231
rect 87432 26228 87460 26268
rect 87984 26268 88892 26296
rect 87984 26228 88012 26268
rect 88886 26256 88892 26268
rect 88944 26256 88950 26308
rect 88150 26228 88156 26240
rect 86911 26200 86945 26228
rect 87432 26200 88012 26228
rect 88111 26200 88156 26228
rect 86911 26197 86923 26200
rect 86865 26191 86923 26197
rect 88150 26188 88156 26200
rect 88208 26188 88214 26240
rect 1104 26138 88872 26160
rect 1104 26086 22898 26138
rect 22950 26086 22962 26138
rect 23014 26086 23026 26138
rect 23078 26086 23090 26138
rect 23142 26086 23154 26138
rect 23206 26086 44846 26138
rect 44898 26086 44910 26138
rect 44962 26086 44974 26138
rect 45026 26086 45038 26138
rect 45090 26086 45102 26138
rect 45154 26086 66794 26138
rect 66846 26086 66858 26138
rect 66910 26086 66922 26138
rect 66974 26086 66986 26138
rect 67038 26086 67050 26138
rect 67102 26086 88872 26138
rect 1104 26064 88872 26086
rect 1397 26027 1455 26033
rect 1397 25993 1409 26027
rect 1443 26024 1455 26027
rect 1486 26024 1492 26036
rect 1443 25996 1492 26024
rect 1443 25993 1455 25996
rect 1397 25987 1455 25993
rect 1486 25984 1492 25996
rect 1544 25984 1550 26036
rect 2774 26024 2780 26036
rect 2735 25996 2780 26024
rect 2774 25984 2780 25996
rect 2832 25984 2838 26036
rect 26694 25984 26700 26036
rect 26752 26024 26758 26036
rect 32214 26024 32220 26036
rect 26752 25996 32220 26024
rect 26752 25984 26758 25996
rect 32214 25984 32220 25996
rect 32272 25984 32278 26036
rect 43993 26027 44051 26033
rect 43993 25993 44005 26027
rect 44039 26024 44051 26027
rect 44726 26024 44732 26036
rect 44039 25996 44732 26024
rect 44039 25993 44051 25996
rect 43993 25987 44051 25993
rect 44726 25984 44732 25996
rect 44784 25984 44790 26036
rect 86126 25984 86132 26036
rect 86184 26024 86190 26036
rect 86770 26024 86776 26036
rect 86184 25996 86776 26024
rect 86184 25984 86190 25996
rect 86770 25984 86776 25996
rect 86828 25984 86834 26036
rect 87506 26024 87512 26036
rect 87467 25996 87512 26024
rect 87506 25984 87512 25996
rect 87564 25984 87570 26036
rect 87690 25984 87696 26036
rect 87748 26024 87754 26036
rect 88061 26027 88119 26033
rect 88061 26024 88073 26027
rect 87748 25996 88073 26024
rect 87748 25984 87754 25996
rect 88061 25993 88073 25996
rect 88107 25993 88119 26027
rect 88061 25987 88119 25993
rect 27893 25959 27951 25965
rect 27893 25925 27905 25959
rect 27939 25956 27951 25959
rect 88150 25956 88156 25968
rect 27939 25928 88156 25956
rect 27939 25925 27951 25928
rect 27893 25919 27951 25925
rect 1581 25891 1639 25897
rect 1581 25857 1593 25891
rect 1627 25888 1639 25891
rect 2590 25888 2596 25900
rect 1627 25860 2596 25888
rect 1627 25857 1639 25860
rect 1581 25851 1639 25857
rect 2590 25848 2596 25860
rect 2648 25848 2654 25900
rect 2682 25848 2688 25900
rect 2740 25888 2746 25900
rect 2961 25891 3019 25897
rect 2740 25860 2785 25888
rect 2740 25848 2746 25860
rect 2961 25857 2973 25891
rect 3007 25888 3019 25891
rect 3786 25888 3792 25900
rect 3007 25860 3792 25888
rect 3007 25857 3019 25860
rect 2961 25851 3019 25857
rect 3786 25848 3792 25860
rect 3844 25848 3850 25900
rect 27341 25891 27399 25897
rect 27341 25857 27353 25891
rect 27387 25888 27399 25891
rect 27908 25888 27936 25919
rect 88150 25916 88156 25928
rect 88208 25916 88214 25968
rect 27387 25860 27936 25888
rect 43809 25891 43867 25897
rect 27387 25857 27399 25860
rect 27341 25851 27399 25857
rect 43809 25857 43821 25891
rect 43855 25888 43867 25891
rect 44634 25888 44640 25900
rect 43855 25860 44640 25888
rect 43855 25857 43867 25860
rect 43809 25851 43867 25857
rect 44634 25848 44640 25860
rect 44692 25848 44698 25900
rect 86770 25848 86776 25900
rect 86828 25888 86834 25900
rect 87693 25891 87751 25897
rect 87693 25888 87705 25891
rect 86828 25860 87705 25888
rect 86828 25848 86834 25860
rect 87693 25857 87705 25860
rect 87739 25857 87751 25891
rect 87693 25851 87751 25857
rect 88245 25891 88303 25897
rect 88245 25857 88257 25891
rect 88291 25857 88303 25891
rect 88245 25851 88303 25857
rect 2225 25823 2283 25829
rect 2225 25789 2237 25823
rect 2271 25820 2283 25823
rect 2700 25820 2728 25848
rect 2271 25792 2728 25820
rect 2271 25789 2283 25792
rect 2225 25783 2283 25789
rect 26786 25780 26792 25832
rect 26844 25820 26850 25832
rect 35342 25820 35348 25832
rect 26844 25792 35348 25820
rect 26844 25780 26850 25792
rect 35342 25780 35348 25792
rect 35400 25780 35406 25832
rect 43254 25780 43260 25832
rect 43312 25820 43318 25832
rect 43625 25823 43683 25829
rect 43625 25820 43637 25823
rect 43312 25792 43637 25820
rect 43312 25780 43318 25792
rect 43625 25789 43637 25792
rect 43671 25789 43683 25823
rect 88260 25820 88288 25851
rect 43625 25783 43683 25789
rect 87156 25792 88288 25820
rect 658 25712 664 25764
rect 716 25752 722 25764
rect 2501 25755 2559 25761
rect 2501 25752 2513 25755
rect 716 25724 2513 25752
rect 716 25712 722 25724
rect 2501 25721 2513 25724
rect 2547 25721 2559 25755
rect 2501 25715 2559 25721
rect 13078 25712 13084 25764
rect 13136 25752 13142 25764
rect 32858 25752 32864 25764
rect 13136 25724 32864 25752
rect 13136 25712 13142 25724
rect 32858 25712 32864 25724
rect 32916 25712 32922 25764
rect 33686 25712 33692 25764
rect 33744 25752 33750 25764
rect 58526 25752 58532 25764
rect 33744 25724 58532 25752
rect 33744 25712 33750 25724
rect 58526 25712 58532 25724
rect 58584 25712 58590 25764
rect 87156 25696 87184 25792
rect 3142 25644 3148 25696
rect 3200 25684 3206 25696
rect 21082 25684 21088 25696
rect 3200 25656 21088 25684
rect 3200 25644 3206 25656
rect 21082 25644 21088 25656
rect 21140 25644 21146 25696
rect 26602 25644 26608 25696
rect 26660 25684 26666 25696
rect 27433 25687 27491 25693
rect 27433 25684 27445 25687
rect 26660 25656 27445 25684
rect 26660 25644 26666 25656
rect 27433 25653 27445 25656
rect 27479 25653 27491 25687
rect 87138 25684 87144 25696
rect 87099 25656 87144 25684
rect 27433 25647 27491 25653
rect 87138 25644 87144 25656
rect 87196 25644 87202 25696
rect 1104 25594 88872 25616
rect 1104 25542 11924 25594
rect 11976 25542 11988 25594
rect 12040 25542 12052 25594
rect 12104 25542 12116 25594
rect 12168 25542 12180 25594
rect 12232 25542 33872 25594
rect 33924 25542 33936 25594
rect 33988 25542 34000 25594
rect 34052 25542 34064 25594
rect 34116 25542 34128 25594
rect 34180 25542 55820 25594
rect 55872 25542 55884 25594
rect 55936 25542 55948 25594
rect 56000 25542 56012 25594
rect 56064 25542 56076 25594
rect 56128 25542 77768 25594
rect 77820 25542 77832 25594
rect 77884 25542 77896 25594
rect 77948 25542 77960 25594
rect 78012 25542 78024 25594
rect 78076 25542 88872 25594
rect 1104 25520 88872 25542
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 1673 25279 1731 25285
rect 1673 25245 1685 25279
rect 1719 25276 1731 25279
rect 1719 25248 6914 25276
rect 1719 25245 1731 25248
rect 1673 25239 1731 25245
rect 6886 25208 6914 25248
rect 17954 25208 17960 25220
rect 6886 25180 17960 25208
rect 17954 25168 17960 25180
rect 18012 25168 18018 25220
rect 87874 25208 87880 25220
rect 87835 25180 87880 25208
rect 87874 25168 87880 25180
rect 87932 25168 87938 25220
rect 87966 25140 87972 25152
rect 87927 25112 87972 25140
rect 87966 25100 87972 25112
rect 88024 25100 88030 25152
rect 1104 25050 88872 25072
rect 1104 24998 22898 25050
rect 22950 24998 22962 25050
rect 23014 24998 23026 25050
rect 23078 24998 23090 25050
rect 23142 24998 23154 25050
rect 23206 24998 44846 25050
rect 44898 24998 44910 25050
rect 44962 24998 44974 25050
rect 45026 24998 45038 25050
rect 45090 24998 45102 25050
rect 45154 24998 66794 25050
rect 66846 24998 66858 25050
rect 66910 24998 66922 25050
rect 66974 24998 66986 25050
rect 67038 24998 67050 25050
rect 67102 24998 88872 25050
rect 1104 24976 88872 24998
rect 88242 24800 88248 24812
rect 88203 24772 88248 24800
rect 88242 24760 88248 24772
rect 88300 24760 88306 24812
rect 1394 24732 1400 24744
rect 1355 24704 1400 24732
rect 1394 24692 1400 24704
rect 1452 24692 1458 24744
rect 1673 24735 1731 24741
rect 1673 24701 1685 24735
rect 1719 24732 1731 24735
rect 1719 24704 6914 24732
rect 1719 24701 1731 24704
rect 1673 24695 1731 24701
rect 6886 24664 6914 24704
rect 22738 24664 22744 24676
rect 6886 24636 22744 24664
rect 22738 24624 22744 24636
rect 22796 24624 22802 24676
rect 88058 24596 88064 24608
rect 88019 24568 88064 24596
rect 88058 24556 88064 24568
rect 88116 24556 88122 24608
rect 1104 24506 88872 24528
rect 1104 24454 11924 24506
rect 11976 24454 11988 24506
rect 12040 24454 12052 24506
rect 12104 24454 12116 24506
rect 12168 24454 12180 24506
rect 12232 24454 33872 24506
rect 33924 24454 33936 24506
rect 33988 24454 34000 24506
rect 34052 24454 34064 24506
rect 34116 24454 34128 24506
rect 34180 24454 55820 24506
rect 55872 24454 55884 24506
rect 55936 24454 55948 24506
rect 56000 24454 56012 24506
rect 56064 24454 56076 24506
rect 56128 24454 77768 24506
rect 77820 24454 77832 24506
rect 77884 24454 77896 24506
rect 77948 24454 77960 24506
rect 78012 24454 78024 24506
rect 78076 24454 88872 24506
rect 1104 24432 88872 24454
rect 53926 24216 53932 24268
rect 53984 24256 53990 24268
rect 63402 24256 63408 24268
rect 53984 24228 63408 24256
rect 53984 24216 53990 24228
rect 63402 24216 63408 24228
rect 63460 24216 63466 24268
rect 35710 24148 35716 24200
rect 35768 24188 35774 24200
rect 64322 24188 64328 24200
rect 35768 24160 64328 24188
rect 35768 24148 35774 24160
rect 64322 24148 64328 24160
rect 64380 24148 64386 24200
rect 86770 24148 86776 24200
rect 86828 24188 86834 24200
rect 88245 24191 88303 24197
rect 88245 24188 88257 24191
rect 86828 24160 88257 24188
rect 86828 24148 86834 24160
rect 88245 24157 88257 24160
rect 88291 24157 88303 24191
rect 88245 24151 88303 24157
rect 10594 24080 10600 24132
rect 10652 24120 10658 24132
rect 56686 24120 56692 24132
rect 10652 24092 56692 24120
rect 10652 24080 10658 24092
rect 56686 24080 56692 24092
rect 56744 24080 56750 24132
rect 88058 24052 88064 24064
rect 88019 24024 88064 24052
rect 88058 24012 88064 24024
rect 88116 24012 88122 24064
rect 1104 23962 88872 23984
rect 1104 23910 22898 23962
rect 22950 23910 22962 23962
rect 23014 23910 23026 23962
rect 23078 23910 23090 23962
rect 23142 23910 23154 23962
rect 23206 23910 44846 23962
rect 44898 23910 44910 23962
rect 44962 23910 44974 23962
rect 45026 23910 45038 23962
rect 45090 23910 45102 23962
rect 45154 23910 66794 23962
rect 66846 23910 66858 23962
rect 66910 23910 66922 23962
rect 66974 23910 66986 23962
rect 67038 23910 67050 23962
rect 67102 23910 88872 23962
rect 1104 23888 88872 23910
rect 86770 23848 86776 23860
rect 86731 23820 86776 23848
rect 86770 23808 86776 23820
rect 86828 23808 86834 23860
rect 1762 23712 1768 23724
rect 1723 23684 1768 23712
rect 1762 23672 1768 23684
rect 1820 23672 1826 23724
rect 17954 23672 17960 23724
rect 18012 23712 18018 23724
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 18012 23684 21833 23712
rect 18012 23672 18018 23684
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 86957 23715 87015 23721
rect 86957 23712 86969 23715
rect 21821 23675 21879 23681
rect 86420 23684 86969 23712
rect 1949 23579 2007 23585
rect 1949 23545 1961 23579
rect 1995 23576 2007 23579
rect 36814 23576 36820 23588
rect 1995 23548 36820 23576
rect 1995 23545 2007 23548
rect 1949 23539 2007 23545
rect 36814 23536 36820 23548
rect 36872 23536 36878 23588
rect 21913 23511 21971 23517
rect 21913 23477 21925 23511
rect 21959 23508 21971 23511
rect 22278 23508 22284 23520
rect 21959 23480 22284 23508
rect 21959 23477 21971 23480
rect 21913 23471 21971 23477
rect 22278 23468 22284 23480
rect 22336 23468 22342 23520
rect 73982 23468 73988 23520
rect 74040 23508 74046 23520
rect 74442 23508 74448 23520
rect 74040 23480 74448 23508
rect 74040 23468 74046 23480
rect 74442 23468 74448 23480
rect 74500 23508 74506 23520
rect 86420 23517 86448 23684
rect 86957 23681 86969 23684
rect 87003 23681 87015 23715
rect 86957 23675 87015 23681
rect 88245 23715 88303 23721
rect 88245 23681 88257 23715
rect 88291 23681 88303 23715
rect 88245 23675 88303 23681
rect 86494 23604 86500 23656
rect 86552 23644 86558 23656
rect 88260 23644 88288 23675
rect 86552 23616 88288 23644
rect 86552 23604 86558 23616
rect 86405 23511 86463 23517
rect 86405 23508 86417 23511
rect 74500 23480 86417 23508
rect 74500 23468 74506 23480
rect 86405 23477 86417 23480
rect 86451 23477 86463 23511
rect 88058 23508 88064 23520
rect 88019 23480 88064 23508
rect 86405 23471 86463 23477
rect 88058 23468 88064 23480
rect 88116 23468 88122 23520
rect 1104 23418 88872 23440
rect 1104 23366 11924 23418
rect 11976 23366 11988 23418
rect 12040 23366 12052 23418
rect 12104 23366 12116 23418
rect 12168 23366 12180 23418
rect 12232 23366 33872 23418
rect 33924 23366 33936 23418
rect 33988 23366 34000 23418
rect 34052 23366 34064 23418
rect 34116 23366 34128 23418
rect 34180 23366 55820 23418
rect 55872 23366 55884 23418
rect 55936 23366 55948 23418
rect 56000 23366 56012 23418
rect 56064 23366 56076 23418
rect 56128 23366 77768 23418
rect 77820 23366 77832 23418
rect 77884 23366 77896 23418
rect 77948 23366 77960 23418
rect 78012 23366 78024 23418
rect 78076 23366 88872 23418
rect 1104 23344 88872 23366
rect 4798 22924 4804 22976
rect 4856 22964 4862 22976
rect 32306 22964 32312 22976
rect 4856 22936 32312 22964
rect 4856 22924 4862 22936
rect 32306 22924 32312 22936
rect 32364 22924 32370 22976
rect 35066 22924 35072 22976
rect 35124 22964 35130 22976
rect 56318 22964 56324 22976
rect 35124 22936 56324 22964
rect 35124 22924 35130 22936
rect 56318 22924 56324 22936
rect 56376 22924 56382 22976
rect 1104 22874 88872 22896
rect 1104 22822 22898 22874
rect 22950 22822 22962 22874
rect 23014 22822 23026 22874
rect 23078 22822 23090 22874
rect 23142 22822 23154 22874
rect 23206 22822 44846 22874
rect 44898 22822 44910 22874
rect 44962 22822 44974 22874
rect 45026 22822 45038 22874
rect 45090 22822 45102 22874
rect 45154 22822 66794 22874
rect 66846 22822 66858 22874
rect 66910 22822 66922 22874
rect 66974 22822 66986 22874
rect 67038 22822 67050 22874
rect 67102 22822 88872 22874
rect 1104 22800 88872 22822
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 36354 22760 36360 22772
rect 6972 22732 36360 22760
rect 6972 22720 6978 22732
rect 36354 22720 36360 22732
rect 36412 22720 36418 22772
rect 54478 22720 54484 22772
rect 54536 22760 54542 22772
rect 71222 22760 71228 22772
rect 54536 22732 71228 22760
rect 54536 22720 54542 22732
rect 71222 22720 71228 22732
rect 71280 22720 71286 22772
rect 36170 22584 36176 22636
rect 36228 22624 36234 22636
rect 38562 22624 38568 22636
rect 36228 22596 38568 22624
rect 36228 22584 36234 22596
rect 38562 22584 38568 22596
rect 38620 22584 38626 22636
rect 73430 22584 73436 22636
rect 73488 22624 73494 22636
rect 73525 22627 73583 22633
rect 73525 22624 73537 22627
rect 73488 22596 73537 22624
rect 73488 22584 73494 22596
rect 73525 22593 73537 22596
rect 73571 22593 73583 22627
rect 88058 22624 88064 22636
rect 88019 22596 88064 22624
rect 73525 22587 73583 22593
rect 88058 22584 88064 22596
rect 88116 22584 88122 22636
rect 1578 22556 1584 22568
rect 1539 22528 1584 22556
rect 1578 22516 1584 22528
rect 1636 22516 1642 22568
rect 73341 22423 73399 22429
rect 73341 22389 73353 22423
rect 73387 22420 73399 22423
rect 86494 22420 86500 22432
rect 73387 22392 86500 22420
rect 73387 22389 73399 22392
rect 73341 22383 73399 22389
rect 86494 22380 86500 22392
rect 86552 22380 86558 22432
rect 88150 22420 88156 22432
rect 88111 22392 88156 22420
rect 88150 22380 88156 22392
rect 88208 22380 88214 22432
rect 1104 22330 88872 22352
rect 1104 22278 11924 22330
rect 11976 22278 11988 22330
rect 12040 22278 12052 22330
rect 12104 22278 12116 22330
rect 12168 22278 12180 22330
rect 12232 22278 33872 22330
rect 33924 22278 33936 22330
rect 33988 22278 34000 22330
rect 34052 22278 34064 22330
rect 34116 22278 34128 22330
rect 34180 22278 55820 22330
rect 55872 22278 55884 22330
rect 55936 22278 55948 22330
rect 56000 22278 56012 22330
rect 56064 22278 56076 22330
rect 56128 22278 77768 22330
rect 77820 22278 77832 22330
rect 77884 22278 77896 22330
rect 77948 22278 77960 22330
rect 78012 22278 78024 22330
rect 78076 22278 88872 22330
rect 1104 22256 88872 22278
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 22012 1639 22015
rect 16482 22012 16488 22024
rect 1627 21984 16488 22012
rect 1627 21981 1639 21984
rect 1581 21975 1639 21981
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 88245 22015 88303 22021
rect 88245 22012 88257 22015
rect 87708 21984 88257 22012
rect 1394 21876 1400 21888
rect 1355 21848 1400 21876
rect 1394 21836 1400 21848
rect 1452 21836 1458 21888
rect 87598 21836 87604 21888
rect 87656 21876 87662 21888
rect 87708 21885 87736 21984
rect 88245 21981 88257 21984
rect 88291 21981 88303 22015
rect 88245 21975 88303 21981
rect 87693 21879 87751 21885
rect 87693 21876 87705 21879
rect 87656 21848 87705 21876
rect 87656 21836 87662 21848
rect 87693 21845 87705 21848
rect 87739 21845 87751 21879
rect 88058 21876 88064 21888
rect 88019 21848 88064 21876
rect 87693 21839 87751 21845
rect 88058 21836 88064 21848
rect 88116 21836 88122 21888
rect 1104 21786 88872 21808
rect 1104 21734 22898 21786
rect 22950 21734 22962 21786
rect 23014 21734 23026 21786
rect 23078 21734 23090 21786
rect 23142 21734 23154 21786
rect 23206 21734 44846 21786
rect 44898 21734 44910 21786
rect 44962 21734 44974 21786
rect 45026 21734 45038 21786
rect 45090 21734 45102 21786
rect 45154 21734 66794 21786
rect 66846 21734 66858 21786
rect 66910 21734 66922 21786
rect 66974 21734 66986 21786
rect 67038 21734 67050 21786
rect 67102 21734 88872 21786
rect 1104 21712 88872 21734
rect 3970 21632 3976 21684
rect 4028 21672 4034 21684
rect 4157 21675 4215 21681
rect 4157 21672 4169 21675
rect 4028 21644 4169 21672
rect 4028 21632 4034 21644
rect 4157 21641 4169 21644
rect 4203 21641 4215 21675
rect 4157 21635 4215 21641
rect 1394 21536 1400 21548
rect 1355 21508 1400 21536
rect 1394 21496 1400 21508
rect 1452 21496 1458 21548
rect 3970 21536 3976 21548
rect 3931 21508 3976 21536
rect 3970 21496 3976 21508
rect 4028 21496 4034 21548
rect 88245 21539 88303 21545
rect 88245 21536 88257 21539
rect 87708 21508 88257 21536
rect 3789 21471 3847 21477
rect 3789 21437 3801 21471
rect 3835 21468 3847 21471
rect 4798 21468 4804 21480
rect 3835 21440 4804 21468
rect 3835 21437 3847 21440
rect 3789 21431 3847 21437
rect 4798 21428 4804 21440
rect 4856 21428 4862 21480
rect 2590 21360 2596 21412
rect 2648 21400 2654 21412
rect 19886 21400 19892 21412
rect 2648 21372 19892 21400
rect 2648 21360 2654 21372
rect 19886 21360 19892 21372
rect 19944 21360 19950 21412
rect 43990 21360 43996 21412
rect 44048 21400 44054 21412
rect 63218 21400 63224 21412
rect 44048 21372 63224 21400
rect 44048 21360 44054 21372
rect 63218 21360 63224 21372
rect 63276 21360 63282 21412
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 87506 21292 87512 21344
rect 87564 21332 87570 21344
rect 87708 21341 87736 21508
rect 88245 21505 88257 21508
rect 88291 21505 88303 21539
rect 88245 21499 88303 21505
rect 87693 21335 87751 21341
rect 87693 21332 87705 21335
rect 87564 21304 87705 21332
rect 87564 21292 87570 21304
rect 87693 21301 87705 21304
rect 87739 21301 87751 21335
rect 88058 21332 88064 21344
rect 88019 21304 88064 21332
rect 87693 21295 87751 21301
rect 88058 21292 88064 21304
rect 88116 21292 88122 21344
rect 1104 21242 88872 21264
rect 1104 21190 11924 21242
rect 11976 21190 11988 21242
rect 12040 21190 12052 21242
rect 12104 21190 12116 21242
rect 12168 21190 12180 21242
rect 12232 21190 33872 21242
rect 33924 21190 33936 21242
rect 33988 21190 34000 21242
rect 34052 21190 34064 21242
rect 34116 21190 34128 21242
rect 34180 21190 55820 21242
rect 55872 21190 55884 21242
rect 55936 21190 55948 21242
rect 56000 21190 56012 21242
rect 56064 21190 56076 21242
rect 56128 21190 77768 21242
rect 77820 21190 77832 21242
rect 77884 21190 77896 21242
rect 77948 21190 77960 21242
rect 78012 21190 78024 21242
rect 78076 21190 88872 21242
rect 1104 21168 88872 21190
rect 1578 21088 1584 21140
rect 1636 21128 1642 21140
rect 57054 21128 57060 21140
rect 1636 21100 57060 21128
rect 1636 21088 1642 21100
rect 57054 21088 57060 21100
rect 57112 21088 57118 21140
rect 84838 20952 84844 21004
rect 84896 20992 84902 21004
rect 87693 20995 87751 21001
rect 87693 20992 87705 20995
rect 84896 20964 87705 20992
rect 84896 20952 84902 20964
rect 87693 20961 87705 20964
rect 87739 20961 87751 20995
rect 87693 20955 87751 20961
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 87414 20924 87420 20936
rect 1627 20896 1992 20924
rect 87375 20896 87420 20924
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 1964 20800 1992 20896
rect 87414 20884 87420 20896
rect 87472 20884 87478 20936
rect 1394 20788 1400 20800
rect 1355 20760 1400 20788
rect 1394 20748 1400 20760
rect 1452 20748 1458 20800
rect 1946 20788 1952 20800
rect 1907 20760 1952 20788
rect 1946 20748 1952 20760
rect 2004 20748 2010 20800
rect 36814 20748 36820 20800
rect 36872 20788 36878 20800
rect 37734 20788 37740 20800
rect 36872 20760 37740 20788
rect 36872 20748 36878 20760
rect 37734 20748 37740 20760
rect 37792 20748 37798 20800
rect 1104 20698 88872 20720
rect 1104 20646 22898 20698
rect 22950 20646 22962 20698
rect 23014 20646 23026 20698
rect 23078 20646 23090 20698
rect 23142 20646 23154 20698
rect 23206 20646 44846 20698
rect 44898 20646 44910 20698
rect 44962 20646 44974 20698
rect 45026 20646 45038 20698
rect 45090 20646 45102 20698
rect 45154 20646 66794 20698
rect 66846 20646 66858 20698
rect 66910 20646 66922 20698
rect 66974 20646 66986 20698
rect 67038 20646 67050 20698
rect 67102 20646 88872 20698
rect 1104 20624 88872 20646
rect 22002 20544 22008 20596
rect 22060 20584 22066 20596
rect 22189 20587 22247 20593
rect 22189 20584 22201 20587
rect 22060 20556 22201 20584
rect 22060 20544 22066 20556
rect 22189 20553 22201 20556
rect 22235 20553 22247 20587
rect 22189 20547 22247 20553
rect 22462 20476 22468 20528
rect 22520 20516 22526 20528
rect 22557 20519 22615 20525
rect 22557 20516 22569 20519
rect 22520 20488 22569 20516
rect 22520 20476 22526 20488
rect 22557 20485 22569 20488
rect 22603 20485 22615 20519
rect 22557 20479 22615 20485
rect 25866 20476 25872 20528
rect 25924 20516 25930 20528
rect 30285 20519 30343 20525
rect 30285 20516 30297 20519
rect 25924 20488 30297 20516
rect 25924 20476 25930 20488
rect 30285 20485 30297 20488
rect 30331 20485 30343 20519
rect 30285 20479 30343 20485
rect 22373 20451 22431 20457
rect 22373 20417 22385 20451
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 22649 20451 22707 20457
rect 22649 20417 22661 20451
rect 22695 20448 22707 20451
rect 23750 20448 23756 20460
rect 22695 20420 23756 20448
rect 22695 20417 22707 20420
rect 22649 20411 22707 20417
rect 22388 20380 22416 20411
rect 23750 20408 23756 20420
rect 23808 20408 23814 20460
rect 30101 20451 30159 20457
rect 30101 20448 30113 20451
rect 24780 20420 30113 20448
rect 24780 20392 24808 20420
rect 30101 20417 30113 20420
rect 30147 20417 30159 20451
rect 30101 20411 30159 20417
rect 30377 20451 30435 20457
rect 30377 20417 30389 20451
rect 30423 20448 30435 20451
rect 30926 20448 30932 20460
rect 30423 20420 30932 20448
rect 30423 20417 30435 20420
rect 30377 20411 30435 20417
rect 30926 20408 30932 20420
rect 30984 20408 30990 20460
rect 24762 20380 24768 20392
rect 22388 20352 24768 20380
rect 24762 20340 24768 20352
rect 24820 20340 24826 20392
rect 29917 20247 29975 20253
rect 29917 20213 29929 20247
rect 29963 20244 29975 20247
rect 88242 20244 88248 20256
rect 29963 20216 88248 20244
rect 29963 20213 29975 20216
rect 29917 20207 29975 20213
rect 88242 20204 88248 20216
rect 88300 20204 88306 20256
rect 1104 20154 88872 20176
rect 1104 20102 11924 20154
rect 11976 20102 11988 20154
rect 12040 20102 12052 20154
rect 12104 20102 12116 20154
rect 12168 20102 12180 20154
rect 12232 20102 33872 20154
rect 33924 20102 33936 20154
rect 33988 20102 34000 20154
rect 34052 20102 34064 20154
rect 34116 20102 34128 20154
rect 34180 20102 55820 20154
rect 55872 20102 55884 20154
rect 55936 20102 55948 20154
rect 56000 20102 56012 20154
rect 56064 20102 56076 20154
rect 56128 20102 77768 20154
rect 77820 20102 77832 20154
rect 77884 20102 77896 20154
rect 77948 20102 77960 20154
rect 78012 20102 78024 20154
rect 78076 20102 88872 20154
rect 1104 20080 88872 20102
rect 57146 20000 57152 20052
rect 57204 20040 57210 20052
rect 59262 20040 59268 20052
rect 57204 20012 59268 20040
rect 57204 20000 57210 20012
rect 59262 20000 59268 20012
rect 59320 20040 59326 20052
rect 88150 20040 88156 20052
rect 59320 20012 88156 20040
rect 59320 20000 59326 20012
rect 88150 20000 88156 20012
rect 88208 20000 88214 20052
rect 38378 19932 38384 19984
rect 38436 19972 38442 19984
rect 83734 19972 83740 19984
rect 38436 19944 83740 19972
rect 38436 19932 38442 19944
rect 83734 19932 83740 19944
rect 83792 19932 83798 19984
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 1670 19836 1676 19848
rect 1631 19808 1676 19836
rect 1670 19796 1676 19808
rect 1728 19796 1734 19848
rect 88245 19839 88303 19845
rect 88245 19836 88257 19839
rect 87708 19808 88257 19836
rect 87708 19712 87736 19808
rect 88245 19805 88257 19808
rect 88291 19805 88303 19839
rect 88245 19799 88303 19805
rect 87690 19700 87696 19712
rect 87651 19672 87696 19700
rect 87690 19660 87696 19672
rect 87748 19660 87754 19712
rect 88058 19700 88064 19712
rect 88019 19672 88064 19700
rect 88058 19660 88064 19672
rect 88116 19660 88122 19712
rect 1104 19610 88872 19632
rect 1104 19558 22898 19610
rect 22950 19558 22962 19610
rect 23014 19558 23026 19610
rect 23078 19558 23090 19610
rect 23142 19558 23154 19610
rect 23206 19558 44846 19610
rect 44898 19558 44910 19610
rect 44962 19558 44974 19610
rect 45026 19558 45038 19610
rect 45090 19558 45102 19610
rect 45154 19558 66794 19610
rect 66846 19558 66858 19610
rect 66910 19558 66922 19610
rect 66974 19558 66986 19610
rect 67038 19558 67050 19610
rect 67102 19558 88872 19610
rect 1104 19536 88872 19558
rect 63862 19456 63868 19508
rect 63920 19496 63926 19508
rect 87690 19496 87696 19508
rect 63920 19468 87696 19496
rect 63920 19456 63926 19468
rect 87690 19456 87696 19468
rect 87748 19456 87754 19508
rect 25866 19428 25872 19440
rect 24964 19400 25872 19428
rect 24964 19372 24992 19400
rect 25866 19388 25872 19400
rect 25924 19428 25930 19440
rect 26237 19431 26295 19437
rect 26237 19428 26249 19431
rect 25924 19400 26249 19428
rect 25924 19388 25930 19400
rect 26237 19397 26249 19400
rect 26283 19397 26295 19431
rect 27982 19428 27988 19440
rect 26237 19391 26295 19397
rect 26344 19400 27988 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 22462 19320 22468 19372
rect 22520 19360 22526 19372
rect 24946 19360 24952 19372
rect 22520 19332 24952 19360
rect 22520 19320 22526 19332
rect 24946 19320 24952 19332
rect 25004 19320 25010 19372
rect 26344 19369 26372 19400
rect 27982 19388 27988 19400
rect 28040 19388 28046 19440
rect 26053 19363 26111 19369
rect 26053 19329 26065 19363
rect 26099 19360 26111 19363
rect 26329 19363 26387 19369
rect 26099 19332 26280 19360
rect 26099 19329 26111 19332
rect 26053 19323 26111 19329
rect 26252 19292 26280 19332
rect 26329 19329 26341 19363
rect 26375 19329 26387 19363
rect 31386 19360 31392 19372
rect 26329 19323 26387 19329
rect 26436 19332 31392 19360
rect 26436 19292 26464 19332
rect 31386 19320 31392 19332
rect 31444 19360 31450 19372
rect 38102 19360 38108 19372
rect 31444 19332 38108 19360
rect 31444 19320 31450 19332
rect 38102 19320 38108 19332
rect 38160 19320 38166 19372
rect 56502 19360 56508 19372
rect 56463 19332 56508 19360
rect 56502 19320 56508 19332
rect 56560 19320 56566 19372
rect 56594 19320 56600 19372
rect 56652 19360 56658 19372
rect 56689 19363 56747 19369
rect 56689 19360 56701 19363
rect 56652 19332 56701 19360
rect 56652 19320 56658 19332
rect 56689 19329 56701 19332
rect 56735 19329 56747 19363
rect 56689 19323 56747 19329
rect 56781 19363 56839 19369
rect 56781 19329 56793 19363
rect 56827 19360 56839 19363
rect 57146 19360 57152 19372
rect 56827 19332 57152 19360
rect 56827 19329 56839 19332
rect 56781 19323 56839 19329
rect 56318 19292 56324 19304
rect 26252 19264 26464 19292
rect 56279 19264 56324 19292
rect 56318 19252 56324 19264
rect 56376 19252 56382 19304
rect 1949 19227 2007 19233
rect 1949 19193 1961 19227
rect 1995 19224 2007 19227
rect 2590 19224 2596 19236
rect 1995 19196 2596 19224
rect 1995 19193 2007 19196
rect 1949 19187 2007 19193
rect 2590 19184 2596 19196
rect 2648 19184 2654 19236
rect 27798 19184 27804 19236
rect 27856 19224 27862 19236
rect 28074 19224 28080 19236
rect 27856 19196 28080 19224
rect 27856 19184 27862 19196
rect 28074 19184 28080 19196
rect 28132 19184 28138 19236
rect 55677 19227 55735 19233
rect 55677 19193 55689 19227
rect 55723 19224 55735 19227
rect 56045 19227 56103 19233
rect 56045 19224 56057 19227
rect 55723 19196 56057 19224
rect 55723 19193 55735 19196
rect 55677 19187 55735 19193
rect 56045 19193 56057 19196
rect 56091 19224 56103 19227
rect 56796 19224 56824 19323
rect 57146 19320 57152 19332
rect 57204 19320 57210 19372
rect 64966 19320 64972 19372
rect 65024 19360 65030 19372
rect 88245 19363 88303 19369
rect 88245 19360 88257 19363
rect 65024 19332 88257 19360
rect 65024 19320 65030 19332
rect 88245 19329 88257 19332
rect 88291 19329 88303 19363
rect 88245 19323 88303 19329
rect 56091 19196 56824 19224
rect 56091 19193 56103 19196
rect 56045 19187 56103 19193
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 25869 19159 25927 19165
rect 25869 19156 25881 19159
rect 4212 19128 25881 19156
rect 4212 19116 4218 19128
rect 25869 19125 25881 19128
rect 25915 19125 25927 19159
rect 25869 19119 25927 19125
rect 27890 19116 27896 19168
rect 27948 19156 27954 19168
rect 28258 19156 28264 19168
rect 27948 19128 28264 19156
rect 27948 19116 27954 19128
rect 28258 19116 28264 19128
rect 28316 19116 28322 19168
rect 57146 19156 57152 19168
rect 57107 19128 57152 19156
rect 57146 19116 57152 19128
rect 57204 19116 57210 19168
rect 88058 19156 88064 19168
rect 88019 19128 88064 19156
rect 88058 19116 88064 19128
rect 88116 19116 88122 19168
rect 1104 19066 88872 19088
rect 1104 19014 11924 19066
rect 11976 19014 11988 19066
rect 12040 19014 12052 19066
rect 12104 19014 12116 19066
rect 12168 19014 12180 19066
rect 12232 19014 33872 19066
rect 33924 19014 33936 19066
rect 33988 19014 34000 19066
rect 34052 19014 34064 19066
rect 34116 19014 34128 19066
rect 34180 19014 55820 19066
rect 55872 19014 55884 19066
rect 55936 19014 55948 19066
rect 56000 19014 56012 19066
rect 56064 19014 56076 19066
rect 56128 19014 77768 19066
rect 77820 19014 77832 19066
rect 77884 19014 77896 19066
rect 77948 19014 77960 19066
rect 78012 19014 78024 19066
rect 78076 19014 88872 19066
rect 1104 18992 88872 19014
rect 24578 18952 24584 18964
rect 24539 18924 24584 18952
rect 24578 18912 24584 18924
rect 24636 18912 24642 18964
rect 26234 18912 26240 18964
rect 26292 18952 26298 18964
rect 27062 18952 27068 18964
rect 26292 18924 27068 18952
rect 26292 18912 26298 18924
rect 27062 18912 27068 18924
rect 27120 18952 27126 18964
rect 33686 18952 33692 18964
rect 27120 18924 33692 18952
rect 27120 18912 27126 18924
rect 33686 18912 33692 18924
rect 33744 18952 33750 18964
rect 34514 18952 34520 18964
rect 33744 18924 34520 18952
rect 33744 18912 33750 18924
rect 34514 18912 34520 18924
rect 34572 18912 34578 18964
rect 56686 18952 56692 18964
rect 56647 18924 56692 18952
rect 56686 18912 56692 18924
rect 56744 18912 56750 18964
rect 34330 18884 34336 18896
rect 25056 18856 34336 18884
rect 24486 18776 24492 18828
rect 24544 18816 24550 18828
rect 25056 18816 25084 18856
rect 34330 18844 34336 18856
rect 34388 18844 34394 18896
rect 57698 18844 57704 18896
rect 57756 18884 57762 18896
rect 70670 18884 70676 18896
rect 57756 18856 70676 18884
rect 57756 18844 57762 18856
rect 70670 18844 70676 18856
rect 70728 18844 70734 18896
rect 24544 18788 25084 18816
rect 24544 18776 24550 18788
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 1949 18751 2007 18757
rect 1949 18748 1961 18751
rect 1627 18720 1961 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 1949 18717 1961 18720
rect 1995 18748 2007 18751
rect 1995 18720 6914 18748
rect 1995 18717 2007 18720
rect 1949 18711 2007 18717
rect 6886 18680 6914 18720
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 24762 18748 24768 18760
rect 22060 18720 24768 18748
rect 22060 18708 22066 18720
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 24946 18748 24952 18760
rect 24907 18720 24952 18748
rect 24946 18708 24952 18720
rect 25004 18708 25010 18760
rect 25056 18757 25084 18788
rect 27798 18776 27804 18828
rect 27856 18816 27862 18828
rect 28077 18819 28135 18825
rect 28077 18816 28089 18819
rect 27856 18788 28089 18816
rect 27856 18776 27862 18788
rect 28077 18785 28089 18788
rect 28123 18785 28135 18819
rect 28077 18779 28135 18785
rect 28261 18819 28319 18825
rect 28261 18785 28273 18819
rect 28307 18785 28319 18819
rect 28261 18779 28319 18785
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18717 25099 18751
rect 25041 18711 25099 18717
rect 27706 18708 27712 18760
rect 27764 18748 27770 18760
rect 28276 18748 28304 18779
rect 48222 18776 48228 18828
rect 48280 18816 48286 18828
rect 48280 18788 60734 18816
rect 48280 18776 48286 18788
rect 27764 18720 28304 18748
rect 27764 18708 27770 18720
rect 35986 18708 35992 18760
rect 36044 18748 36050 18760
rect 36173 18751 36231 18757
rect 36173 18748 36185 18751
rect 36044 18720 36185 18748
rect 36044 18708 36050 18720
rect 36173 18717 36185 18720
rect 36219 18717 36231 18751
rect 36173 18711 36231 18717
rect 47765 18751 47823 18757
rect 47765 18717 47777 18751
rect 47811 18748 47823 18751
rect 48038 18748 48044 18760
rect 47811 18720 48044 18748
rect 47811 18717 47823 18720
rect 47765 18711 47823 18717
rect 48038 18708 48044 18720
rect 48096 18708 48102 18760
rect 55950 18708 55956 18760
rect 56008 18748 56014 18760
rect 56502 18748 56508 18760
rect 56008 18720 56508 18748
rect 56008 18708 56014 18720
rect 56502 18708 56508 18720
rect 56560 18748 56566 18760
rect 56873 18751 56931 18757
rect 56873 18748 56885 18751
rect 56560 18720 56885 18748
rect 56560 18708 56566 18720
rect 56873 18717 56885 18720
rect 56919 18748 56931 18751
rect 56962 18748 56968 18760
rect 56919 18720 56968 18748
rect 56919 18717 56931 18720
rect 56873 18711 56931 18717
rect 56962 18708 56968 18720
rect 57020 18708 57026 18760
rect 60706 18748 60734 18788
rect 73522 18748 73528 18760
rect 60706 18720 73528 18748
rect 73522 18708 73528 18720
rect 73580 18708 73586 18760
rect 88242 18748 88248 18760
rect 88203 18720 88248 18748
rect 88242 18708 88248 18720
rect 88300 18708 88306 18760
rect 6886 18652 39068 18680
rect 1394 18612 1400 18624
rect 1355 18584 1400 18612
rect 1394 18572 1400 18584
rect 1452 18572 1458 18624
rect 27617 18615 27675 18621
rect 27617 18581 27629 18615
rect 27663 18612 27675 18615
rect 27890 18612 27896 18624
rect 27663 18584 27896 18612
rect 27663 18581 27675 18584
rect 27617 18575 27675 18581
rect 27890 18572 27896 18584
rect 27948 18572 27954 18624
rect 27985 18615 28043 18621
rect 27985 18581 27997 18615
rect 28031 18612 28043 18615
rect 28258 18612 28264 18624
rect 28031 18584 28264 18612
rect 28031 18581 28043 18584
rect 27985 18575 28043 18581
rect 28258 18572 28264 18584
rect 28316 18572 28322 18624
rect 35710 18572 35716 18624
rect 35768 18612 35774 18624
rect 35989 18615 36047 18621
rect 35989 18612 36001 18615
rect 35768 18584 36001 18612
rect 35768 18572 35774 18584
rect 35989 18581 36001 18584
rect 36035 18581 36047 18615
rect 39040 18612 39068 18652
rect 39114 18640 39120 18692
rect 39172 18680 39178 18692
rect 50154 18680 50160 18692
rect 39172 18652 50160 18680
rect 39172 18640 39178 18652
rect 50154 18640 50160 18652
rect 50212 18640 50218 18692
rect 57149 18683 57207 18689
rect 57149 18649 57161 18683
rect 57195 18680 57207 18683
rect 59170 18680 59176 18692
rect 57195 18652 59176 18680
rect 57195 18649 57207 18652
rect 57149 18643 57207 18649
rect 59170 18640 59176 18652
rect 59228 18680 59234 18692
rect 59228 18652 60734 18680
rect 59228 18640 59234 18652
rect 41230 18612 41236 18624
rect 39040 18584 41236 18612
rect 35989 18575 36047 18581
rect 41230 18572 41236 18584
rect 41288 18572 41294 18624
rect 47581 18615 47639 18621
rect 47581 18581 47593 18615
rect 47627 18612 47639 18615
rect 47670 18612 47676 18624
rect 47627 18584 47676 18612
rect 47627 18581 47639 18584
rect 47581 18575 47639 18581
rect 47670 18572 47676 18584
rect 47728 18572 47734 18624
rect 56226 18572 56232 18624
rect 56284 18612 56290 18624
rect 56594 18612 56600 18624
rect 56284 18584 56600 18612
rect 56284 18572 56290 18584
rect 56594 18572 56600 18584
rect 56652 18612 56658 18624
rect 57057 18615 57115 18621
rect 57057 18612 57069 18615
rect 56652 18584 57069 18612
rect 56652 18572 56658 18584
rect 57057 18581 57069 18584
rect 57103 18581 57115 18615
rect 60706 18612 60734 18652
rect 68002 18640 68008 18692
rect 68060 18680 68066 18692
rect 71958 18680 71964 18692
rect 68060 18652 71964 18680
rect 68060 18640 68066 18652
rect 71958 18640 71964 18652
rect 72016 18640 72022 18692
rect 78950 18612 78956 18624
rect 60706 18584 78956 18612
rect 57057 18575 57115 18581
rect 78950 18572 78956 18584
rect 79008 18572 79014 18624
rect 88058 18612 88064 18624
rect 88019 18584 88064 18612
rect 88058 18572 88064 18584
rect 88116 18572 88122 18624
rect 1104 18522 88872 18544
rect 1104 18470 22898 18522
rect 22950 18470 22962 18522
rect 23014 18470 23026 18522
rect 23078 18470 23090 18522
rect 23142 18470 23154 18522
rect 23206 18470 44846 18522
rect 44898 18470 44910 18522
rect 44962 18470 44974 18522
rect 45026 18470 45038 18522
rect 45090 18470 45102 18522
rect 45154 18470 66794 18522
rect 66846 18470 66858 18522
rect 66910 18470 66922 18522
rect 66974 18470 66986 18522
rect 67038 18470 67050 18522
rect 67102 18470 88872 18522
rect 1104 18448 88872 18470
rect 25958 18368 25964 18420
rect 26016 18408 26022 18420
rect 26145 18411 26203 18417
rect 26145 18408 26157 18411
rect 26016 18380 26157 18408
rect 26016 18368 26022 18380
rect 26145 18377 26157 18380
rect 26191 18377 26203 18411
rect 26145 18371 26203 18377
rect 27985 18411 28043 18417
rect 27985 18377 27997 18411
rect 28031 18377 28043 18411
rect 27985 18371 28043 18377
rect 28445 18411 28503 18417
rect 28445 18377 28457 18411
rect 28491 18408 28503 18411
rect 28534 18408 28540 18420
rect 28491 18380 28540 18408
rect 28491 18377 28503 18380
rect 28445 18371 28503 18377
rect 1854 18300 1860 18352
rect 1912 18340 1918 18352
rect 23845 18343 23903 18349
rect 23845 18340 23857 18343
rect 1912 18312 23857 18340
rect 1912 18300 1918 18312
rect 23845 18309 23857 18312
rect 23891 18340 23903 18343
rect 24673 18343 24731 18349
rect 24673 18340 24685 18343
rect 23891 18312 24685 18340
rect 23891 18309 23903 18312
rect 23845 18303 23903 18309
rect 24673 18309 24685 18312
rect 24719 18309 24731 18343
rect 26970 18340 26976 18352
rect 24673 18303 24731 18309
rect 24780 18312 26976 18340
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 12342 18272 12348 18284
rect 1627 18244 12348 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 20806 18232 20812 18284
rect 20864 18272 20870 18284
rect 23750 18272 23756 18284
rect 20864 18244 23756 18272
rect 20864 18232 20870 18244
rect 23750 18232 23756 18244
rect 23808 18272 23814 18284
rect 24581 18275 24639 18281
rect 24581 18272 24593 18275
rect 23808 18244 24593 18272
rect 23808 18232 23814 18244
rect 24581 18241 24593 18244
rect 24627 18272 24639 18275
rect 24780 18272 24808 18312
rect 26970 18300 26976 18312
rect 27028 18300 27034 18352
rect 24627 18244 24808 18272
rect 26053 18275 26111 18281
rect 24627 18241 24639 18244
rect 24581 18235 24639 18241
rect 26053 18241 26065 18275
rect 26099 18272 26111 18275
rect 27430 18272 27436 18284
rect 26099 18244 27436 18272
rect 26099 18241 26111 18244
rect 26053 18235 26111 18241
rect 27430 18232 27436 18244
rect 27488 18232 27494 18284
rect 27617 18275 27675 18281
rect 27617 18241 27629 18275
rect 27663 18272 27675 18275
rect 28000 18272 28028 18371
rect 28534 18368 28540 18380
rect 28592 18368 28598 18420
rect 33965 18411 34023 18417
rect 33965 18377 33977 18411
rect 34011 18377 34023 18411
rect 35986 18408 35992 18420
rect 35947 18380 35992 18408
rect 33965 18371 34023 18377
rect 27663 18244 28028 18272
rect 27663 18241 27675 18244
rect 27617 18235 27675 18241
rect 28074 18232 28080 18284
rect 28132 18272 28138 18284
rect 28350 18272 28356 18284
rect 28132 18244 28356 18272
rect 28132 18232 28138 18244
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 29273 18275 29331 18281
rect 29273 18272 29285 18275
rect 28460 18244 29285 18272
rect 24765 18207 24823 18213
rect 24765 18173 24777 18207
rect 24811 18204 24823 18207
rect 26234 18204 26240 18216
rect 24811 18176 26240 18204
rect 24811 18173 24823 18176
rect 24765 18167 24823 18173
rect 26234 18164 26240 18176
rect 26292 18164 26298 18216
rect 26329 18207 26387 18213
rect 26329 18173 26341 18207
rect 26375 18204 26387 18207
rect 27706 18204 27712 18216
rect 26375 18176 27712 18204
rect 26375 18173 26387 18176
rect 26329 18167 26387 18173
rect 27706 18164 27712 18176
rect 27764 18164 27770 18216
rect 27890 18164 27896 18216
rect 27948 18204 27954 18216
rect 28460 18204 28488 18244
rect 29273 18241 29285 18244
rect 29319 18241 29331 18275
rect 29273 18235 29331 18241
rect 33597 18275 33655 18281
rect 33597 18241 33609 18275
rect 33643 18272 33655 18275
rect 33980 18272 34008 18371
rect 35986 18368 35992 18380
rect 36044 18368 36050 18420
rect 43530 18408 43536 18420
rect 36280 18380 43536 18408
rect 34425 18343 34483 18349
rect 34425 18309 34437 18343
rect 34471 18340 34483 18343
rect 36280 18340 36308 18380
rect 43530 18368 43536 18380
rect 43588 18368 43594 18420
rect 48038 18408 48044 18420
rect 47999 18380 48044 18408
rect 48038 18368 48044 18380
rect 48096 18368 48102 18420
rect 48222 18368 48228 18420
rect 48280 18408 48286 18420
rect 48317 18411 48375 18417
rect 48317 18408 48329 18411
rect 48280 18380 48329 18408
rect 48280 18368 48286 18380
rect 48317 18377 48329 18380
rect 48363 18377 48375 18411
rect 48317 18371 48375 18377
rect 48961 18411 49019 18417
rect 48961 18377 48973 18411
rect 49007 18408 49019 18411
rect 49142 18408 49148 18420
rect 49007 18380 49148 18408
rect 49007 18377 49019 18380
rect 48961 18371 49019 18377
rect 49142 18368 49148 18380
rect 49200 18368 49206 18420
rect 49326 18408 49332 18420
rect 49287 18380 49332 18408
rect 49326 18368 49332 18380
rect 49384 18368 49390 18420
rect 52914 18368 52920 18420
rect 52972 18408 52978 18420
rect 54941 18411 54999 18417
rect 54941 18408 54953 18411
rect 52972 18380 54953 18408
rect 52972 18368 52978 18380
rect 54941 18377 54953 18380
rect 54987 18377 54999 18411
rect 54941 18371 54999 18377
rect 55309 18411 55367 18417
rect 55309 18377 55321 18411
rect 55355 18408 55367 18411
rect 56137 18411 56195 18417
rect 56137 18408 56149 18411
rect 55355 18380 56149 18408
rect 55355 18377 55367 18380
rect 55309 18371 55367 18377
rect 56137 18377 56149 18380
rect 56183 18408 56195 18411
rect 56226 18408 56232 18420
rect 56183 18380 56232 18408
rect 56183 18377 56195 18380
rect 56137 18371 56195 18377
rect 56226 18368 56232 18380
rect 56284 18368 56290 18420
rect 67450 18408 67456 18420
rect 67411 18380 67456 18408
rect 67450 18368 67456 18380
rect 67508 18368 67514 18420
rect 76374 18408 76380 18420
rect 67560 18380 76380 18408
rect 36446 18340 36452 18352
rect 34471 18312 36308 18340
rect 36407 18312 36452 18340
rect 34471 18309 34483 18312
rect 34425 18303 34483 18309
rect 36446 18300 36452 18312
rect 36504 18300 36510 18352
rect 39482 18300 39488 18352
rect 39540 18340 39546 18352
rect 41506 18340 41512 18352
rect 39540 18312 41512 18340
rect 39540 18300 39546 18312
rect 41506 18300 41512 18312
rect 41564 18300 41570 18352
rect 46198 18300 46204 18352
rect 46256 18340 46262 18352
rect 46256 18312 54688 18340
rect 46256 18300 46262 18312
rect 34330 18272 34336 18284
rect 33643 18244 34008 18272
rect 34243 18244 34336 18272
rect 33643 18241 33655 18244
rect 33597 18235 33655 18241
rect 34330 18232 34336 18244
rect 34388 18272 34394 18284
rect 35621 18275 35679 18281
rect 34388 18244 34652 18272
rect 34388 18232 34394 18244
rect 28626 18204 28632 18216
rect 27948 18176 28488 18204
rect 28587 18176 28632 18204
rect 27948 18164 27954 18176
rect 28626 18164 28632 18176
rect 28684 18164 28690 18216
rect 34514 18204 34520 18216
rect 34475 18176 34520 18204
rect 34514 18164 34520 18176
rect 34572 18164 34578 18216
rect 34624 18204 34652 18244
rect 35621 18241 35633 18275
rect 35667 18272 35679 18275
rect 35986 18272 35992 18284
rect 35667 18244 35992 18272
rect 35667 18241 35679 18244
rect 35621 18235 35679 18241
rect 35986 18232 35992 18244
rect 36044 18232 36050 18284
rect 36357 18275 36415 18281
rect 36357 18241 36369 18275
rect 36403 18272 36415 18275
rect 36814 18272 36820 18284
rect 36403 18244 36820 18272
rect 36403 18241 36415 18244
rect 36357 18235 36415 18241
rect 36814 18232 36820 18244
rect 36872 18232 36878 18284
rect 41877 18275 41935 18281
rect 41877 18241 41889 18275
rect 41923 18272 41935 18275
rect 42426 18272 42432 18284
rect 41923 18244 42432 18272
rect 41923 18241 41935 18244
rect 41877 18235 41935 18241
rect 42426 18232 42432 18244
rect 42484 18232 42490 18284
rect 44542 18232 44548 18284
rect 44600 18272 44606 18284
rect 45005 18275 45063 18281
rect 45005 18272 45017 18275
rect 44600 18244 45017 18272
rect 44600 18232 44606 18244
rect 45005 18241 45017 18244
rect 45051 18241 45063 18275
rect 45005 18235 45063 18241
rect 47762 18232 47768 18284
rect 47820 18272 47826 18284
rect 47857 18275 47915 18281
rect 47857 18272 47869 18275
rect 47820 18244 47869 18272
rect 47820 18232 47826 18244
rect 47857 18241 47869 18244
rect 47903 18272 47915 18275
rect 48222 18272 48228 18284
rect 47903 18244 48228 18272
rect 47903 18241 47915 18244
rect 47857 18235 47915 18241
rect 48222 18232 48228 18244
rect 48280 18232 48286 18284
rect 48777 18275 48835 18281
rect 48777 18241 48789 18275
rect 48823 18272 48835 18275
rect 48866 18272 48872 18284
rect 48823 18244 48872 18272
rect 48823 18241 48835 18244
rect 48777 18235 48835 18241
rect 48866 18232 48872 18244
rect 48924 18232 48930 18284
rect 49053 18275 49111 18281
rect 49053 18241 49065 18275
rect 49099 18272 49111 18275
rect 49326 18272 49332 18284
rect 49099 18244 49332 18272
rect 49099 18241 49111 18244
rect 49053 18235 49111 18241
rect 49326 18232 49332 18244
rect 49384 18272 49390 18284
rect 51810 18272 51816 18284
rect 49384 18244 51816 18272
rect 49384 18232 49390 18244
rect 51810 18232 51816 18244
rect 51868 18232 51874 18284
rect 54573 18275 54631 18281
rect 54573 18241 54585 18275
rect 54619 18241 54631 18275
rect 54660 18272 54688 18312
rect 54754 18300 54760 18352
rect 54812 18340 54818 18352
rect 55769 18343 55827 18349
rect 55769 18340 55781 18343
rect 54812 18312 55781 18340
rect 54812 18300 54818 18312
rect 55769 18309 55781 18312
rect 55815 18309 55827 18343
rect 67560 18340 67588 18380
rect 76374 18368 76380 18380
rect 76432 18368 76438 18420
rect 55769 18303 55827 18309
rect 55876 18312 67588 18340
rect 69477 18343 69535 18349
rect 55122 18272 55128 18284
rect 54660 18244 55128 18272
rect 54573 18235 54631 18241
rect 36262 18204 36268 18216
rect 34624 18176 36268 18204
rect 36262 18164 36268 18176
rect 36320 18164 36326 18216
rect 36633 18207 36691 18213
rect 36633 18173 36645 18207
rect 36679 18204 36691 18207
rect 36722 18204 36728 18216
rect 36679 18176 36728 18204
rect 36679 18173 36691 18176
rect 36633 18167 36691 18173
rect 36722 18164 36728 18176
rect 36780 18164 36786 18216
rect 44266 18164 44272 18216
rect 44324 18204 44330 18216
rect 47673 18207 47731 18213
rect 47673 18204 47685 18207
rect 44324 18176 47685 18204
rect 44324 18164 44330 18176
rect 47673 18173 47685 18176
rect 47719 18204 47731 18207
rect 51166 18204 51172 18216
rect 47719 18176 51172 18204
rect 47719 18173 47731 18176
rect 47673 18167 47731 18173
rect 51166 18164 51172 18176
rect 51224 18164 51230 18216
rect 54588 18204 54616 18235
rect 55122 18232 55128 18244
rect 55180 18232 55186 18284
rect 55398 18272 55404 18284
rect 55311 18244 55404 18272
rect 55398 18232 55404 18244
rect 55456 18272 55462 18284
rect 55876 18272 55904 18312
rect 69477 18309 69489 18343
rect 69523 18340 69535 18343
rect 78122 18340 78128 18352
rect 69523 18312 78128 18340
rect 69523 18309 69535 18312
rect 69477 18303 69535 18309
rect 78122 18300 78128 18312
rect 78180 18300 78186 18352
rect 55456 18244 55904 18272
rect 55456 18232 55462 18244
rect 55950 18232 55956 18284
rect 56008 18272 56014 18284
rect 56229 18275 56287 18281
rect 56008 18244 56053 18272
rect 56008 18232 56014 18244
rect 56229 18241 56241 18275
rect 56275 18272 56287 18275
rect 56318 18272 56324 18284
rect 56275 18244 56324 18272
rect 56275 18241 56287 18244
rect 56229 18235 56287 18241
rect 56318 18232 56324 18244
rect 56376 18272 56382 18284
rect 64874 18272 64880 18284
rect 56376 18244 64880 18272
rect 56376 18232 56382 18244
rect 64874 18232 64880 18244
rect 64932 18232 64938 18284
rect 67361 18275 67419 18281
rect 67361 18241 67373 18275
rect 67407 18272 67419 18275
rect 69198 18272 69204 18284
rect 67407 18244 69204 18272
rect 67407 18241 67419 18244
rect 67361 18235 67419 18241
rect 69198 18232 69204 18244
rect 69256 18232 69262 18284
rect 69385 18275 69443 18281
rect 69385 18241 69397 18275
rect 69431 18272 69443 18275
rect 69750 18272 69756 18284
rect 69431 18244 69756 18272
rect 69431 18241 69443 18244
rect 69385 18235 69443 18241
rect 69750 18232 69756 18244
rect 69808 18232 69814 18284
rect 70486 18272 70492 18284
rect 70447 18244 70492 18272
rect 70486 18232 70492 18244
rect 70544 18232 70550 18284
rect 70581 18275 70639 18281
rect 70581 18241 70593 18275
rect 70627 18272 70639 18275
rect 70627 18244 80054 18272
rect 70627 18241 70639 18244
rect 70581 18235 70639 18241
rect 55674 18204 55680 18216
rect 54588 18176 55680 18204
rect 55674 18164 55680 18176
rect 55732 18164 55738 18216
rect 60366 18204 60372 18216
rect 55775 18176 60372 18204
rect 7466 18096 7472 18148
rect 7524 18136 7530 18148
rect 48593 18139 48651 18145
rect 48593 18136 48605 18139
rect 7524 18108 48605 18136
rect 7524 18096 7530 18108
rect 48593 18105 48605 18108
rect 48639 18105 48651 18139
rect 48593 18099 48651 18105
rect 49602 18096 49608 18148
rect 49660 18136 49666 18148
rect 51074 18136 51080 18148
rect 49660 18108 51080 18136
rect 49660 18096 49666 18108
rect 51074 18096 51080 18108
rect 51132 18096 51138 18148
rect 53834 18096 53840 18148
rect 53892 18136 53898 18148
rect 53892 18108 54524 18136
rect 53892 18096 53898 18108
rect 1394 18068 1400 18080
rect 1355 18040 1400 18068
rect 1394 18028 1400 18040
rect 1452 18028 1458 18080
rect 24213 18071 24271 18077
rect 24213 18037 24225 18071
rect 24259 18068 24271 18071
rect 24946 18068 24952 18080
rect 24259 18040 24952 18068
rect 24259 18037 24271 18040
rect 24213 18031 24271 18037
rect 24946 18028 24952 18040
rect 25004 18028 25010 18080
rect 25685 18071 25743 18077
rect 25685 18037 25697 18071
rect 25731 18068 25743 18071
rect 26234 18068 26240 18080
rect 25731 18040 26240 18068
rect 25731 18037 25743 18040
rect 25685 18031 25743 18037
rect 26234 18028 26240 18040
rect 26292 18028 26298 18080
rect 27433 18071 27491 18077
rect 27433 18037 27445 18071
rect 27479 18068 27491 18071
rect 27614 18068 27620 18080
rect 27479 18040 27620 18068
rect 27479 18037 27491 18040
rect 27433 18031 27491 18037
rect 27614 18028 27620 18040
rect 27672 18028 27678 18080
rect 27798 18028 27804 18080
rect 27856 18068 27862 18080
rect 29089 18071 29147 18077
rect 29089 18068 29101 18071
rect 27856 18040 29101 18068
rect 27856 18028 27862 18040
rect 29089 18037 29101 18040
rect 29135 18037 29147 18071
rect 29089 18031 29147 18037
rect 33413 18071 33471 18077
rect 33413 18037 33425 18071
rect 33459 18068 33471 18071
rect 34974 18068 34980 18080
rect 33459 18040 34980 18068
rect 33459 18037 33471 18040
rect 33413 18031 33471 18037
rect 34974 18028 34980 18040
rect 35032 18028 35038 18080
rect 35437 18071 35495 18077
rect 35437 18037 35449 18071
rect 35483 18068 35495 18071
rect 36630 18068 36636 18080
rect 35483 18040 36636 18068
rect 35483 18037 35495 18040
rect 35437 18031 35495 18037
rect 36630 18028 36636 18040
rect 36688 18028 36694 18080
rect 41693 18071 41751 18077
rect 41693 18037 41705 18071
rect 41739 18068 41751 18071
rect 41782 18068 41788 18080
rect 41739 18040 41788 18068
rect 41739 18037 41751 18040
rect 41693 18031 41751 18037
rect 41782 18028 41788 18040
rect 41840 18028 41846 18080
rect 44821 18071 44879 18077
rect 44821 18037 44833 18071
rect 44867 18068 44879 18071
rect 45186 18068 45192 18080
rect 44867 18040 45192 18068
rect 44867 18037 44879 18040
rect 44821 18031 44879 18037
rect 45186 18028 45192 18040
rect 45244 18028 45250 18080
rect 54386 18068 54392 18080
rect 54347 18040 54392 18068
rect 54386 18028 54392 18040
rect 54444 18028 54450 18080
rect 54496 18068 54524 18108
rect 55122 18096 55128 18148
rect 55180 18136 55186 18148
rect 55775 18136 55803 18176
rect 60366 18164 60372 18176
rect 60424 18164 60430 18216
rect 60550 18164 60556 18216
rect 60608 18204 60614 18216
rect 61378 18204 61384 18216
rect 60608 18176 61384 18204
rect 60608 18164 60614 18176
rect 61378 18164 61384 18176
rect 61436 18164 61442 18216
rect 67545 18207 67603 18213
rect 67545 18204 67557 18207
rect 67376 18176 67557 18204
rect 67376 18148 67404 18176
rect 67545 18173 67557 18176
rect 67591 18173 67603 18207
rect 67545 18167 67603 18173
rect 69290 18164 69296 18216
rect 69348 18204 69354 18216
rect 69569 18207 69627 18213
rect 69569 18204 69581 18207
rect 69348 18176 69581 18204
rect 69348 18164 69354 18176
rect 69569 18173 69581 18176
rect 69615 18204 69627 18207
rect 70026 18204 70032 18216
rect 69615 18176 70032 18204
rect 69615 18173 69627 18176
rect 69569 18167 69627 18173
rect 70026 18164 70032 18176
rect 70084 18164 70090 18216
rect 70670 18204 70676 18216
rect 70631 18176 70676 18204
rect 70670 18164 70676 18176
rect 70728 18164 70734 18216
rect 80026 18204 80054 18244
rect 88058 18204 88064 18216
rect 80026 18176 88064 18204
rect 88058 18164 88064 18176
rect 88116 18164 88122 18216
rect 55180 18108 55803 18136
rect 55180 18096 55186 18108
rect 57974 18096 57980 18148
rect 58032 18136 58038 18148
rect 58710 18136 58716 18148
rect 58032 18108 58716 18136
rect 58032 18096 58038 18108
rect 58710 18096 58716 18108
rect 58768 18096 58774 18148
rect 67358 18096 67364 18148
rect 67416 18096 67422 18148
rect 70210 18096 70216 18148
rect 70268 18136 70274 18148
rect 70854 18136 70860 18148
rect 70268 18108 70860 18136
rect 70268 18096 70274 18108
rect 70854 18096 70860 18108
rect 70912 18096 70918 18148
rect 56318 18068 56324 18080
rect 54496 18040 56324 18068
rect 56318 18028 56324 18040
rect 56376 18068 56382 18080
rect 62758 18068 62764 18080
rect 56376 18040 62764 18068
rect 56376 18028 56382 18040
rect 62758 18028 62764 18040
rect 62816 18028 62822 18080
rect 66993 18071 67051 18077
rect 66993 18037 67005 18071
rect 67039 18068 67051 18071
rect 68094 18068 68100 18080
rect 67039 18040 68100 18068
rect 67039 18037 67051 18040
rect 66993 18031 67051 18037
rect 68094 18028 68100 18040
rect 68152 18028 68158 18080
rect 69014 18068 69020 18080
rect 68975 18040 69020 18068
rect 69014 18028 69020 18040
rect 69072 18028 69078 18080
rect 70121 18071 70179 18077
rect 70121 18037 70133 18071
rect 70167 18068 70179 18071
rect 70946 18068 70952 18080
rect 70167 18040 70952 18068
rect 70167 18037 70179 18040
rect 70121 18031 70179 18037
rect 70946 18028 70952 18040
rect 71004 18028 71010 18080
rect 1104 17978 88872 18000
rect 1104 17926 11924 17978
rect 11976 17926 11988 17978
rect 12040 17926 12052 17978
rect 12104 17926 12116 17978
rect 12168 17926 12180 17978
rect 12232 17926 33872 17978
rect 33924 17926 33936 17978
rect 33988 17926 34000 17978
rect 34052 17926 34064 17978
rect 34116 17926 34128 17978
rect 34180 17926 55820 17978
rect 55872 17926 55884 17978
rect 55936 17926 55948 17978
rect 56000 17926 56012 17978
rect 56064 17926 56076 17978
rect 56128 17926 77768 17978
rect 77820 17926 77832 17978
rect 77884 17926 77896 17978
rect 77948 17926 77960 17978
rect 78012 17926 78024 17978
rect 78076 17926 88872 17978
rect 1104 17904 88872 17926
rect 1946 17824 1952 17876
rect 2004 17864 2010 17876
rect 12526 17864 12532 17876
rect 2004 17836 12532 17864
rect 2004 17824 2010 17836
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12636 17836 28304 17864
rect 2866 17756 2872 17808
rect 2924 17796 2930 17808
rect 12636 17796 12664 17836
rect 2924 17768 12664 17796
rect 24765 17799 24823 17805
rect 2924 17756 2930 17768
rect 24765 17765 24777 17799
rect 24811 17765 24823 17799
rect 28276 17796 28304 17836
rect 28994 17824 29000 17876
rect 29052 17864 29058 17876
rect 29052 17836 31892 17864
rect 29052 17824 29058 17836
rect 28276 17768 28396 17796
rect 24765 17759 24823 17765
rect 2038 17688 2044 17740
rect 2096 17728 2102 17740
rect 12434 17728 12440 17740
rect 2096 17700 12440 17728
rect 2096 17688 2102 17700
rect 12434 17688 12440 17700
rect 12492 17688 12498 17740
rect 24780 17728 24808 17759
rect 25317 17731 25375 17737
rect 24780 17700 25268 17728
rect 2682 17620 2688 17672
rect 2740 17660 2746 17672
rect 12526 17660 12532 17672
rect 2740 17632 12532 17660
rect 2740 17620 2746 17632
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 12618 17620 12624 17672
rect 12676 17660 12682 17672
rect 24946 17660 24952 17672
rect 12676 17632 24808 17660
rect 24907 17632 24952 17660
rect 12676 17620 12682 17632
rect 4062 17552 4068 17604
rect 4120 17592 4126 17604
rect 24670 17592 24676 17604
rect 4120 17564 12434 17592
rect 4120 17552 4126 17564
rect 12406 17524 12434 17564
rect 12636 17564 24676 17592
rect 12636 17524 12664 17564
rect 24670 17552 24676 17564
rect 24728 17552 24734 17604
rect 12406 17496 12664 17524
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 24578 17524 24584 17536
rect 12768 17496 24584 17524
rect 12768 17484 12774 17496
rect 24578 17484 24584 17496
rect 24636 17484 24642 17536
rect 24780 17524 24808 17632
rect 24946 17620 24952 17632
rect 25004 17620 25010 17672
rect 25240 17660 25268 17700
rect 25317 17697 25329 17731
rect 25363 17728 25375 17731
rect 25774 17728 25780 17740
rect 25363 17700 25780 17728
rect 25363 17697 25375 17700
rect 25317 17691 25375 17697
rect 25774 17688 25780 17700
rect 25832 17688 25838 17740
rect 27338 17688 27344 17740
rect 27396 17728 27402 17740
rect 27614 17728 27620 17740
rect 27396 17700 27441 17728
rect 27575 17700 27620 17728
rect 27396 17688 27402 17700
rect 27614 17688 27620 17700
rect 27672 17688 27678 17740
rect 25593 17663 25651 17669
rect 25593 17660 25605 17663
rect 25240 17632 25605 17660
rect 25593 17629 25605 17632
rect 25639 17629 25651 17663
rect 27154 17660 27160 17672
rect 25593 17623 25651 17629
rect 26252 17632 27160 17660
rect 26252 17524 26280 17632
rect 27154 17620 27160 17632
rect 27212 17620 27218 17672
rect 28368 17660 28396 17768
rect 28442 17756 28448 17808
rect 28500 17796 28506 17808
rect 31754 17796 31760 17808
rect 28500 17768 31760 17796
rect 28500 17756 28506 17768
rect 31754 17756 31760 17768
rect 31812 17756 31818 17808
rect 31864 17796 31892 17836
rect 31938 17824 31944 17876
rect 31996 17864 32002 17876
rect 31996 17836 40816 17864
rect 31996 17824 32002 17836
rect 36081 17799 36139 17805
rect 31864 17768 34560 17796
rect 28534 17688 28540 17740
rect 28592 17728 28598 17740
rect 28721 17731 28779 17737
rect 28721 17728 28733 17731
rect 28592 17700 28733 17728
rect 28592 17688 28598 17700
rect 28721 17697 28733 17700
rect 28767 17728 28779 17731
rect 31110 17728 31116 17740
rect 28767 17700 31116 17728
rect 28767 17697 28779 17700
rect 28721 17691 28779 17697
rect 31110 17688 31116 17700
rect 31168 17688 31174 17740
rect 31202 17688 31208 17740
rect 31260 17728 31266 17740
rect 32125 17731 32183 17737
rect 32125 17728 32137 17731
rect 31260 17700 32137 17728
rect 31260 17688 31266 17700
rect 32125 17697 32137 17700
rect 32171 17697 32183 17731
rect 32125 17691 32183 17697
rect 32309 17731 32367 17737
rect 32309 17697 32321 17731
rect 32355 17728 32367 17731
rect 32398 17728 32404 17740
rect 32355 17700 32404 17728
rect 32355 17697 32367 17700
rect 32309 17691 32367 17697
rect 32398 17688 32404 17700
rect 32456 17688 32462 17740
rect 33413 17663 33471 17669
rect 33413 17660 33425 17663
rect 27264 17632 28304 17660
rect 28368 17632 33425 17660
rect 26970 17592 26976 17604
rect 26883 17564 26976 17592
rect 26970 17552 26976 17564
rect 27028 17592 27034 17604
rect 27264 17592 27292 17632
rect 27028 17564 27292 17592
rect 27028 17552 27034 17564
rect 24780 17496 26280 17524
rect 26326 17484 26332 17536
rect 26384 17524 26390 17536
rect 28074 17524 28080 17536
rect 26384 17496 28080 17524
rect 26384 17484 26390 17496
rect 28074 17484 28080 17496
rect 28132 17484 28138 17536
rect 28276 17524 28304 17632
rect 33413 17629 33425 17632
rect 33459 17629 33471 17663
rect 33594 17660 33600 17672
rect 33555 17632 33600 17660
rect 33413 17623 33471 17629
rect 33594 17620 33600 17632
rect 33652 17620 33658 17672
rect 33873 17663 33931 17669
rect 33873 17629 33885 17663
rect 33919 17660 33931 17663
rect 34422 17660 34428 17672
rect 33919 17632 34428 17660
rect 33919 17629 33931 17632
rect 33873 17623 33931 17629
rect 34422 17620 34428 17632
rect 34480 17620 34486 17672
rect 28350 17552 28356 17604
rect 28408 17592 28414 17604
rect 31938 17592 31944 17604
rect 28408 17564 31944 17592
rect 28408 17552 28414 17564
rect 31938 17552 31944 17564
rect 31996 17552 32002 17604
rect 32122 17552 32128 17604
rect 32180 17592 32186 17604
rect 34532 17592 34560 17768
rect 36081 17765 36093 17799
rect 36127 17796 36139 17799
rect 36262 17796 36268 17808
rect 36127 17768 36268 17796
rect 36127 17765 36139 17768
rect 36081 17759 36139 17765
rect 36262 17756 36268 17768
rect 36320 17756 36326 17808
rect 37550 17756 37556 17808
rect 37608 17796 37614 17808
rect 40494 17796 40500 17808
rect 37608 17768 40500 17796
rect 37608 17756 37614 17768
rect 40494 17756 40500 17768
rect 40552 17756 40558 17808
rect 40788 17796 40816 17836
rect 41506 17824 41512 17876
rect 41564 17864 41570 17876
rect 46198 17864 46204 17876
rect 41564 17836 46204 17864
rect 41564 17824 41570 17836
rect 46198 17824 46204 17836
rect 46256 17824 46262 17876
rect 46290 17824 46296 17876
rect 46348 17864 46354 17876
rect 48774 17864 48780 17876
rect 46348 17836 48636 17864
rect 48735 17836 48780 17864
rect 46348 17824 46354 17836
rect 41325 17799 41383 17805
rect 41325 17796 41337 17799
rect 40788 17768 41337 17796
rect 37826 17688 37832 17740
rect 37884 17728 37890 17740
rect 40678 17728 40684 17740
rect 37884 17700 40684 17728
rect 37884 17688 37890 17700
rect 40678 17688 40684 17700
rect 40736 17688 40742 17740
rect 40788 17737 40816 17768
rect 41325 17765 41337 17768
rect 41371 17765 41383 17799
rect 41325 17759 41383 17765
rect 42889 17799 42947 17805
rect 42889 17765 42901 17799
rect 42935 17765 42947 17799
rect 44542 17796 44548 17808
rect 44503 17768 44548 17796
rect 42889 17759 42947 17765
rect 40773 17731 40831 17737
rect 40773 17697 40785 17731
rect 40819 17697 40831 17731
rect 40773 17691 40831 17697
rect 40957 17731 41015 17737
rect 40957 17697 40969 17731
rect 41003 17728 41015 17731
rect 41414 17728 41420 17740
rect 41003 17700 41420 17728
rect 41003 17697 41015 17700
rect 40957 17691 41015 17697
rect 41414 17688 41420 17700
rect 41472 17688 41478 17740
rect 34698 17660 34704 17672
rect 34659 17632 34704 17660
rect 34698 17620 34704 17632
rect 34756 17660 34762 17672
rect 36541 17663 36599 17669
rect 36541 17660 36553 17663
rect 34756 17632 36553 17660
rect 34756 17620 34762 17632
rect 36541 17629 36553 17632
rect 36587 17629 36599 17663
rect 36541 17623 36599 17629
rect 36630 17620 36636 17672
rect 36688 17660 36694 17672
rect 36797 17663 36855 17669
rect 36797 17660 36809 17663
rect 36688 17632 36809 17660
rect 36688 17620 36694 17632
rect 36797 17629 36809 17632
rect 36843 17629 36855 17663
rect 41322 17660 41328 17672
rect 36797 17623 36855 17629
rect 36924 17632 41328 17660
rect 34790 17592 34796 17604
rect 32180 17564 33916 17592
rect 34532 17564 34796 17592
rect 32180 17552 32186 17564
rect 30006 17524 30012 17536
rect 28276 17496 30012 17524
rect 30006 17484 30012 17496
rect 30064 17484 30070 17536
rect 30834 17484 30840 17536
rect 30892 17524 30898 17536
rect 31665 17527 31723 17533
rect 31665 17524 31677 17527
rect 30892 17496 31677 17524
rect 30892 17484 30898 17496
rect 31665 17493 31677 17496
rect 31711 17493 31723 17527
rect 31665 17487 31723 17493
rect 32033 17527 32091 17533
rect 32033 17493 32045 17527
rect 32079 17524 32091 17527
rect 32490 17524 32496 17536
rect 32079 17496 32496 17524
rect 32079 17493 32091 17496
rect 32033 17487 32091 17493
rect 32490 17484 32496 17496
rect 32548 17484 32554 17536
rect 33778 17524 33784 17536
rect 33739 17496 33784 17524
rect 33778 17484 33784 17496
rect 33836 17484 33842 17536
rect 33888 17524 33916 17564
rect 34790 17552 34796 17564
rect 34848 17552 34854 17604
rect 34974 17601 34980 17604
rect 34968 17592 34980 17601
rect 34935 17564 34980 17592
rect 34968 17555 34980 17564
rect 34974 17552 34980 17555
rect 35032 17552 35038 17604
rect 36924 17592 36952 17632
rect 41322 17620 41328 17632
rect 41380 17620 41386 17672
rect 41506 17660 41512 17672
rect 41467 17632 41512 17660
rect 41506 17620 41512 17632
rect 41564 17620 41570 17672
rect 41616 17632 42748 17660
rect 40681 17595 40739 17601
rect 35084 17564 36952 17592
rect 37016 17564 40632 17592
rect 35084 17524 35112 17564
rect 33888 17496 35112 17524
rect 35158 17484 35164 17536
rect 35216 17524 35222 17536
rect 37016 17524 37044 17564
rect 35216 17496 37044 17524
rect 37921 17527 37979 17533
rect 35216 17484 35222 17496
rect 37921 17493 37933 17527
rect 37967 17524 37979 17527
rect 38194 17524 38200 17536
rect 37967 17496 38200 17524
rect 37967 17493 37979 17496
rect 37921 17487 37979 17493
rect 38194 17484 38200 17496
rect 38252 17484 38258 17536
rect 40218 17484 40224 17536
rect 40276 17524 40282 17536
rect 40313 17527 40371 17533
rect 40313 17524 40325 17527
rect 40276 17496 40325 17524
rect 40276 17484 40282 17496
rect 40313 17493 40325 17496
rect 40359 17493 40371 17527
rect 40604 17524 40632 17564
rect 40681 17561 40693 17595
rect 40727 17592 40739 17595
rect 41414 17592 41420 17604
rect 40727 17564 41420 17592
rect 40727 17561 40739 17564
rect 40681 17555 40739 17561
rect 41414 17552 41420 17564
rect 41472 17552 41478 17604
rect 41616 17524 41644 17632
rect 41782 17601 41788 17604
rect 41776 17592 41788 17601
rect 41743 17564 41788 17592
rect 41776 17555 41788 17564
rect 41782 17552 41788 17555
rect 41840 17552 41846 17604
rect 42720 17592 42748 17632
rect 42794 17620 42800 17672
rect 42852 17660 42858 17672
rect 42904 17660 42932 17759
rect 44542 17756 44548 17768
rect 44600 17756 44606 17808
rect 45462 17796 45468 17808
rect 45423 17768 45468 17796
rect 45462 17756 45468 17768
rect 45520 17756 45526 17808
rect 47489 17799 47547 17805
rect 47489 17765 47501 17799
rect 47535 17765 47547 17799
rect 48608 17796 48636 17836
rect 48774 17824 48780 17836
rect 48832 17824 48838 17876
rect 50154 17864 50160 17876
rect 50115 17836 50160 17864
rect 50154 17824 50160 17836
rect 50212 17824 50218 17876
rect 51074 17824 51080 17876
rect 51132 17864 51138 17876
rect 60550 17864 60556 17876
rect 51132 17836 60556 17864
rect 51132 17824 51138 17836
rect 60550 17824 60556 17836
rect 60608 17824 60614 17876
rect 62758 17824 62764 17876
rect 62816 17864 62822 17876
rect 70210 17864 70216 17876
rect 62816 17836 70216 17864
rect 62816 17824 62822 17836
rect 70210 17824 70216 17836
rect 70268 17824 70274 17876
rect 48608 17768 50476 17796
rect 47489 17759 47547 17765
rect 43257 17731 43315 17737
rect 43257 17697 43269 17731
rect 43303 17728 43315 17731
rect 43438 17728 43444 17740
rect 43303 17700 43444 17728
rect 43303 17697 43315 17700
rect 43257 17691 43315 17697
rect 43438 17688 43444 17700
rect 43496 17688 43502 17740
rect 47504 17728 47532 17759
rect 48866 17728 48872 17740
rect 44376 17700 47532 17728
rect 48779 17700 48872 17728
rect 43165 17663 43223 17669
rect 43165 17660 43177 17663
rect 42852 17632 43177 17660
rect 42852 17620 42858 17632
rect 43165 17629 43177 17632
rect 43211 17629 43223 17663
rect 43165 17623 43223 17629
rect 43346 17620 43352 17672
rect 43404 17660 43410 17672
rect 44266 17660 44272 17672
rect 43404 17632 44272 17660
rect 43404 17620 43410 17632
rect 44266 17620 44272 17632
rect 44324 17620 44330 17672
rect 44376 17669 44404 17700
rect 48866 17688 48872 17700
rect 48924 17728 48930 17740
rect 50448 17728 50476 17768
rect 54294 17756 54300 17808
rect 54352 17796 54358 17808
rect 55306 17796 55312 17808
rect 54352 17768 55312 17796
rect 54352 17756 54358 17768
rect 55306 17756 55312 17768
rect 55364 17796 55370 17808
rect 55364 17768 55536 17796
rect 55364 17756 55370 17768
rect 53006 17728 53012 17740
rect 48924 17700 50384 17728
rect 50448 17700 53012 17728
rect 48924 17688 48930 17700
rect 44361 17663 44419 17669
rect 44361 17629 44373 17663
rect 44407 17629 44419 17663
rect 45646 17660 45652 17672
rect 45607 17632 45652 17660
rect 44361 17623 44419 17629
rect 44376 17592 44404 17623
rect 45646 17620 45652 17632
rect 45704 17620 45710 17672
rect 45922 17660 45928 17672
rect 45883 17632 45928 17660
rect 45922 17620 45928 17632
rect 45980 17620 45986 17672
rect 46934 17660 46940 17672
rect 46895 17632 46940 17660
rect 46934 17620 46940 17632
rect 46992 17620 46998 17672
rect 47210 17660 47216 17672
rect 47171 17632 47216 17660
rect 47210 17620 47216 17632
rect 47268 17620 47274 17672
rect 47357 17663 47415 17669
rect 47357 17629 47369 17663
rect 47403 17660 47415 17663
rect 48130 17660 48136 17672
rect 47403 17632 47992 17660
rect 48091 17632 48136 17660
rect 47403 17629 47415 17632
rect 47357 17623 47415 17629
rect 42720 17564 44404 17592
rect 46566 17552 46572 17604
rect 46624 17592 46630 17604
rect 47121 17595 47179 17601
rect 47121 17592 47133 17595
rect 46624 17564 47133 17592
rect 46624 17552 46630 17564
rect 47121 17561 47133 17564
rect 47167 17561 47179 17595
rect 47854 17592 47860 17604
rect 47121 17555 47179 17561
rect 47320 17564 47860 17592
rect 40604 17496 41644 17524
rect 40313 17487 40371 17493
rect 41690 17484 41696 17536
rect 41748 17524 41754 17536
rect 45833 17527 45891 17533
rect 45833 17524 45845 17527
rect 41748 17496 45845 17524
rect 41748 17484 41754 17496
rect 45833 17493 45845 17496
rect 45879 17524 45891 17527
rect 47320 17524 47348 17564
rect 47854 17552 47860 17564
rect 47912 17552 47918 17604
rect 47964 17592 47992 17632
rect 48130 17620 48136 17632
rect 48188 17620 48194 17672
rect 48222 17620 48228 17672
rect 48280 17660 48286 17672
rect 48409 17663 48467 17669
rect 48409 17660 48421 17663
rect 48280 17632 48421 17660
rect 48280 17620 48286 17632
rect 48409 17629 48421 17632
rect 48455 17629 48467 17663
rect 48884 17660 48912 17688
rect 48961 17663 49019 17669
rect 48961 17660 48973 17663
rect 48884 17632 48973 17660
rect 48409 17623 48467 17629
rect 48961 17629 48973 17632
rect 49007 17629 49019 17663
rect 49142 17660 49148 17672
rect 49103 17632 49148 17660
rect 48961 17623 49019 17629
rect 49142 17620 49148 17632
rect 49200 17620 49206 17672
rect 49234 17620 49240 17672
rect 49292 17660 49298 17672
rect 50356 17669 50384 17700
rect 53006 17688 53012 17700
rect 53064 17688 53070 17740
rect 53098 17688 53104 17740
rect 53156 17728 53162 17740
rect 55398 17728 55404 17740
rect 53156 17700 55404 17728
rect 53156 17688 53162 17700
rect 55398 17688 55404 17700
rect 55456 17688 55462 17740
rect 50341 17663 50399 17669
rect 49292 17632 49337 17660
rect 49292 17620 49298 17632
rect 50341 17629 50353 17663
rect 50387 17660 50399 17663
rect 50522 17660 50528 17672
rect 50387 17632 50528 17660
rect 50387 17629 50399 17632
rect 50341 17623 50399 17629
rect 50522 17620 50528 17632
rect 50580 17620 50586 17672
rect 50617 17663 50675 17669
rect 50617 17629 50629 17663
rect 50663 17660 50675 17663
rect 52178 17660 52184 17672
rect 50663 17632 52184 17660
rect 50663 17629 50675 17632
rect 50617 17623 50675 17629
rect 52178 17620 52184 17632
rect 52236 17620 52242 17672
rect 53282 17660 53288 17672
rect 53243 17632 53288 17660
rect 53282 17620 53288 17632
rect 53340 17620 53346 17672
rect 53561 17663 53619 17669
rect 53561 17629 53573 17663
rect 53607 17660 53619 17663
rect 53926 17660 53932 17672
rect 53607 17632 53932 17660
rect 53607 17629 53619 17632
rect 53561 17623 53619 17629
rect 53926 17620 53932 17632
rect 53984 17620 53990 17672
rect 54110 17660 54116 17672
rect 54071 17632 54116 17660
rect 54110 17620 54116 17632
rect 54168 17620 54174 17672
rect 54389 17663 54447 17669
rect 54389 17629 54401 17663
rect 54435 17660 54447 17663
rect 54570 17660 54576 17672
rect 54435 17632 54576 17660
rect 54435 17629 54447 17632
rect 54389 17623 54447 17629
rect 54570 17620 54576 17632
rect 54628 17620 54634 17672
rect 54662 17620 54668 17672
rect 54720 17660 54726 17672
rect 55306 17660 55312 17672
rect 54720 17632 55312 17660
rect 54720 17620 54726 17632
rect 55306 17620 55312 17632
rect 55364 17620 55370 17672
rect 55508 17669 55536 17768
rect 56410 17756 56416 17808
rect 56468 17796 56474 17808
rect 60458 17796 60464 17808
rect 56468 17768 60464 17796
rect 56468 17756 56474 17768
rect 60458 17756 60464 17768
rect 60516 17756 60522 17808
rect 60642 17756 60648 17808
rect 60700 17796 60706 17808
rect 61010 17796 61016 17808
rect 60700 17768 61016 17796
rect 60700 17756 60706 17768
rect 61010 17756 61016 17768
rect 61068 17756 61074 17808
rect 61102 17756 61108 17808
rect 61160 17796 61166 17808
rect 64506 17796 64512 17808
rect 61160 17768 64512 17796
rect 61160 17756 61166 17768
rect 64506 17756 64512 17768
rect 64564 17756 64570 17808
rect 64969 17799 65027 17805
rect 64969 17765 64981 17799
rect 65015 17796 65027 17799
rect 65518 17796 65524 17808
rect 65015 17768 65524 17796
rect 65015 17765 65027 17768
rect 64969 17759 65027 17765
rect 65518 17756 65524 17768
rect 65576 17756 65582 17808
rect 67913 17799 67971 17805
rect 67913 17765 67925 17799
rect 67959 17796 67971 17799
rect 68462 17796 68468 17808
rect 67959 17768 68468 17796
rect 67959 17765 67971 17768
rect 67913 17759 67971 17765
rect 68462 17756 68468 17768
rect 68520 17756 68526 17808
rect 55674 17728 55680 17740
rect 55635 17700 55680 17728
rect 55674 17688 55680 17700
rect 55732 17688 55738 17740
rect 55968 17700 58204 17728
rect 55493 17663 55551 17669
rect 55493 17629 55505 17663
rect 55539 17629 55551 17663
rect 55493 17623 55551 17629
rect 55582 17620 55588 17672
rect 55640 17660 55646 17672
rect 55968 17660 55996 17700
rect 55640 17632 55996 17660
rect 55640 17620 55646 17632
rect 56042 17620 56048 17672
rect 56100 17660 56106 17672
rect 56229 17663 56287 17669
rect 56100 17632 56145 17660
rect 56100 17620 56106 17632
rect 56229 17629 56241 17663
rect 56275 17660 56287 17663
rect 56318 17660 56324 17672
rect 56275 17632 56324 17660
rect 56275 17629 56287 17632
rect 56229 17623 56287 17629
rect 56318 17620 56324 17632
rect 56376 17620 56382 17672
rect 56413 17663 56471 17669
rect 56413 17629 56425 17663
rect 56459 17660 56471 17663
rect 56965 17663 57023 17669
rect 56965 17660 56977 17663
rect 56459 17632 56977 17660
rect 56459 17629 56471 17632
rect 56413 17623 56471 17629
rect 56965 17629 56977 17632
rect 57011 17629 57023 17663
rect 56965 17623 57023 17629
rect 53098 17592 53104 17604
rect 47964 17564 53104 17592
rect 53098 17552 53104 17564
rect 53156 17552 53162 17604
rect 58176 17592 58204 17700
rect 58881 17700 60780 17728
rect 58710 17660 58716 17672
rect 58671 17632 58716 17660
rect 58710 17620 58716 17632
rect 58768 17620 58774 17672
rect 58881 17669 58909 17700
rect 58851 17663 58909 17669
rect 58851 17629 58863 17663
rect 58897 17629 58909 17663
rect 58851 17623 58909 17629
rect 58986 17620 58992 17672
rect 59044 17660 59050 17672
rect 59127 17663 59185 17669
rect 59044 17632 59089 17660
rect 59044 17620 59050 17632
rect 59127 17629 59139 17663
rect 59173 17660 59185 17663
rect 59262 17660 59268 17672
rect 59173 17632 59268 17660
rect 59173 17629 59185 17632
rect 59127 17623 59185 17629
rect 59262 17620 59268 17632
rect 59320 17620 59326 17672
rect 59906 17620 59912 17672
rect 59964 17660 59970 17672
rect 60001 17663 60059 17669
rect 60001 17660 60013 17663
rect 59964 17632 60013 17660
rect 59964 17620 59970 17632
rect 60001 17629 60013 17632
rect 60047 17629 60059 17663
rect 60752 17660 60780 17700
rect 60826 17688 60832 17740
rect 60884 17728 60890 17740
rect 61657 17731 61715 17737
rect 61657 17728 61669 17731
rect 60884 17700 61669 17728
rect 60884 17688 60890 17700
rect 61657 17697 61669 17700
rect 61703 17697 61715 17731
rect 61657 17691 61715 17697
rect 61562 17660 61568 17672
rect 60752 17632 61568 17660
rect 60001 17623 60059 17629
rect 61562 17620 61568 17632
rect 61620 17620 61626 17672
rect 61672 17660 61700 17691
rect 62758 17688 62764 17740
rect 62816 17728 62822 17740
rect 68557 17731 68615 17737
rect 68557 17728 68569 17731
rect 62816 17700 65656 17728
rect 62816 17688 62822 17700
rect 62390 17660 62396 17672
rect 61672 17632 62396 17660
rect 62390 17620 62396 17632
rect 62448 17620 62454 17672
rect 62482 17620 62488 17672
rect 62540 17660 62546 17672
rect 62669 17663 62727 17669
rect 62669 17660 62681 17663
rect 62540 17632 62681 17660
rect 62540 17620 62546 17632
rect 62669 17629 62681 17632
rect 62715 17629 62727 17663
rect 65150 17660 65156 17672
rect 65111 17632 65156 17660
rect 62669 17623 62727 17629
rect 65150 17620 65156 17632
rect 65208 17620 65214 17672
rect 65628 17669 65656 17700
rect 67606 17700 68569 17728
rect 65613 17663 65671 17669
rect 65613 17629 65625 17663
rect 65659 17660 65671 17663
rect 67606 17660 67634 17700
rect 68557 17697 68569 17700
rect 68603 17728 68615 17731
rect 68603 17700 69152 17728
rect 68603 17697 68615 17700
rect 68557 17691 68615 17697
rect 68094 17660 68100 17672
rect 65659 17632 67634 17660
rect 68055 17632 68100 17660
rect 65659 17629 65671 17632
rect 65613 17623 65671 17629
rect 68094 17620 68100 17632
rect 68152 17620 68158 17672
rect 68462 17620 68468 17672
rect 68520 17660 68526 17672
rect 68833 17663 68891 17669
rect 68833 17660 68845 17663
rect 68520 17632 68845 17660
rect 68520 17620 68526 17632
rect 68833 17629 68845 17632
rect 68879 17629 68891 17663
rect 69124 17660 69152 17700
rect 69198 17688 69204 17740
rect 69256 17728 69262 17740
rect 69937 17731 69995 17737
rect 69937 17728 69949 17731
rect 69256 17700 69949 17728
rect 69256 17688 69262 17700
rect 69937 17697 69949 17700
rect 69983 17697 69995 17731
rect 69937 17691 69995 17697
rect 69658 17660 69664 17672
rect 69124 17632 69664 17660
rect 68833 17623 68891 17629
rect 69658 17620 69664 17632
rect 69716 17620 69722 17672
rect 70946 17660 70952 17672
rect 70907 17632 70952 17660
rect 70946 17620 70952 17632
rect 71004 17620 71010 17672
rect 53208 17564 56916 17592
rect 58176 17564 59216 17592
rect 45879 17496 47348 17524
rect 45879 17493 45891 17496
rect 45833 17487 45891 17493
rect 47394 17484 47400 17536
rect 47452 17524 47458 17536
rect 47949 17527 48007 17533
rect 47949 17524 47961 17527
rect 47452 17496 47961 17524
rect 47452 17484 47458 17496
rect 47949 17493 47961 17496
rect 47995 17493 48007 17527
rect 47949 17487 48007 17493
rect 48317 17527 48375 17533
rect 48317 17493 48329 17527
rect 48363 17524 48375 17527
rect 48958 17524 48964 17536
rect 48363 17496 48964 17524
rect 48363 17493 48375 17496
rect 48317 17487 48375 17493
rect 48958 17484 48964 17496
rect 49016 17484 49022 17536
rect 49142 17484 49148 17536
rect 49200 17524 49206 17536
rect 50525 17527 50583 17533
rect 50525 17524 50537 17527
rect 49200 17496 50537 17524
rect 49200 17484 49206 17496
rect 50525 17493 50537 17496
rect 50571 17524 50583 17527
rect 53208 17524 53236 17564
rect 53374 17524 53380 17536
rect 53432 17533 53438 17536
rect 50571 17496 53236 17524
rect 53341 17496 53380 17524
rect 50571 17493 50583 17496
rect 50525 17487 50583 17493
rect 53374 17484 53380 17496
rect 53432 17487 53441 17533
rect 53469 17527 53527 17533
rect 53469 17493 53481 17527
rect 53515 17524 53527 17527
rect 53558 17524 53564 17536
rect 53515 17496 53564 17524
rect 53515 17493 53527 17496
rect 53469 17487 53527 17493
rect 53432 17484 53438 17487
rect 53558 17484 53564 17496
rect 53616 17484 53622 17536
rect 53650 17484 53656 17536
rect 53708 17524 53714 17536
rect 53929 17527 53987 17533
rect 53929 17524 53941 17527
rect 53708 17496 53941 17524
rect 53708 17484 53714 17496
rect 53929 17493 53941 17496
rect 53975 17493 53987 17527
rect 53929 17487 53987 17493
rect 54297 17527 54355 17533
rect 54297 17493 54309 17527
rect 54343 17524 54355 17527
rect 56410 17524 56416 17536
rect 54343 17496 56416 17524
rect 54343 17493 54355 17496
rect 54297 17487 54355 17493
rect 56410 17484 56416 17496
rect 56468 17484 56474 17536
rect 56594 17484 56600 17536
rect 56652 17524 56658 17536
rect 56781 17527 56839 17533
rect 56781 17524 56793 17527
rect 56652 17496 56793 17524
rect 56652 17484 56658 17496
rect 56781 17493 56793 17496
rect 56827 17493 56839 17527
rect 56888 17524 56916 17564
rect 59078 17524 59084 17536
rect 56888 17496 59084 17524
rect 56781 17487 56839 17493
rect 59078 17484 59084 17496
rect 59136 17484 59142 17536
rect 59188 17524 59216 17564
rect 59354 17552 59360 17604
rect 59412 17592 59418 17604
rect 60642 17592 60648 17604
rect 59412 17564 60648 17592
rect 59412 17552 59418 17564
rect 60642 17552 60648 17564
rect 60700 17552 60706 17604
rect 60826 17592 60832 17604
rect 60787 17564 60832 17592
rect 60826 17552 60832 17564
rect 60884 17592 60890 17604
rect 61473 17595 61531 17601
rect 61473 17592 61485 17595
rect 60884 17564 61485 17592
rect 60884 17552 60890 17564
rect 61473 17561 61485 17564
rect 61519 17561 61531 17595
rect 62114 17592 62120 17604
rect 61473 17555 61531 17561
rect 61580 17564 62120 17592
rect 59265 17527 59323 17533
rect 59265 17524 59277 17527
rect 59188 17496 59277 17524
rect 59265 17493 59277 17496
rect 59311 17524 59323 17527
rect 59722 17524 59728 17536
rect 59311 17496 59728 17524
rect 59311 17493 59323 17496
rect 59265 17487 59323 17493
rect 59722 17484 59728 17496
rect 59780 17484 59786 17536
rect 59817 17527 59875 17533
rect 59817 17493 59829 17527
rect 59863 17524 59875 17527
rect 60366 17524 60372 17536
rect 59863 17496 60372 17524
rect 59863 17493 59875 17496
rect 59817 17487 59875 17493
rect 60366 17484 60372 17496
rect 60424 17484 60430 17536
rect 60918 17524 60924 17536
rect 60879 17496 60924 17524
rect 60918 17484 60924 17496
rect 60976 17484 60982 17536
rect 61010 17484 61016 17536
rect 61068 17524 61074 17536
rect 61580 17524 61608 17564
rect 62114 17552 62120 17564
rect 62172 17552 62178 17604
rect 62209 17595 62267 17601
rect 62209 17561 62221 17595
rect 62255 17592 62267 17595
rect 62255 17564 65104 17592
rect 62255 17561 62267 17564
rect 62209 17555 62267 17561
rect 62574 17524 62580 17536
rect 61068 17496 61608 17524
rect 62535 17496 62580 17524
rect 61068 17484 61074 17496
rect 62574 17484 62580 17496
rect 62632 17484 62638 17536
rect 65076 17524 65104 17564
rect 65518 17552 65524 17604
rect 65576 17592 65582 17604
rect 65858 17595 65916 17601
rect 65858 17592 65870 17595
rect 65576 17564 65870 17592
rect 65576 17552 65582 17564
rect 65858 17561 65870 17564
rect 65904 17561 65916 17595
rect 65858 17555 65916 17561
rect 65996 17564 67634 17592
rect 65996 17524 66024 17564
rect 65076 17496 66024 17524
rect 66714 17484 66720 17536
rect 66772 17524 66778 17536
rect 66993 17527 67051 17533
rect 66993 17524 67005 17527
rect 66772 17496 67005 17524
rect 66772 17484 66778 17496
rect 66993 17493 67005 17496
rect 67039 17493 67051 17527
rect 67606 17524 67634 17564
rect 68278 17552 68284 17604
rect 68336 17592 68342 17604
rect 68554 17592 68560 17604
rect 68336 17564 68560 17592
rect 68336 17552 68342 17564
rect 68554 17552 68560 17564
rect 68612 17552 68618 17604
rect 75178 17592 75184 17604
rect 69492 17564 75184 17592
rect 69492 17524 69520 17564
rect 75178 17552 75184 17564
rect 75236 17552 75242 17604
rect 67606 17496 69520 17524
rect 66993 17487 67051 17493
rect 69566 17484 69572 17536
rect 69624 17524 69630 17536
rect 70486 17524 70492 17536
rect 69624 17496 70492 17524
rect 69624 17484 69630 17496
rect 70486 17484 70492 17496
rect 70544 17484 70550 17536
rect 70762 17524 70768 17536
rect 70723 17496 70768 17524
rect 70762 17484 70768 17496
rect 70820 17484 70826 17536
rect 1104 17434 88872 17456
rect 1104 17382 22898 17434
rect 22950 17382 22962 17434
rect 23014 17382 23026 17434
rect 23078 17382 23090 17434
rect 23142 17382 23154 17434
rect 23206 17382 44846 17434
rect 44898 17382 44910 17434
rect 44962 17382 44974 17434
rect 45026 17382 45038 17434
rect 45090 17382 45102 17434
rect 45154 17382 66794 17434
rect 66846 17382 66858 17434
rect 66910 17382 66922 17434
rect 66974 17382 66986 17434
rect 67038 17382 67050 17434
rect 67102 17382 88872 17434
rect 1104 17360 88872 17382
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12492 17292 22692 17320
rect 12492 17280 12498 17292
rect 22370 17252 22376 17264
rect 6886 17224 22376 17252
rect 1762 17184 1768 17196
rect 1723 17156 1768 17184
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17116 2007 17119
rect 6886 17116 6914 17224
rect 22370 17212 22376 17224
rect 22428 17212 22434 17264
rect 22664 17252 22692 17292
rect 22738 17280 22744 17332
rect 22796 17320 22802 17332
rect 23201 17323 23259 17329
rect 23201 17320 23213 17323
rect 22796 17292 23213 17320
rect 22796 17280 22802 17292
rect 23201 17289 23213 17292
rect 23247 17320 23259 17323
rect 24029 17323 24087 17329
rect 24029 17320 24041 17323
rect 23247 17292 24041 17320
rect 23247 17289 23259 17292
rect 23201 17283 23259 17289
rect 24029 17289 24041 17292
rect 24075 17289 24087 17323
rect 28350 17320 28356 17332
rect 24029 17283 24087 17289
rect 24136 17292 28356 17320
rect 24136 17252 24164 17292
rect 28350 17280 28356 17292
rect 28408 17280 28414 17332
rect 30006 17280 30012 17332
rect 30064 17320 30070 17332
rect 30064 17292 80054 17320
rect 30064 17280 30070 17292
rect 22664 17224 24164 17252
rect 24670 17212 24676 17264
rect 24728 17252 24734 17264
rect 27516 17255 27574 17261
rect 24728 17224 26372 17252
rect 24728 17212 24734 17224
rect 23934 17184 23940 17196
rect 23895 17156 23940 17184
rect 23934 17144 23940 17156
rect 23992 17144 23998 17196
rect 24946 17184 24952 17196
rect 24907 17156 24952 17184
rect 24946 17144 24952 17156
rect 25004 17144 25010 17196
rect 26234 17184 26240 17196
rect 26195 17156 26240 17184
rect 26234 17144 26240 17156
rect 26292 17144 26298 17196
rect 26344 17184 26372 17224
rect 27516 17221 27528 17255
rect 27562 17252 27574 17255
rect 27798 17252 27804 17264
rect 27562 17224 27804 17252
rect 27562 17221 27574 17224
rect 27516 17215 27574 17221
rect 27798 17212 27804 17224
rect 27856 17212 27862 17264
rect 32122 17252 32128 17264
rect 27908 17224 32128 17252
rect 27908 17184 27936 17224
rect 32122 17212 32128 17224
rect 32180 17212 32186 17264
rect 32214 17212 32220 17264
rect 32272 17252 32278 17264
rect 32585 17255 32643 17261
rect 32585 17252 32597 17255
rect 32272 17224 32597 17252
rect 32272 17212 32278 17224
rect 32585 17221 32597 17224
rect 32631 17221 32643 17255
rect 32585 17215 32643 17221
rect 32766 17212 32772 17264
rect 32824 17252 32830 17264
rect 35710 17261 35716 17264
rect 35704 17252 35716 17261
rect 32824 17224 34008 17252
rect 35671 17224 35716 17252
rect 32824 17212 32830 17224
rect 26344 17156 27936 17184
rect 28074 17144 28080 17196
rect 28132 17184 28138 17196
rect 31665 17187 31723 17193
rect 28132 17156 28304 17184
rect 28132 17144 28138 17156
rect 1995 17088 6914 17116
rect 1995 17085 2007 17088
rect 1949 17079 2007 17085
rect 24210 17076 24216 17128
rect 24268 17116 24274 17128
rect 24670 17116 24676 17128
rect 24268 17088 24676 17116
rect 24268 17076 24274 17088
rect 24670 17076 24676 17088
rect 24728 17076 24734 17128
rect 26970 17076 26976 17128
rect 27028 17116 27034 17128
rect 27246 17116 27252 17128
rect 27028 17088 27252 17116
rect 27028 17076 27034 17088
rect 27246 17076 27252 17088
rect 27304 17076 27310 17128
rect 23569 17051 23627 17057
rect 23569 17017 23581 17051
rect 23615 17048 23627 17051
rect 24946 17048 24952 17060
rect 23615 17020 24952 17048
rect 23615 17017 23627 17020
rect 23569 17011 23627 17017
rect 24946 17008 24952 17020
rect 25004 17008 25010 17060
rect 28276 17048 28304 17156
rect 31665 17153 31677 17187
rect 31711 17184 31723 17187
rect 32493 17187 32551 17193
rect 31711 17156 31984 17184
rect 31711 17153 31723 17156
rect 31665 17147 31723 17153
rect 28350 17076 28356 17128
rect 28408 17116 28414 17128
rect 31754 17116 31760 17128
rect 28408 17088 31760 17116
rect 28408 17076 28414 17088
rect 31754 17076 31760 17088
rect 31812 17076 31818 17128
rect 31956 17048 31984 17156
rect 32493 17153 32505 17187
rect 32539 17184 32551 17187
rect 32674 17184 32680 17196
rect 32539 17156 32680 17184
rect 32539 17153 32551 17156
rect 32493 17147 32551 17153
rect 32674 17144 32680 17156
rect 32732 17144 32738 17196
rect 33594 17184 33600 17196
rect 33555 17156 33600 17184
rect 33594 17144 33600 17156
rect 33652 17144 33658 17196
rect 33778 17184 33784 17196
rect 33739 17156 33784 17184
rect 33778 17144 33784 17156
rect 33836 17144 33842 17196
rect 33873 17187 33931 17193
rect 33873 17153 33885 17187
rect 33919 17153 33931 17187
rect 33980 17184 34008 17224
rect 35704 17215 35716 17224
rect 35710 17212 35716 17215
rect 35768 17212 35774 17264
rect 37826 17252 37832 17264
rect 37787 17224 37832 17252
rect 37826 17212 37832 17224
rect 37884 17212 37890 17264
rect 39482 17252 39488 17264
rect 37936 17224 39488 17252
rect 37550 17184 37556 17196
rect 33980 17156 37556 17184
rect 33873 17147 33931 17153
rect 32030 17076 32036 17128
rect 32088 17116 32094 17128
rect 32088 17088 32260 17116
rect 32088 17076 32094 17088
rect 32125 17051 32183 17057
rect 32125 17048 32137 17051
rect 28276 17020 31754 17048
rect 31956 17020 32137 17048
rect 24765 16983 24823 16989
rect 24765 16949 24777 16983
rect 24811 16980 24823 16983
rect 25682 16980 25688 16992
rect 24811 16952 25688 16980
rect 24811 16949 24823 16952
rect 24765 16943 24823 16949
rect 25682 16940 25688 16952
rect 25740 16940 25746 16992
rect 26053 16983 26111 16989
rect 26053 16949 26065 16983
rect 26099 16980 26111 16983
rect 26234 16980 26240 16992
rect 26099 16952 26240 16980
rect 26099 16949 26111 16952
rect 26053 16943 26111 16949
rect 26234 16940 26240 16952
rect 26292 16940 26298 16992
rect 28534 16940 28540 16992
rect 28592 16980 28598 16992
rect 28629 16983 28687 16989
rect 28629 16980 28641 16983
rect 28592 16952 28641 16980
rect 28592 16940 28598 16952
rect 28629 16949 28641 16952
rect 28675 16949 28687 16983
rect 31478 16980 31484 16992
rect 31439 16952 31484 16980
rect 28629 16943 28687 16949
rect 31478 16940 31484 16952
rect 31536 16940 31542 16992
rect 31726 16980 31754 17020
rect 32125 17017 32137 17020
rect 32171 17017 32183 17051
rect 32232 17048 32260 17088
rect 32398 17076 32404 17128
rect 32456 17116 32462 17128
rect 32766 17116 32772 17128
rect 32456 17088 32772 17116
rect 32456 17076 32462 17088
rect 32766 17076 32772 17088
rect 32824 17076 32830 17128
rect 33888 17116 33916 17147
rect 37550 17144 37556 17156
rect 37608 17144 37614 17196
rect 37642 17144 37648 17196
rect 37700 17184 37706 17196
rect 37936 17184 37964 17224
rect 39482 17212 39488 17224
rect 39540 17212 39546 17264
rect 41506 17252 41512 17264
rect 39592 17224 41512 17252
rect 38194 17184 38200 17196
rect 37700 17156 37964 17184
rect 38155 17156 38200 17184
rect 37700 17144 37706 17156
rect 38194 17144 38200 17156
rect 38252 17144 38258 17196
rect 39592 17193 39620 17224
rect 41506 17212 41512 17224
rect 41564 17252 41570 17264
rect 41874 17252 41880 17264
rect 41564 17224 41880 17252
rect 41564 17212 41570 17224
rect 41874 17212 41880 17224
rect 41932 17212 41938 17264
rect 42886 17252 42892 17264
rect 42847 17224 42892 17252
rect 42886 17212 42892 17224
rect 42944 17212 42950 17264
rect 44726 17252 44732 17264
rect 43732 17224 44732 17252
rect 39577 17187 39635 17193
rect 39577 17153 39589 17187
rect 39623 17153 39635 17187
rect 39577 17147 39635 17153
rect 39844 17187 39902 17193
rect 39844 17153 39856 17187
rect 39890 17184 39902 17187
rect 40126 17184 40132 17196
rect 39890 17156 40132 17184
rect 39890 17153 39902 17156
rect 39844 17147 39902 17153
rect 40126 17144 40132 17156
rect 40184 17144 40190 17196
rect 41230 17184 41236 17196
rect 41191 17156 41236 17184
rect 41230 17144 41236 17156
rect 41288 17184 41294 17196
rect 41782 17184 41788 17196
rect 41288 17156 41788 17184
rect 41288 17144 41294 17156
rect 41782 17144 41788 17156
rect 41840 17144 41846 17196
rect 42242 17144 42248 17196
rect 42300 17184 42306 17196
rect 42794 17184 42800 17196
rect 42300 17156 42656 17184
rect 42755 17156 42800 17184
rect 42300 17144 42306 17156
rect 34330 17116 34336 17128
rect 32876 17088 34336 17116
rect 32876 17048 32904 17088
rect 34330 17076 34336 17088
rect 34388 17076 34394 17128
rect 35434 17116 35440 17128
rect 34716 17088 35440 17116
rect 34716 17060 34744 17088
rect 35434 17076 35440 17088
rect 35492 17076 35498 17128
rect 41601 17119 41659 17125
rect 41601 17085 41613 17119
rect 41647 17085 41659 17119
rect 41601 17079 41659 17085
rect 32232 17020 32904 17048
rect 32125 17011 32183 17017
rect 33042 17008 33048 17060
rect 33100 17048 33106 17060
rect 34698 17048 34704 17060
rect 33100 17020 34704 17048
rect 33100 17008 33106 17020
rect 34698 17008 34704 17020
rect 34756 17008 34762 17060
rect 36446 17008 36452 17060
rect 36504 17048 36510 17060
rect 39574 17048 39580 17060
rect 36504 17020 39580 17048
rect 36504 17008 36510 17020
rect 39574 17008 39580 17020
rect 39632 17008 39638 17060
rect 40957 17051 41015 17057
rect 40957 17017 40969 17051
rect 41003 17048 41015 17051
rect 41414 17048 41420 17060
rect 41003 17020 41420 17048
rect 41003 17017 41015 17020
rect 40957 17011 41015 17017
rect 41414 17008 41420 17020
rect 41472 17008 41478 17060
rect 41616 17048 41644 17079
rect 41690 17076 41696 17128
rect 41748 17116 41754 17128
rect 42628 17116 42656 17156
rect 42794 17144 42800 17156
rect 42852 17144 42858 17196
rect 43533 17187 43591 17193
rect 43533 17153 43545 17187
rect 43579 17184 43591 17187
rect 43622 17184 43628 17196
rect 43579 17156 43628 17184
rect 43579 17153 43591 17156
rect 43533 17147 43591 17153
rect 43622 17144 43628 17156
rect 43680 17144 43686 17196
rect 43732 17193 43760 17224
rect 44726 17212 44732 17224
rect 44784 17212 44790 17264
rect 45738 17252 45744 17264
rect 44836 17224 45744 17252
rect 44836 17193 44864 17224
rect 45738 17212 45744 17224
rect 45796 17252 45802 17264
rect 45796 17224 47624 17252
rect 45796 17212 45802 17224
rect 45094 17193 45100 17196
rect 43717 17187 43775 17193
rect 43717 17153 43729 17187
rect 43763 17153 43775 17187
rect 43717 17147 43775 17153
rect 43809 17187 43867 17193
rect 43809 17153 43821 17187
rect 43855 17153 43867 17187
rect 43809 17147 43867 17153
rect 44821 17187 44879 17193
rect 44821 17153 44833 17187
rect 44867 17153 44879 17187
rect 45088 17184 45100 17193
rect 45055 17156 45100 17184
rect 44821 17147 44879 17153
rect 45088 17147 45100 17156
rect 42981 17119 43039 17125
rect 42981 17116 42993 17119
rect 41748 17088 42564 17116
rect 42628 17088 42993 17116
rect 41748 17076 41754 17088
rect 42426 17048 42432 17060
rect 41616 17020 42104 17048
rect 42387 17020 42432 17048
rect 33413 16983 33471 16989
rect 33413 16980 33425 16983
rect 31726 16952 33425 16980
rect 33413 16949 33425 16952
rect 33459 16949 33471 16983
rect 36814 16980 36820 16992
rect 36775 16952 36820 16980
rect 33413 16943 33471 16949
rect 36814 16940 36820 16952
rect 36872 16940 36878 16992
rect 38289 16983 38347 16989
rect 38289 16949 38301 16983
rect 38335 16980 38347 16983
rect 40310 16980 40316 16992
rect 38335 16952 40316 16980
rect 38335 16949 38347 16952
rect 38289 16943 38347 16949
rect 40310 16940 40316 16952
rect 40368 16940 40374 16992
rect 41506 16940 41512 16992
rect 41564 16980 41570 16992
rect 41969 16983 42027 16989
rect 41969 16980 41981 16983
rect 41564 16952 41981 16980
rect 41564 16940 41570 16952
rect 41969 16949 41981 16952
rect 42015 16949 42027 16983
rect 42076 16980 42104 17020
rect 42426 17008 42432 17020
rect 42484 17008 42490 17060
rect 42536 17048 42564 17088
rect 42981 17085 42993 17088
rect 43027 17085 43039 17119
rect 42981 17079 43039 17085
rect 43070 17076 43076 17128
rect 43128 17116 43134 17128
rect 43824 17116 43852 17147
rect 45094 17144 45100 17147
rect 45152 17144 45158 17196
rect 46566 17184 46572 17196
rect 46527 17156 46572 17184
rect 46566 17144 46572 17156
rect 46624 17144 46630 17196
rect 46750 17184 46756 17196
rect 46711 17156 46756 17184
rect 46750 17144 46756 17156
rect 46808 17144 46814 17196
rect 46937 17187 46995 17193
rect 46937 17153 46949 17187
rect 46983 17153 46995 17187
rect 46937 17147 46995 17153
rect 46952 17116 46980 17147
rect 47026 17144 47032 17196
rect 47084 17184 47090 17196
rect 47596 17193 47624 17224
rect 47946 17212 47952 17264
rect 48004 17252 48010 17264
rect 53650 17252 53656 17264
rect 48004 17224 53420 17252
rect 53611 17224 53656 17252
rect 48004 17212 48010 17224
rect 47581 17187 47639 17193
rect 47084 17156 47129 17184
rect 47084 17144 47090 17156
rect 47581 17153 47593 17187
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 47670 17144 47676 17196
rect 47728 17184 47734 17196
rect 47837 17187 47895 17193
rect 47837 17184 47849 17187
rect 47728 17156 47849 17184
rect 47728 17144 47734 17156
rect 47837 17153 47849 17156
rect 47883 17153 47895 17187
rect 47837 17147 47895 17153
rect 48314 17144 48320 17196
rect 48372 17184 48378 17196
rect 48774 17184 48780 17196
rect 48372 17156 48780 17184
rect 48372 17144 48378 17156
rect 48774 17144 48780 17156
rect 48832 17144 48838 17196
rect 49694 17184 49700 17196
rect 49655 17156 49700 17184
rect 49694 17144 49700 17156
rect 49752 17144 49758 17196
rect 49878 17184 49884 17196
rect 49839 17156 49884 17184
rect 49878 17144 49884 17156
rect 49936 17144 49942 17196
rect 49973 17187 50031 17193
rect 49973 17153 49985 17187
rect 50019 17184 50031 17187
rect 50522 17184 50528 17196
rect 50019 17156 50528 17184
rect 50019 17153 50031 17156
rect 49973 17147 50031 17153
rect 50522 17144 50528 17156
rect 50580 17144 50586 17196
rect 50798 17144 50804 17196
rect 50856 17184 50862 17196
rect 50985 17187 51043 17193
rect 50856 17156 50901 17184
rect 50856 17144 50862 17156
rect 50985 17153 50997 17187
rect 51031 17184 51043 17187
rect 51537 17187 51595 17193
rect 51537 17184 51549 17187
rect 51031 17156 51549 17184
rect 51031 17153 51043 17156
rect 50985 17147 51043 17153
rect 51537 17153 51549 17156
rect 51583 17153 51595 17187
rect 51537 17147 51595 17153
rect 52917 17187 52975 17193
rect 52917 17153 52929 17187
rect 52963 17184 52975 17187
rect 52963 17156 53328 17184
rect 52963 17153 52975 17156
rect 52917 17147 52975 17153
rect 49418 17116 49424 17128
rect 43128 17088 43852 17116
rect 46216 17088 46980 17116
rect 48608 17088 49424 17116
rect 43128 17076 43134 17088
rect 42536 17020 43760 17048
rect 43346 16980 43352 16992
rect 42076 16952 43352 16980
rect 41969 16943 42027 16949
rect 43346 16940 43352 16952
rect 43404 16940 43410 16992
rect 43533 16983 43591 16989
rect 43533 16949 43545 16983
rect 43579 16980 43591 16983
rect 43622 16980 43628 16992
rect 43579 16952 43628 16980
rect 43579 16949 43591 16952
rect 43533 16943 43591 16949
rect 43622 16940 43628 16952
rect 43680 16940 43686 16992
rect 43732 16980 43760 17020
rect 43806 17008 43812 17060
rect 43864 17048 43870 17060
rect 44818 17048 44824 17060
rect 43864 17020 44824 17048
rect 43864 17008 43870 17020
rect 44818 17008 44824 17020
rect 44876 17008 44882 17060
rect 46216 17057 46244 17088
rect 46201 17051 46259 17057
rect 46201 17017 46213 17051
rect 46247 17017 46259 17051
rect 46201 17011 46259 17017
rect 46290 17008 46296 17060
rect 46348 17048 46354 17060
rect 46348 17020 46980 17048
rect 46348 17008 46354 17020
rect 46842 16980 46848 16992
rect 43732 16952 46848 16980
rect 46842 16940 46848 16952
rect 46900 16940 46906 16992
rect 46952 16980 46980 17020
rect 48608 16980 48636 17088
rect 49418 17076 49424 17088
rect 49476 17076 49482 17128
rect 49712 17116 49740 17144
rect 50154 17116 50160 17128
rect 49712 17088 50160 17116
rect 50154 17076 50160 17088
rect 50212 17076 50218 17128
rect 50617 17119 50675 17125
rect 50617 17085 50629 17119
rect 50663 17116 50675 17119
rect 51074 17116 51080 17128
rect 50663 17088 51080 17116
rect 50663 17085 50675 17088
rect 50617 17079 50675 17085
rect 51074 17076 51080 17088
rect 51132 17076 51138 17128
rect 51184 17088 53236 17116
rect 48958 17048 48964 17060
rect 48919 17020 48964 17048
rect 48958 17008 48964 17020
rect 49016 17008 49022 17060
rect 49513 17051 49571 17057
rect 49513 17017 49525 17051
rect 49559 17048 49571 17051
rect 49602 17048 49608 17060
rect 49559 17020 49608 17048
rect 49559 17017 49571 17020
rect 49513 17011 49571 17017
rect 49602 17008 49608 17020
rect 49660 17008 49666 17060
rect 49970 17008 49976 17060
rect 50028 17048 50034 17060
rect 51184 17048 51212 17088
rect 53101 17051 53159 17057
rect 53101 17048 53113 17051
rect 50028 17020 51212 17048
rect 51276 17020 53113 17048
rect 50028 17008 50034 17020
rect 46952 16952 48636 16980
rect 50341 16983 50399 16989
rect 50341 16949 50353 16983
rect 50387 16980 50399 16983
rect 50798 16980 50804 16992
rect 50387 16952 50804 16980
rect 50387 16949 50399 16952
rect 50341 16943 50399 16949
rect 50798 16940 50804 16952
rect 50856 16940 50862 16992
rect 50982 16940 50988 16992
rect 51040 16980 51046 16992
rect 51276 16980 51304 17020
rect 53101 17017 53113 17020
rect 53147 17017 53159 17051
rect 53101 17011 53159 17017
rect 51040 16952 51304 16980
rect 51040 16940 51046 16952
rect 51350 16940 51356 16992
rect 51408 16980 51414 16992
rect 53208 16980 53236 17088
rect 53300 17048 53328 17156
rect 53392 17116 53420 17224
rect 53650 17212 53656 17224
rect 53708 17212 53714 17264
rect 54202 17252 54208 17264
rect 53852 17224 54208 17252
rect 53466 17144 53472 17196
rect 53524 17184 53530 17196
rect 53852 17193 53880 17224
rect 54202 17212 54208 17224
rect 54260 17212 54266 17264
rect 54386 17261 54392 17264
rect 54380 17252 54392 17261
rect 54347 17224 54392 17252
rect 54380 17215 54392 17224
rect 54386 17212 54392 17215
rect 54444 17212 54450 17264
rect 54478 17212 54484 17264
rect 54536 17252 54542 17264
rect 54536 17224 58388 17252
rect 54536 17212 54542 17224
rect 53745 17187 53803 17193
rect 53524 17156 53569 17184
rect 53524 17144 53530 17156
rect 53745 17153 53757 17187
rect 53791 17153 53803 17187
rect 53745 17147 53803 17153
rect 53837 17187 53895 17193
rect 53837 17153 53849 17187
rect 53883 17153 53895 17187
rect 53837 17147 53895 17153
rect 53760 17116 53788 17147
rect 53926 17144 53932 17196
rect 53984 17184 53990 17196
rect 53984 17156 56272 17184
rect 53984 17144 53990 17156
rect 53392 17088 53788 17116
rect 54113 17119 54171 17125
rect 54113 17085 54125 17119
rect 54159 17085 54171 17119
rect 54113 17079 54171 17085
rect 53742 17048 53748 17060
rect 53300 17020 53748 17048
rect 53742 17008 53748 17020
rect 53800 17008 53806 17060
rect 53834 17008 53840 17060
rect 53892 17048 53898 17060
rect 54021 17051 54079 17057
rect 54021 17048 54033 17051
rect 53892 17020 54033 17048
rect 53892 17008 53898 17020
rect 54021 17017 54033 17020
rect 54067 17017 54079 17051
rect 54021 17011 54079 17017
rect 53926 16980 53932 16992
rect 51408 16952 51453 16980
rect 53208 16952 53932 16980
rect 51408 16940 51414 16952
rect 53926 16940 53932 16952
rect 53984 16940 53990 16992
rect 54128 16980 54156 17079
rect 55306 17076 55312 17128
rect 55364 17116 55370 17128
rect 56042 17116 56048 17128
rect 55364 17088 56048 17116
rect 55364 17076 55370 17088
rect 56042 17076 56048 17088
rect 56100 17116 56106 17128
rect 56137 17119 56195 17125
rect 56137 17116 56149 17119
rect 56100 17088 56149 17116
rect 56100 17076 56106 17088
rect 56137 17085 56149 17088
rect 56183 17085 56195 17119
rect 56244 17116 56272 17156
rect 56318 17144 56324 17196
rect 56376 17184 56382 17196
rect 56376 17156 56421 17184
rect 56376 17144 56382 17156
rect 56778 17144 56784 17196
rect 56836 17184 56842 17196
rect 57698 17184 57704 17196
rect 56836 17156 57704 17184
rect 56836 17144 56842 17156
rect 57698 17144 57704 17156
rect 57756 17144 57762 17196
rect 57882 17184 57888 17196
rect 57843 17156 57888 17184
rect 57882 17144 57888 17156
rect 57940 17144 57946 17196
rect 58066 17184 58072 17196
rect 58027 17156 58072 17184
rect 58066 17144 58072 17156
rect 58124 17144 58130 17196
rect 58158 17144 58164 17196
rect 58216 17184 58222 17196
rect 58360 17184 58388 17224
rect 58526 17212 58532 17264
rect 58584 17252 58590 17264
rect 58713 17255 58771 17261
rect 58713 17252 58725 17255
rect 58584 17224 58725 17252
rect 58584 17212 58590 17224
rect 58713 17221 58725 17224
rect 58759 17221 58771 17255
rect 59906 17252 59912 17264
rect 59867 17224 59912 17252
rect 58713 17215 58771 17221
rect 59906 17212 59912 17224
rect 59964 17212 59970 17264
rect 62666 17252 62672 17264
rect 60292 17224 62672 17252
rect 58802 17184 58808 17196
rect 58216 17156 58261 17184
rect 58360 17156 58808 17184
rect 58216 17144 58222 17156
rect 58802 17144 58808 17156
rect 58860 17144 58866 17196
rect 58894 17144 58900 17196
rect 58952 17184 58958 17196
rect 59081 17187 59139 17193
rect 58952 17156 58997 17184
rect 58952 17144 58958 17156
rect 59081 17153 59093 17187
rect 59127 17153 59139 17187
rect 59081 17147 59139 17153
rect 59173 17187 59231 17193
rect 59173 17153 59185 17187
rect 59219 17184 59231 17187
rect 59219 17156 59676 17184
rect 59219 17153 59231 17156
rect 59173 17147 59231 17153
rect 58618 17116 58624 17128
rect 56244 17088 58624 17116
rect 56137 17079 56195 17085
rect 58618 17076 58624 17088
rect 58676 17076 58682 17128
rect 59096 17116 59124 17147
rect 59262 17116 59268 17128
rect 59096 17088 59268 17116
rect 59262 17076 59268 17088
rect 59320 17076 59326 17128
rect 59538 17116 59544 17128
rect 59499 17088 59544 17116
rect 59538 17076 59544 17088
rect 59596 17076 59602 17128
rect 59648 17116 59676 17156
rect 59722 17144 59728 17196
rect 59780 17184 59786 17196
rect 60292 17193 60320 17224
rect 62666 17212 62672 17224
rect 62724 17212 62730 17264
rect 63129 17255 63187 17261
rect 63129 17221 63141 17255
rect 63175 17252 63187 17255
rect 64414 17252 64420 17264
rect 63175 17224 64420 17252
rect 63175 17221 63187 17224
rect 63129 17215 63187 17221
rect 64414 17212 64420 17224
rect 64472 17212 64478 17264
rect 65153 17255 65211 17261
rect 65153 17252 65165 17255
rect 64524 17224 65165 17252
rect 60277 17187 60335 17193
rect 59780 17156 59825 17184
rect 59780 17144 59786 17156
rect 60277 17153 60289 17187
rect 60323 17153 60335 17187
rect 60277 17147 60335 17153
rect 60366 17144 60372 17196
rect 60424 17184 60430 17196
rect 60533 17187 60591 17193
rect 60533 17184 60545 17187
rect 60424 17156 60545 17184
rect 60424 17144 60430 17156
rect 60533 17153 60545 17156
rect 60579 17153 60591 17187
rect 62114 17184 62120 17196
rect 62075 17156 62120 17184
rect 60533 17147 60591 17153
rect 62114 17144 62120 17156
rect 62172 17144 62178 17196
rect 62390 17144 62396 17196
rect 62448 17184 62454 17196
rect 63313 17187 63371 17193
rect 63313 17184 63325 17187
rect 62448 17156 63325 17184
rect 62448 17144 62454 17156
rect 63313 17153 63325 17156
rect 63359 17153 63371 17187
rect 63494 17184 63500 17196
rect 63455 17156 63500 17184
rect 63313 17147 63371 17153
rect 63494 17144 63500 17156
rect 63552 17144 63558 17196
rect 63589 17187 63647 17193
rect 63589 17153 63601 17187
rect 63635 17184 63647 17187
rect 63678 17184 63684 17196
rect 63635 17156 63684 17184
rect 63635 17153 63647 17156
rect 63589 17147 63647 17153
rect 63678 17144 63684 17156
rect 63736 17144 63742 17196
rect 64524 17193 64552 17224
rect 65153 17221 65165 17224
rect 65199 17221 65211 17255
rect 69382 17252 69388 17264
rect 65153 17215 65211 17221
rect 65260 17224 69388 17252
rect 64509 17187 64567 17193
rect 64509 17153 64521 17187
rect 64555 17153 64567 17187
rect 64509 17147 64567 17153
rect 64782 17144 64788 17196
rect 64840 17184 64846 17196
rect 64877 17187 64935 17193
rect 64877 17184 64889 17187
rect 64840 17156 64889 17184
rect 64840 17144 64846 17156
rect 64877 17153 64889 17156
rect 64923 17153 64935 17187
rect 64877 17147 64935 17153
rect 64966 17144 64972 17196
rect 65024 17184 65030 17196
rect 65024 17156 65069 17184
rect 65024 17144 65030 17156
rect 59814 17116 59820 17128
rect 59648 17088 59820 17116
rect 59814 17076 59820 17088
rect 59872 17116 59878 17128
rect 59998 17116 60004 17128
rect 59872 17088 60004 17116
rect 59872 17076 59878 17088
rect 59998 17076 60004 17088
rect 60056 17076 60062 17128
rect 61378 17076 61384 17128
rect 61436 17116 61442 17128
rect 64690 17116 64696 17128
rect 61436 17088 64696 17116
rect 61436 17076 61442 17088
rect 64690 17076 64696 17088
rect 64748 17076 64754 17128
rect 65260 17116 65288 17224
rect 69382 17212 69388 17224
rect 69440 17212 69446 17264
rect 70670 17212 70676 17264
rect 70728 17252 70734 17264
rect 80026 17252 80054 17292
rect 87598 17252 87604 17264
rect 70728 17224 73844 17252
rect 80026 17224 87604 17252
rect 70728 17212 70734 17224
rect 66165 17188 66223 17193
rect 66165 17187 66392 17188
rect 66165 17153 66177 17187
rect 66211 17184 66392 17187
rect 66714 17184 66720 17196
rect 66211 17160 66720 17184
rect 66211 17153 66223 17160
rect 66364 17156 66720 17160
rect 66165 17147 66223 17153
rect 66714 17144 66720 17156
rect 66772 17184 66778 17196
rect 66901 17187 66959 17193
rect 66901 17184 66913 17187
rect 66772 17156 66913 17184
rect 66772 17144 66778 17156
rect 66901 17153 66913 17156
rect 66947 17153 66959 17187
rect 66901 17147 66959 17153
rect 66990 17144 66996 17196
rect 67048 17184 67054 17196
rect 68925 17187 68983 17193
rect 67048 17156 67093 17184
rect 67048 17144 67054 17156
rect 68925 17153 68937 17187
rect 68971 17184 68983 17187
rect 69014 17184 69020 17196
rect 68971 17156 69020 17184
rect 68971 17153 68983 17156
rect 68925 17147 68983 17153
rect 69014 17144 69020 17156
rect 69072 17144 69078 17196
rect 69106 17144 69112 17196
rect 69164 17184 69170 17196
rect 69937 17187 69995 17193
rect 69164 17156 69796 17184
rect 69164 17144 69170 17156
rect 65076 17088 65288 17116
rect 66257 17119 66315 17125
rect 55122 17008 55128 17060
rect 55180 17048 55186 17060
rect 55861 17051 55919 17057
rect 55861 17048 55873 17051
rect 55180 17020 55873 17048
rect 55180 17008 55186 17020
rect 55861 17017 55873 17020
rect 55907 17048 55919 17051
rect 56318 17048 56324 17060
rect 55907 17020 56324 17048
rect 55907 17017 55919 17020
rect 55861 17011 55919 17017
rect 56318 17008 56324 17020
rect 56376 17048 56382 17060
rect 60274 17048 60280 17060
rect 56376 17020 60280 17048
rect 56376 17008 56382 17020
rect 60274 17008 60280 17020
rect 60332 17008 60338 17060
rect 65076 17048 65104 17088
rect 66257 17085 66269 17119
rect 66303 17085 66315 17119
rect 66438 17116 66444 17128
rect 66399 17088 66444 17116
rect 66257 17079 66315 17085
rect 61488 17020 65104 17048
rect 55214 16980 55220 16992
rect 54128 16952 55220 16980
rect 55214 16940 55220 16952
rect 55272 16940 55278 16992
rect 55306 16940 55312 16992
rect 55364 16980 55370 16992
rect 55493 16983 55551 16989
rect 55493 16980 55505 16983
rect 55364 16952 55505 16980
rect 55364 16940 55370 16952
rect 55493 16949 55505 16952
rect 55539 16949 55551 16983
rect 56502 16980 56508 16992
rect 56463 16952 56508 16980
rect 55493 16943 55551 16949
rect 56502 16940 56508 16952
rect 56560 16940 56566 16992
rect 57885 16983 57943 16989
rect 57885 16949 57897 16983
rect 57931 16980 57943 16983
rect 59262 16980 59268 16992
rect 57931 16952 59268 16980
rect 57931 16949 57943 16952
rect 57885 16943 57943 16949
rect 59262 16940 59268 16952
rect 59320 16940 59326 16992
rect 60642 16940 60648 16992
rect 60700 16980 60706 16992
rect 61488 16980 61516 17020
rect 65150 17008 65156 17060
rect 65208 17048 65214 17060
rect 65797 17051 65855 17057
rect 65797 17048 65809 17051
rect 65208 17020 65809 17048
rect 65208 17008 65214 17020
rect 65797 17017 65809 17020
rect 65843 17017 65855 17051
rect 66272 17048 66300 17079
rect 66438 17076 66444 17088
rect 66496 17076 66502 17128
rect 66530 17076 66536 17128
rect 66588 17116 66594 17128
rect 69658 17116 69664 17128
rect 66588 17088 68968 17116
rect 69619 17088 69664 17116
rect 66588 17076 66594 17088
rect 68554 17048 68560 17060
rect 65797 17011 65855 17017
rect 66180 17020 68560 17048
rect 61654 16980 61660 16992
rect 60700 16952 61516 16980
rect 61615 16952 61660 16980
rect 60700 16940 60706 16952
rect 61654 16940 61660 16952
rect 61712 16940 61718 16992
rect 62209 16983 62267 16989
rect 62209 16949 62221 16983
rect 62255 16980 62267 16983
rect 62574 16980 62580 16992
rect 62255 16952 62580 16980
rect 62255 16949 62267 16952
rect 62209 16943 62267 16949
rect 62574 16940 62580 16952
rect 62632 16980 62638 16992
rect 64230 16980 64236 16992
rect 62632 16952 64236 16980
rect 62632 16940 62638 16952
rect 64230 16940 64236 16952
rect 64288 16940 64294 16992
rect 64325 16983 64383 16989
rect 64325 16949 64337 16983
rect 64371 16980 64383 16983
rect 65334 16980 65340 16992
rect 64371 16952 65340 16980
rect 64371 16949 64383 16952
rect 64325 16943 64383 16949
rect 65334 16940 65340 16952
rect 65392 16940 65398 16992
rect 65521 16983 65579 16989
rect 65521 16949 65533 16983
rect 65567 16980 65579 16983
rect 66180 16980 66208 17020
rect 68554 17008 68560 17020
rect 68612 17008 68618 17060
rect 68646 17008 68652 17060
rect 68704 17048 68710 17060
rect 68741 17051 68799 17057
rect 68741 17048 68753 17051
rect 68704 17020 68753 17048
rect 68704 17008 68710 17020
rect 68741 17017 68753 17020
rect 68787 17017 68799 17051
rect 68741 17011 68799 17017
rect 65567 16952 66208 16980
rect 68940 16980 68968 17088
rect 69658 17076 69664 17088
rect 69716 17076 69722 17128
rect 69768 17116 69796 17156
rect 69937 17153 69949 17187
rect 69983 17184 69995 17187
rect 70762 17184 70768 17196
rect 69983 17156 70768 17184
rect 69983 17153 69995 17156
rect 69937 17147 69995 17153
rect 70762 17144 70768 17156
rect 70820 17144 70826 17196
rect 73816 17193 73844 17224
rect 87598 17212 87604 17224
rect 87656 17212 87662 17264
rect 73801 17187 73859 17193
rect 73801 17153 73813 17187
rect 73847 17153 73859 17187
rect 88245 17187 88303 17193
rect 88245 17184 88257 17187
rect 73801 17147 73859 17153
rect 84166 17156 88257 17184
rect 70394 17116 70400 17128
rect 69768 17088 70400 17116
rect 70394 17076 70400 17088
rect 70452 17076 70458 17128
rect 70578 17076 70584 17128
rect 70636 17116 70642 17128
rect 71041 17119 71099 17125
rect 71041 17116 71053 17119
rect 70636 17088 71053 17116
rect 70636 17076 70642 17088
rect 71041 17085 71053 17088
rect 71087 17116 71099 17119
rect 71314 17116 71320 17128
rect 71087 17088 71320 17116
rect 71087 17085 71099 17088
rect 71041 17079 71099 17085
rect 71314 17076 71320 17088
rect 71372 17076 71378 17128
rect 84166 17116 84194 17156
rect 88245 17153 88257 17156
rect 88291 17153 88303 17187
rect 88245 17147 88303 17153
rect 73632 17088 84194 17116
rect 73632 17057 73660 17088
rect 73617 17051 73675 17057
rect 70964 17020 71268 17048
rect 70964 16980 70992 17020
rect 68940 16952 70992 16980
rect 71240 16980 71268 17020
rect 73617 17017 73629 17051
rect 73663 17017 73675 17051
rect 87046 17048 87052 17060
rect 73617 17011 73675 17017
rect 80026 17020 87052 17048
rect 80026 16980 80054 17020
rect 87046 17008 87052 17020
rect 87104 17008 87110 17060
rect 88058 17048 88064 17060
rect 88019 17020 88064 17048
rect 88058 17008 88064 17020
rect 88116 17008 88122 17060
rect 71240 16952 80054 16980
rect 65567 16949 65579 16952
rect 65521 16943 65579 16949
rect 1104 16890 88872 16912
rect 1104 16838 11924 16890
rect 11976 16838 11988 16890
rect 12040 16838 12052 16890
rect 12104 16838 12116 16890
rect 12168 16838 12180 16890
rect 12232 16838 33872 16890
rect 33924 16838 33936 16890
rect 33988 16838 34000 16890
rect 34052 16838 34064 16890
rect 34116 16838 34128 16890
rect 34180 16838 55820 16890
rect 55872 16838 55884 16890
rect 55936 16838 55948 16890
rect 56000 16838 56012 16890
rect 56064 16838 56076 16890
rect 56128 16838 77768 16890
rect 77820 16838 77832 16890
rect 77884 16838 77896 16890
rect 77948 16838 77960 16890
rect 78012 16838 78024 16890
rect 78076 16838 88872 16890
rect 1104 16816 88872 16838
rect 20070 16776 20076 16788
rect 20031 16748 20076 16776
rect 20070 16736 20076 16748
rect 20128 16736 20134 16788
rect 21082 16736 21088 16788
rect 21140 16776 21146 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 21140 16748 21189 16776
rect 21140 16736 21146 16748
rect 21177 16745 21189 16748
rect 21223 16745 21235 16779
rect 21177 16739 21235 16745
rect 21634 16736 21640 16788
rect 21692 16776 21698 16788
rect 61378 16776 61384 16788
rect 21692 16748 61384 16776
rect 21692 16736 21698 16748
rect 61378 16736 61384 16748
rect 61436 16736 61442 16788
rect 61562 16736 61568 16788
rect 61620 16776 61626 16788
rect 62301 16779 62359 16785
rect 62301 16776 62313 16779
rect 61620 16748 62313 16776
rect 61620 16736 61626 16748
rect 62301 16745 62313 16748
rect 62347 16745 62359 16779
rect 62301 16739 62359 16745
rect 62390 16736 62396 16788
rect 62448 16776 62454 16788
rect 63494 16776 63500 16788
rect 62448 16748 63500 16776
rect 62448 16736 62454 16748
rect 63494 16736 63500 16748
rect 63552 16736 63558 16788
rect 64322 16736 64328 16788
rect 64380 16776 64386 16788
rect 64693 16779 64751 16785
rect 64693 16776 64705 16779
rect 64380 16748 64705 16776
rect 64380 16736 64386 16748
rect 64693 16745 64705 16748
rect 64739 16745 64751 16779
rect 64693 16739 64751 16745
rect 65628 16748 67634 16776
rect 28629 16711 28687 16717
rect 28629 16677 28641 16711
rect 28675 16708 28687 16711
rect 28718 16708 28724 16720
rect 28675 16680 28724 16708
rect 28675 16677 28687 16680
rect 28629 16671 28687 16677
rect 28718 16668 28724 16680
rect 28776 16668 28782 16720
rect 32766 16668 32772 16720
rect 32824 16708 32830 16720
rect 36446 16708 36452 16720
rect 32824 16680 36452 16708
rect 32824 16668 32830 16680
rect 36446 16668 36452 16680
rect 36504 16668 36510 16720
rect 36722 16708 36728 16720
rect 36556 16680 36728 16708
rect 20901 16643 20959 16649
rect 20456 16612 20760 16640
rect 1581 16575 1639 16581
rect 1581 16541 1593 16575
rect 1627 16572 1639 16575
rect 2958 16572 2964 16584
rect 1627 16544 2964 16572
rect 1627 16541 1639 16544
rect 1581 16535 1639 16541
rect 2958 16532 2964 16544
rect 3016 16532 3022 16584
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16572 20315 16575
rect 20456 16572 20484 16612
rect 20303 16544 20484 16572
rect 20303 16541 20315 16544
rect 20257 16535 20315 16541
rect 20530 16532 20536 16584
rect 20588 16572 20594 16584
rect 20732 16572 20760 16612
rect 20901 16609 20913 16643
rect 20947 16640 20959 16643
rect 20947 16612 21680 16640
rect 20947 16609 20959 16612
rect 20901 16603 20959 16609
rect 21652 16584 21680 16612
rect 25774 16600 25780 16652
rect 25832 16640 25838 16652
rect 26053 16643 26111 16649
rect 26053 16640 26065 16643
rect 25832 16612 26065 16640
rect 25832 16600 25838 16612
rect 26053 16609 26065 16612
rect 26099 16609 26111 16643
rect 26053 16603 26111 16609
rect 28166 16600 28172 16652
rect 28224 16640 28230 16652
rect 28261 16643 28319 16649
rect 28261 16640 28273 16643
rect 28224 16612 28273 16640
rect 28224 16600 28230 16612
rect 28261 16609 28273 16612
rect 28307 16609 28319 16643
rect 28261 16603 28319 16609
rect 32858 16600 32864 16652
rect 32916 16640 32922 16652
rect 33597 16643 33655 16649
rect 33597 16640 33609 16643
rect 32916 16612 33609 16640
rect 32916 16600 32922 16612
rect 33597 16609 33609 16612
rect 33643 16609 33655 16643
rect 33597 16603 33655 16609
rect 33689 16643 33747 16649
rect 33689 16609 33701 16643
rect 33735 16609 33747 16643
rect 33689 16603 33747 16609
rect 21358 16572 21364 16584
rect 20588 16544 20633 16572
rect 20732 16544 21364 16572
rect 20588 16532 20594 16544
rect 21358 16532 21364 16544
rect 21416 16532 21422 16584
rect 21634 16572 21640 16584
rect 21595 16544 21640 16572
rect 21634 16532 21640 16544
rect 21692 16532 21698 16584
rect 25685 16575 25743 16581
rect 25685 16541 25697 16575
rect 25731 16572 25743 16575
rect 25958 16572 25964 16584
rect 25731 16544 25964 16572
rect 25731 16541 25743 16544
rect 25685 16535 25743 16541
rect 25958 16532 25964 16544
rect 26016 16532 26022 16584
rect 26326 16581 26332 16584
rect 26320 16535 26332 16581
rect 26326 16532 26332 16535
rect 26384 16532 26390 16584
rect 28442 16572 28448 16584
rect 28403 16544 28448 16572
rect 28442 16532 28448 16544
rect 28500 16532 28506 16584
rect 30834 16572 30840 16584
rect 30795 16544 30840 16572
rect 30834 16532 30840 16544
rect 30892 16532 30898 16584
rect 31110 16532 31116 16584
rect 31168 16572 31174 16584
rect 31205 16575 31263 16581
rect 31205 16572 31217 16575
rect 31168 16544 31217 16572
rect 31168 16532 31174 16544
rect 31205 16541 31217 16544
rect 31251 16541 31263 16575
rect 31205 16535 31263 16541
rect 33318 16532 33324 16584
rect 33376 16572 33382 16584
rect 33704 16572 33732 16603
rect 33778 16600 33784 16652
rect 33836 16640 33842 16652
rect 36354 16640 36360 16652
rect 33836 16612 35940 16640
rect 36315 16612 36360 16640
rect 33836 16600 33842 16612
rect 35912 16584 35940 16612
rect 36354 16600 36360 16612
rect 36412 16600 36418 16652
rect 36556 16649 36584 16680
rect 36722 16668 36728 16680
rect 36780 16708 36786 16720
rect 40037 16711 40095 16717
rect 36780 16680 39988 16708
rect 36780 16668 36786 16680
rect 36541 16643 36599 16649
rect 36541 16609 36553 16643
rect 36587 16609 36599 16643
rect 36541 16603 36599 16609
rect 36814 16600 36820 16652
rect 36872 16640 36878 16652
rect 38746 16640 38752 16652
rect 36872 16612 38608 16640
rect 36872 16600 36878 16612
rect 35345 16575 35403 16581
rect 35345 16572 35357 16575
rect 33376 16544 33732 16572
rect 34716 16544 35357 16572
rect 33376 16532 33382 16544
rect 34716 16516 34744 16544
rect 35345 16541 35357 16544
rect 35391 16541 35403 16575
rect 35345 16535 35403 16541
rect 35894 16532 35900 16584
rect 35952 16532 35958 16584
rect 36265 16575 36323 16581
rect 36265 16541 36277 16575
rect 36311 16572 36323 16575
rect 38194 16572 38200 16584
rect 36311 16544 38200 16572
rect 36311 16541 36323 16544
rect 36265 16535 36323 16541
rect 38194 16532 38200 16544
rect 38252 16532 38258 16584
rect 38580 16581 38608 16612
rect 38672 16612 38752 16640
rect 38565 16575 38623 16581
rect 38565 16541 38577 16575
rect 38611 16541 38623 16575
rect 38565 16535 38623 16541
rect 20441 16507 20499 16513
rect 20441 16473 20453 16507
rect 20487 16504 20499 16507
rect 21545 16507 21603 16513
rect 21545 16504 21557 16507
rect 20487 16476 21557 16504
rect 20487 16473 20499 16476
rect 20441 16467 20499 16473
rect 21545 16473 21557 16476
rect 21591 16504 21603 16507
rect 26142 16504 26148 16516
rect 21591 16476 26148 16504
rect 21591 16473 21603 16476
rect 21545 16467 21603 16473
rect 26142 16464 26148 16476
rect 26200 16464 26206 16516
rect 28626 16504 28632 16516
rect 26436 16476 28632 16504
rect 1394 16436 1400 16448
rect 1355 16408 1400 16436
rect 1394 16396 1400 16408
rect 1452 16396 1458 16448
rect 25314 16396 25320 16448
rect 25372 16436 25378 16448
rect 25501 16439 25559 16445
rect 25501 16436 25513 16439
rect 25372 16408 25513 16436
rect 25372 16396 25378 16408
rect 25501 16405 25513 16408
rect 25547 16405 25559 16439
rect 25501 16399 25559 16405
rect 25590 16396 25596 16448
rect 25648 16436 25654 16448
rect 26436 16436 26464 16476
rect 28626 16464 28632 16476
rect 28684 16464 28690 16516
rect 31478 16513 31484 16516
rect 31472 16504 31484 16513
rect 31439 16476 31484 16504
rect 31472 16467 31484 16476
rect 31478 16464 31484 16467
rect 31536 16464 31542 16516
rect 32858 16504 32864 16516
rect 31726 16476 32864 16504
rect 27430 16436 27436 16448
rect 25648 16408 26464 16436
rect 27391 16408 27436 16436
rect 25648 16396 25654 16408
rect 27430 16396 27436 16408
rect 27488 16396 27494 16448
rect 29178 16396 29184 16448
rect 29236 16436 29242 16448
rect 29730 16436 29736 16448
rect 29236 16408 29736 16436
rect 29236 16396 29242 16408
rect 29730 16396 29736 16408
rect 29788 16396 29794 16448
rect 30650 16436 30656 16448
rect 30611 16408 30656 16436
rect 30650 16396 30656 16408
rect 30708 16396 30714 16448
rect 30742 16396 30748 16448
rect 30800 16436 30806 16448
rect 31726 16436 31754 16476
rect 32858 16464 32864 16476
rect 32916 16464 32922 16516
rect 33505 16507 33563 16513
rect 33505 16473 33517 16507
rect 33551 16504 33563 16507
rect 34698 16504 34704 16516
rect 33551 16476 34704 16504
rect 33551 16473 33563 16476
rect 33505 16467 33563 16473
rect 34698 16464 34704 16476
rect 34756 16464 34762 16516
rect 35912 16504 35940 16532
rect 38013 16507 38071 16513
rect 38013 16504 38025 16507
rect 35912 16476 38025 16504
rect 38013 16473 38025 16476
rect 38059 16504 38071 16507
rect 38672 16504 38700 16612
rect 38746 16600 38752 16612
rect 38804 16600 38810 16652
rect 39960 16640 39988 16680
rect 40037 16677 40049 16711
rect 40083 16708 40095 16711
rect 40126 16708 40132 16720
rect 40083 16680 40132 16708
rect 40083 16677 40095 16680
rect 40037 16671 40095 16677
rect 40126 16668 40132 16680
rect 40184 16668 40190 16720
rect 40310 16668 40316 16720
rect 40368 16708 40374 16720
rect 41690 16708 41696 16720
rect 40368 16680 41696 16708
rect 40368 16668 40374 16680
rect 41690 16668 41696 16680
rect 41748 16668 41754 16720
rect 42978 16668 42984 16720
rect 43036 16708 43042 16720
rect 45922 16708 45928 16720
rect 43036 16680 45928 16708
rect 43036 16668 43042 16680
rect 45922 16668 45928 16680
rect 45980 16668 45986 16720
rect 46569 16711 46627 16717
rect 46569 16677 46581 16711
rect 46615 16708 46627 16711
rect 46934 16708 46940 16720
rect 46615 16680 46940 16708
rect 46615 16677 46627 16680
rect 46569 16671 46627 16677
rect 46934 16668 46940 16680
rect 46992 16668 46998 16720
rect 47762 16708 47768 16720
rect 47723 16680 47768 16708
rect 47762 16668 47768 16680
rect 47820 16668 47826 16720
rect 47854 16668 47860 16720
rect 47912 16708 47918 16720
rect 50062 16708 50068 16720
rect 47912 16680 50068 16708
rect 47912 16668 47918 16680
rect 50062 16668 50068 16680
rect 50120 16668 50126 16720
rect 51258 16668 51264 16720
rect 51316 16708 51322 16720
rect 52822 16708 52828 16720
rect 51316 16680 52828 16708
rect 51316 16668 51322 16680
rect 52822 16668 52828 16680
rect 52880 16668 52886 16720
rect 52917 16711 52975 16717
rect 52917 16677 52929 16711
rect 52963 16708 52975 16711
rect 55122 16708 55128 16720
rect 52963 16680 55128 16708
rect 52963 16677 52975 16680
rect 52917 16671 52975 16677
rect 55122 16668 55128 16680
rect 55180 16668 55186 16720
rect 57793 16711 57851 16717
rect 57793 16677 57805 16711
rect 57839 16708 57851 16711
rect 58710 16708 58716 16720
rect 57839 16680 58716 16708
rect 57839 16677 57851 16680
rect 57793 16671 57851 16677
rect 58710 16668 58716 16680
rect 58768 16668 58774 16720
rect 59262 16668 59268 16720
rect 59320 16708 59326 16720
rect 62022 16708 62028 16720
rect 59320 16680 62028 16708
rect 59320 16668 59326 16680
rect 62022 16668 62028 16680
rect 62080 16668 62086 16720
rect 63034 16668 63040 16720
rect 63092 16708 63098 16720
rect 64138 16708 64144 16720
rect 63092 16680 64144 16708
rect 63092 16668 63098 16680
rect 64138 16668 64144 16680
rect 64196 16708 64202 16720
rect 64782 16708 64788 16720
rect 64196 16680 64788 16708
rect 64196 16668 64202 16680
rect 64782 16668 64788 16680
rect 64840 16668 64846 16720
rect 47026 16640 47032 16652
rect 39960 16612 41736 16640
rect 41708 16584 41736 16612
rect 44100 16612 47032 16640
rect 40218 16572 40224 16584
rect 40179 16544 40224 16572
rect 40218 16532 40224 16544
rect 40276 16532 40282 16584
rect 41506 16572 41512 16584
rect 41467 16544 41512 16572
rect 41506 16532 41512 16544
rect 41564 16532 41570 16584
rect 41690 16532 41696 16584
rect 41748 16532 41754 16584
rect 41874 16532 41880 16584
rect 41932 16572 41938 16584
rect 42702 16572 42708 16584
rect 41932 16544 42708 16572
rect 41932 16532 41938 16544
rect 42702 16532 42708 16544
rect 42760 16532 42766 16584
rect 44100 16581 44128 16612
rect 47026 16600 47032 16612
rect 47084 16640 47090 16652
rect 48222 16640 48228 16652
rect 47084 16612 48228 16640
rect 47084 16600 47090 16612
rect 48222 16600 48228 16612
rect 48280 16640 48286 16652
rect 48280 16600 48314 16640
rect 49786 16600 49792 16652
rect 49844 16640 49850 16652
rect 50157 16643 50215 16649
rect 50157 16640 50169 16643
rect 49844 16612 50169 16640
rect 49844 16600 49850 16612
rect 50157 16609 50169 16612
rect 50203 16609 50215 16643
rect 50157 16603 50215 16609
rect 51166 16600 51172 16652
rect 51224 16640 51230 16652
rect 53466 16640 53472 16652
rect 51224 16612 53472 16640
rect 51224 16600 51230 16612
rect 53466 16600 53472 16612
rect 53524 16600 53530 16652
rect 54297 16643 54355 16649
rect 54297 16640 54309 16643
rect 53668 16612 54309 16640
rect 43809 16575 43867 16581
rect 43809 16541 43821 16575
rect 43855 16541 43867 16575
rect 43809 16535 43867 16541
rect 44085 16575 44143 16581
rect 44085 16541 44097 16575
rect 44131 16541 44143 16575
rect 46750 16572 46756 16584
rect 44085 16535 44143 16541
rect 44744 16544 46756 16572
rect 42122 16507 42180 16513
rect 42122 16504 42134 16507
rect 38059 16476 38700 16504
rect 41340 16476 42134 16504
rect 38059 16473 38071 16476
rect 38013 16467 38071 16473
rect 30800 16408 31754 16436
rect 32585 16439 32643 16445
rect 30800 16396 30806 16408
rect 32585 16405 32597 16439
rect 32631 16436 32643 16439
rect 32674 16436 32680 16448
rect 32631 16408 32680 16436
rect 32631 16405 32643 16408
rect 32585 16399 32643 16405
rect 32674 16396 32680 16408
rect 32732 16396 32738 16448
rect 33134 16436 33140 16448
rect 33095 16408 33140 16436
rect 33134 16396 33140 16408
rect 33192 16396 33198 16448
rect 35437 16439 35495 16445
rect 35437 16405 35449 16439
rect 35483 16436 35495 16439
rect 35526 16436 35532 16448
rect 35483 16408 35532 16436
rect 35483 16405 35495 16408
rect 35437 16399 35495 16405
rect 35526 16396 35532 16408
rect 35584 16396 35590 16448
rect 35897 16439 35955 16445
rect 35897 16405 35909 16439
rect 35943 16436 35955 16439
rect 35986 16436 35992 16448
rect 35943 16408 35992 16436
rect 35943 16405 35955 16408
rect 35897 16399 35955 16405
rect 35986 16396 35992 16408
rect 36044 16396 36050 16448
rect 37550 16396 37556 16448
rect 37608 16436 37614 16448
rect 38105 16439 38163 16445
rect 38105 16436 38117 16439
rect 37608 16408 38117 16436
rect 37608 16396 37614 16408
rect 38105 16405 38117 16408
rect 38151 16405 38163 16439
rect 38654 16436 38660 16448
rect 38615 16408 38660 16436
rect 38105 16399 38163 16405
rect 38654 16396 38660 16408
rect 38712 16396 38718 16448
rect 41340 16445 41368 16476
rect 42122 16473 42134 16476
rect 42168 16473 42180 16507
rect 43824 16504 43852 16535
rect 44744 16516 44772 16544
rect 46750 16532 46756 16544
rect 46808 16532 46814 16584
rect 46842 16532 46848 16584
rect 46900 16572 46906 16584
rect 47210 16572 47216 16584
rect 46900 16544 46945 16572
rect 47171 16544 47216 16572
rect 46900 16532 46906 16544
rect 47210 16532 47216 16544
rect 47268 16532 47274 16584
rect 47394 16572 47400 16584
rect 47355 16544 47400 16572
rect 47394 16532 47400 16544
rect 47452 16532 47458 16584
rect 47578 16572 47584 16584
rect 47636 16581 47642 16584
rect 47544 16544 47584 16572
rect 47578 16532 47584 16544
rect 47636 16535 47644 16581
rect 48286 16572 48314 16600
rect 50246 16572 50252 16584
rect 48286 16544 50252 16572
rect 47636 16532 47642 16535
rect 50246 16532 50252 16544
rect 50304 16532 50310 16584
rect 50424 16575 50482 16581
rect 50424 16541 50436 16575
rect 50470 16572 50482 16575
rect 51350 16572 51356 16584
rect 50470 16544 51356 16572
rect 50470 16541 50482 16544
rect 50424 16535 50482 16541
rect 51350 16532 51356 16544
rect 51408 16532 51414 16584
rect 52362 16572 52368 16584
rect 52323 16544 52368 16572
rect 52362 16532 52368 16544
rect 52420 16532 52426 16584
rect 52546 16572 52552 16584
rect 52507 16544 52552 16572
rect 52546 16532 52552 16544
rect 52604 16532 52610 16584
rect 52730 16532 52736 16584
rect 52788 16581 52794 16584
rect 52788 16572 52796 16581
rect 53374 16572 53380 16584
rect 52788 16544 52833 16572
rect 53335 16544 53380 16572
rect 52788 16535 52796 16544
rect 52788 16532 52794 16535
rect 53374 16532 53380 16544
rect 53432 16532 53438 16584
rect 53561 16575 53619 16581
rect 53561 16541 53573 16575
rect 53607 16572 53619 16575
rect 53668 16572 53696 16612
rect 54297 16609 54309 16612
rect 54343 16609 54355 16643
rect 54297 16603 54355 16609
rect 54404 16612 55168 16640
rect 53607 16544 53696 16572
rect 53745 16575 53803 16581
rect 53607 16541 53619 16544
rect 53561 16535 53619 16541
rect 53745 16541 53757 16575
rect 53791 16541 53803 16575
rect 53745 16535 53803 16541
rect 44726 16504 44732 16516
rect 42122 16467 42180 16473
rect 43272 16476 43760 16504
rect 43824 16476 44732 16504
rect 41325 16439 41383 16445
rect 41325 16405 41337 16439
rect 41371 16405 41383 16439
rect 41325 16399 41383 16405
rect 41782 16396 41788 16448
rect 41840 16436 41846 16448
rect 43162 16436 43168 16448
rect 41840 16408 43168 16436
rect 41840 16396 41846 16408
rect 43162 16396 43168 16408
rect 43220 16396 43226 16448
rect 43272 16445 43300 16476
rect 43257 16439 43315 16445
rect 43257 16405 43269 16439
rect 43303 16405 43315 16439
rect 43257 16399 43315 16405
rect 43346 16396 43352 16448
rect 43404 16436 43410 16448
rect 43625 16439 43683 16445
rect 43625 16436 43637 16439
rect 43404 16408 43637 16436
rect 43404 16396 43410 16408
rect 43625 16405 43637 16408
rect 43671 16405 43683 16439
rect 43732 16436 43760 16476
rect 44726 16464 44732 16476
rect 44784 16464 44790 16516
rect 46569 16507 46627 16513
rect 46569 16473 46581 16507
rect 46615 16504 46627 16507
rect 47118 16504 47124 16516
rect 46615 16476 47124 16504
rect 46615 16473 46627 16476
rect 46569 16467 46627 16473
rect 47118 16464 47124 16476
rect 47176 16464 47182 16516
rect 47302 16464 47308 16516
rect 47360 16504 47366 16516
rect 47489 16507 47547 16513
rect 47489 16504 47501 16507
rect 47360 16476 47501 16504
rect 47360 16464 47366 16476
rect 47489 16473 47501 16476
rect 47535 16504 47547 16507
rect 50890 16504 50896 16516
rect 47535 16476 50896 16504
rect 47535 16473 47547 16476
rect 47489 16467 47547 16473
rect 50890 16464 50896 16476
rect 50948 16464 50954 16516
rect 50982 16464 50988 16516
rect 51040 16504 51046 16516
rect 51074 16504 51080 16516
rect 51040 16476 51080 16504
rect 51040 16464 51046 16476
rect 51074 16464 51080 16476
rect 51132 16464 51138 16516
rect 51994 16504 52000 16516
rect 51552 16476 52000 16504
rect 43993 16439 44051 16445
rect 43993 16436 44005 16439
rect 43732 16408 44005 16436
rect 43625 16399 43683 16405
rect 43993 16405 44005 16408
rect 44039 16405 44051 16439
rect 43993 16399 44051 16405
rect 44818 16396 44824 16448
rect 44876 16436 44882 16448
rect 46658 16436 46664 16448
rect 44876 16408 46664 16436
rect 44876 16396 44882 16408
rect 46658 16396 46664 16408
rect 46716 16396 46722 16448
rect 46753 16439 46811 16445
rect 46753 16405 46765 16439
rect 46799 16436 46811 16439
rect 47762 16436 47768 16448
rect 46799 16408 47768 16436
rect 46799 16405 46811 16408
rect 46753 16399 46811 16405
rect 47762 16396 47768 16408
rect 47820 16396 47826 16448
rect 48222 16396 48228 16448
rect 48280 16436 48286 16448
rect 50246 16436 50252 16448
rect 48280 16408 50252 16436
rect 48280 16396 48286 16408
rect 50246 16396 50252 16408
rect 50304 16396 50310 16448
rect 50338 16396 50344 16448
rect 50396 16436 50402 16448
rect 51442 16436 51448 16448
rect 50396 16408 51448 16436
rect 50396 16396 50402 16408
rect 51442 16396 51448 16408
rect 51500 16396 51506 16448
rect 51552 16445 51580 16476
rect 51994 16464 52000 16476
rect 52052 16464 52058 16516
rect 52454 16464 52460 16516
rect 52512 16504 52518 16516
rect 52641 16507 52699 16513
rect 52641 16504 52653 16507
rect 52512 16476 52653 16504
rect 52512 16464 52518 16476
rect 52641 16473 52653 16476
rect 52687 16473 52699 16507
rect 52641 16467 52699 16473
rect 53098 16464 53104 16516
rect 53156 16504 53162 16516
rect 53653 16507 53711 16513
rect 53653 16504 53665 16507
rect 53156 16476 53665 16504
rect 53156 16464 53162 16476
rect 53653 16473 53665 16476
rect 53699 16473 53711 16507
rect 53653 16467 53711 16473
rect 51537 16439 51595 16445
rect 51537 16405 51549 16439
rect 51583 16405 51595 16439
rect 51537 16399 51595 16405
rect 51626 16396 51632 16448
rect 51684 16436 51690 16448
rect 53760 16436 53788 16535
rect 53926 16532 53932 16584
rect 53984 16572 53990 16584
rect 54404 16572 54432 16612
rect 53984 16544 54432 16572
rect 54481 16575 54539 16581
rect 53984 16532 53990 16544
rect 54481 16541 54493 16575
rect 54527 16541 54539 16575
rect 54754 16572 54760 16584
rect 54715 16544 54760 16572
rect 54481 16535 54539 16541
rect 54110 16464 54116 16516
rect 54168 16504 54174 16516
rect 54386 16504 54392 16516
rect 54168 16476 54392 16504
rect 54168 16464 54174 16476
rect 54386 16464 54392 16476
rect 54444 16504 54450 16516
rect 54496 16504 54524 16535
rect 54754 16532 54760 16544
rect 54812 16532 54818 16584
rect 55140 16572 55168 16612
rect 55214 16600 55220 16652
rect 55272 16640 55278 16652
rect 55309 16643 55367 16649
rect 55309 16640 55321 16643
rect 55272 16612 55321 16640
rect 55272 16600 55278 16612
rect 55309 16609 55321 16612
rect 55355 16609 55367 16643
rect 58894 16640 58900 16652
rect 55309 16603 55367 16609
rect 56336 16612 58900 16640
rect 56336 16572 56364 16612
rect 58894 16600 58900 16612
rect 58952 16600 58958 16652
rect 59357 16643 59415 16649
rect 59357 16609 59369 16643
rect 59403 16640 59415 16643
rect 59906 16640 59912 16652
rect 59403 16612 59912 16640
rect 59403 16609 59415 16612
rect 59357 16603 59415 16609
rect 59906 16600 59912 16612
rect 59964 16600 59970 16652
rect 65242 16640 65248 16652
rect 64892 16612 65248 16640
rect 55140 16544 56364 16572
rect 56502 16532 56508 16584
rect 56560 16572 56566 16584
rect 57241 16575 57299 16581
rect 57241 16572 57253 16575
rect 56560 16544 57253 16572
rect 56560 16532 56566 16544
rect 57241 16541 57253 16544
rect 57287 16541 57299 16575
rect 58069 16575 58127 16581
rect 58069 16572 58081 16575
rect 57241 16535 57299 16541
rect 57348 16544 58081 16572
rect 54444 16476 54524 16504
rect 54665 16507 54723 16513
rect 54444 16464 54450 16476
rect 54665 16473 54677 16507
rect 54711 16504 54723 16507
rect 55306 16504 55312 16516
rect 54711 16476 55312 16504
rect 54711 16473 54723 16476
rect 54665 16467 54723 16473
rect 55306 16464 55312 16476
rect 55364 16464 55370 16516
rect 55576 16507 55634 16513
rect 55576 16473 55588 16507
rect 55622 16504 55634 16507
rect 56594 16504 56600 16516
rect 55622 16476 56600 16504
rect 55622 16473 55634 16476
rect 55576 16467 55634 16473
rect 56594 16464 56600 16476
rect 56652 16464 56658 16516
rect 56870 16464 56876 16516
rect 56928 16504 56934 16516
rect 57348 16504 57376 16544
rect 58069 16541 58081 16544
rect 58115 16541 58127 16575
rect 58621 16575 58679 16581
rect 58621 16572 58633 16575
rect 58069 16535 58127 16541
rect 58176 16544 58633 16572
rect 56928 16476 57376 16504
rect 57793 16507 57851 16513
rect 56928 16464 56934 16476
rect 57793 16473 57805 16507
rect 57839 16504 57851 16507
rect 57882 16504 57888 16516
rect 57839 16476 57888 16504
rect 57839 16473 57851 16476
rect 57793 16467 57851 16473
rect 57882 16464 57888 16476
rect 57940 16464 57946 16516
rect 58176 16504 58204 16544
rect 58621 16541 58633 16544
rect 58667 16541 58679 16575
rect 58621 16535 58679 16541
rect 58713 16575 58771 16581
rect 58713 16541 58725 16575
rect 58759 16541 58771 16575
rect 58713 16535 58771 16541
rect 60553 16575 60611 16581
rect 60553 16541 60565 16575
rect 60599 16572 60611 16575
rect 60826 16572 60832 16584
rect 60599 16544 60832 16572
rect 60599 16541 60611 16544
rect 60553 16535 60611 16541
rect 58434 16504 58440 16516
rect 57992 16476 58204 16504
rect 58395 16476 58440 16504
rect 51684 16408 53788 16436
rect 53929 16439 53987 16445
rect 51684 16396 51690 16408
rect 53929 16405 53941 16439
rect 53975 16436 53987 16439
rect 54294 16436 54300 16448
rect 53975 16408 54300 16436
rect 53975 16405 53987 16408
rect 53929 16399 53987 16405
rect 54294 16396 54300 16408
rect 54352 16396 54358 16448
rect 56410 16396 56416 16448
rect 56468 16436 56474 16448
rect 56689 16439 56747 16445
rect 56689 16436 56701 16439
rect 56468 16408 56701 16436
rect 56468 16396 56474 16408
rect 56689 16405 56701 16408
rect 56735 16405 56747 16439
rect 56689 16399 56747 16405
rect 56778 16396 56784 16448
rect 56836 16436 56842 16448
rect 57057 16439 57115 16445
rect 57057 16436 57069 16439
rect 56836 16408 57069 16436
rect 56836 16396 56842 16408
rect 57057 16405 57069 16408
rect 57103 16405 57115 16439
rect 57057 16399 57115 16405
rect 57330 16396 57336 16448
rect 57388 16436 57394 16448
rect 57992 16445 58020 16476
rect 58434 16464 58440 16476
rect 58492 16464 58498 16516
rect 57977 16439 58035 16445
rect 57977 16436 57989 16439
rect 57388 16408 57989 16436
rect 57388 16396 57394 16408
rect 57977 16405 57989 16408
rect 58023 16405 58035 16439
rect 58526 16436 58532 16448
rect 58584 16445 58590 16448
rect 58493 16408 58532 16436
rect 57977 16399 58035 16405
rect 58526 16396 58532 16408
rect 58584 16399 58593 16445
rect 58728 16436 58756 16535
rect 60826 16532 60832 16544
rect 60884 16572 60890 16584
rect 61010 16572 61016 16584
rect 60884 16544 61016 16572
rect 60884 16532 60890 16544
rect 61010 16532 61016 16544
rect 61068 16532 61074 16584
rect 61102 16532 61108 16584
rect 61160 16572 61166 16584
rect 61381 16575 61439 16581
rect 61160 16544 61253 16572
rect 61160 16532 61166 16544
rect 61381 16541 61393 16575
rect 61427 16572 61439 16575
rect 62485 16575 62543 16581
rect 61427 16544 61608 16572
rect 61427 16541 61439 16544
rect 61381 16535 61439 16541
rect 59078 16464 59084 16516
rect 59136 16504 59142 16516
rect 59173 16507 59231 16513
rect 59173 16504 59185 16507
rect 59136 16476 59185 16504
rect 59136 16464 59142 16476
rect 59173 16473 59185 16476
rect 59219 16473 59231 16507
rect 59173 16467 59231 16473
rect 59262 16464 59268 16516
rect 59320 16504 59326 16516
rect 59817 16507 59875 16513
rect 59817 16504 59829 16507
rect 59320 16476 59829 16504
rect 59320 16464 59326 16476
rect 59817 16473 59829 16476
rect 59863 16473 59875 16507
rect 59817 16467 59875 16473
rect 60001 16507 60059 16513
rect 60001 16473 60013 16507
rect 60047 16504 60059 16507
rect 60090 16504 60096 16516
rect 60047 16476 60096 16504
rect 60047 16473 60059 16476
rect 60001 16467 60059 16473
rect 60090 16464 60096 16476
rect 60148 16464 60154 16516
rect 60734 16464 60740 16516
rect 60792 16504 60798 16516
rect 61120 16504 61148 16532
rect 60792 16476 61148 16504
rect 60792 16464 60798 16476
rect 61194 16464 61200 16516
rect 61252 16504 61258 16516
rect 61580 16504 61608 16544
rect 62485 16541 62497 16575
rect 62531 16572 62543 16575
rect 62574 16572 62580 16584
rect 62531 16544 62580 16572
rect 62531 16541 62543 16544
rect 62485 16535 62543 16541
rect 62574 16532 62580 16544
rect 62632 16532 62638 16584
rect 62758 16572 62764 16584
rect 62719 16544 62764 16572
rect 62758 16532 62764 16544
rect 62816 16532 62822 16584
rect 64892 16581 64920 16612
rect 65242 16600 65248 16612
rect 65300 16600 65306 16652
rect 65518 16600 65524 16652
rect 65576 16640 65582 16652
rect 65628 16649 65656 16748
rect 65613 16643 65671 16649
rect 65613 16640 65625 16643
rect 65576 16612 65625 16640
rect 65576 16600 65582 16612
rect 65613 16609 65625 16612
rect 65659 16609 65671 16643
rect 67606 16640 67634 16748
rect 68554 16736 68560 16788
rect 68612 16776 68618 16788
rect 87322 16776 87328 16788
rect 68612 16748 87328 16776
rect 68612 16736 68618 16748
rect 87322 16736 87328 16748
rect 87380 16736 87386 16788
rect 69382 16668 69388 16720
rect 69440 16708 69446 16720
rect 77110 16708 77116 16720
rect 69440 16680 77116 16708
rect 69440 16668 69446 16680
rect 77110 16668 77116 16680
rect 77168 16668 77174 16720
rect 68373 16643 68431 16649
rect 68373 16640 68385 16643
rect 67606 16612 68385 16640
rect 65613 16603 65671 16609
rect 68373 16609 68385 16612
rect 68419 16609 68431 16643
rect 71130 16640 71136 16652
rect 71091 16612 71136 16640
rect 68373 16603 68431 16609
rect 63221 16575 63279 16581
rect 63221 16572 63233 16575
rect 62868 16544 63233 16572
rect 61252 16476 61608 16504
rect 61252 16464 61258 16476
rect 60182 16436 60188 16448
rect 58728 16408 60188 16436
rect 58584 16396 58590 16399
rect 60182 16396 60188 16408
rect 60240 16396 60246 16448
rect 60642 16396 60648 16448
rect 60700 16436 60706 16448
rect 61580 16436 61608 16476
rect 61654 16464 61660 16516
rect 61712 16504 61718 16516
rect 62669 16507 62727 16513
rect 62669 16504 62681 16507
rect 61712 16476 62681 16504
rect 61712 16464 61718 16476
rect 62669 16473 62681 16476
rect 62715 16473 62727 16507
rect 62669 16467 62727 16473
rect 62868 16436 62896 16544
rect 63221 16541 63233 16544
rect 63267 16572 63279 16575
rect 63865 16575 63923 16581
rect 63865 16572 63877 16575
rect 63267 16544 63877 16572
rect 63267 16541 63279 16544
rect 63221 16535 63279 16541
rect 63865 16541 63877 16544
rect 63911 16541 63923 16575
rect 63865 16535 63923 16541
rect 64049 16575 64107 16581
rect 64049 16541 64061 16575
rect 64095 16572 64107 16575
rect 64877 16575 64935 16581
rect 64877 16572 64889 16575
rect 64095 16544 64889 16572
rect 64095 16541 64107 16544
rect 64049 16535 64107 16541
rect 64877 16541 64889 16544
rect 64923 16541 64935 16575
rect 64877 16535 64935 16541
rect 65153 16575 65211 16581
rect 65153 16541 65165 16575
rect 65199 16541 65211 16575
rect 65153 16535 65211 16541
rect 63126 16464 63132 16516
rect 63184 16504 63190 16516
rect 64064 16504 64092 16535
rect 63184 16476 64092 16504
rect 65168 16504 65196 16535
rect 65334 16532 65340 16584
rect 65392 16572 65398 16584
rect 65869 16575 65927 16581
rect 65869 16572 65881 16575
rect 65392 16544 65881 16572
rect 65392 16532 65398 16544
rect 65869 16541 65881 16544
rect 65915 16541 65927 16575
rect 68388 16572 68416 16603
rect 71130 16600 71136 16612
rect 71188 16600 71194 16652
rect 71501 16643 71559 16649
rect 71501 16609 71513 16643
rect 71547 16640 71559 16643
rect 73062 16640 73068 16652
rect 71547 16612 73068 16640
rect 71547 16609 71559 16612
rect 71501 16603 71559 16609
rect 73062 16600 73068 16612
rect 73120 16600 73126 16652
rect 68922 16572 68928 16584
rect 68388 16544 68928 16572
rect 65869 16535 65927 16541
rect 68922 16532 68928 16544
rect 68980 16532 68986 16584
rect 70305 16575 70363 16581
rect 70305 16541 70317 16575
rect 70351 16572 70363 16575
rect 70762 16572 70768 16584
rect 70351 16544 70768 16572
rect 70351 16541 70363 16544
rect 70305 16535 70363 16541
rect 70762 16532 70768 16544
rect 70820 16532 70826 16584
rect 71314 16572 71320 16584
rect 71275 16544 71320 16572
rect 71314 16532 71320 16544
rect 71372 16532 71378 16584
rect 87874 16532 87880 16584
rect 87932 16572 87938 16584
rect 88245 16575 88303 16581
rect 88245 16572 88257 16575
rect 87932 16544 88257 16572
rect 87932 16532 87938 16544
rect 88245 16541 88257 16544
rect 88291 16541 88303 16575
rect 88245 16535 88303 16541
rect 68646 16513 68652 16516
rect 68640 16504 68652 16513
rect 65168 16476 67634 16504
rect 68607 16476 68652 16504
rect 63184 16464 63190 16476
rect 63310 16436 63316 16448
rect 60700 16408 60745 16436
rect 61580 16408 62896 16436
rect 63271 16408 63316 16436
rect 60700 16396 60706 16408
rect 63310 16396 63316 16408
rect 63368 16396 63374 16448
rect 65061 16439 65119 16445
rect 65061 16405 65073 16439
rect 65107 16436 65119 16439
rect 65334 16436 65340 16448
rect 65107 16408 65340 16436
rect 65107 16405 65119 16408
rect 65061 16399 65119 16405
rect 65334 16396 65340 16408
rect 65392 16396 65398 16448
rect 65978 16396 65984 16448
rect 66036 16436 66042 16448
rect 66993 16439 67051 16445
rect 66993 16436 67005 16439
rect 66036 16408 67005 16436
rect 66036 16396 66042 16408
rect 66993 16405 67005 16408
rect 67039 16405 67051 16439
rect 67606 16436 67634 16476
rect 68640 16467 68652 16476
rect 68646 16464 68652 16467
rect 68704 16464 68710 16516
rect 68370 16436 68376 16448
rect 67606 16408 68376 16436
rect 66993 16399 67051 16405
rect 68370 16396 68376 16408
rect 68428 16436 68434 16448
rect 68554 16436 68560 16448
rect 68428 16408 68560 16436
rect 68428 16396 68434 16408
rect 68554 16396 68560 16408
rect 68612 16396 68618 16448
rect 69750 16436 69756 16448
rect 69711 16408 69756 16436
rect 69750 16396 69756 16408
rect 69808 16396 69814 16448
rect 70118 16436 70124 16448
rect 70079 16408 70124 16436
rect 70118 16396 70124 16408
rect 70176 16396 70182 16448
rect 88058 16436 88064 16448
rect 88019 16408 88064 16436
rect 88058 16396 88064 16408
rect 88116 16396 88122 16448
rect 1104 16346 88872 16368
rect 1104 16294 22898 16346
rect 22950 16294 22962 16346
rect 23014 16294 23026 16346
rect 23078 16294 23090 16346
rect 23142 16294 23154 16346
rect 23206 16294 44846 16346
rect 44898 16294 44910 16346
rect 44962 16294 44974 16346
rect 45026 16294 45038 16346
rect 45090 16294 45102 16346
rect 45154 16294 66794 16346
rect 66846 16294 66858 16346
rect 66910 16294 66922 16346
rect 66974 16294 66986 16346
rect 67038 16294 67050 16346
rect 67102 16294 88872 16346
rect 1104 16272 88872 16294
rect 2958 16232 2964 16244
rect 2919 16204 2964 16232
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 20254 16192 20260 16244
rect 20312 16232 20318 16244
rect 21821 16235 21879 16241
rect 21821 16232 21833 16235
rect 20312 16204 21833 16232
rect 20312 16192 20318 16204
rect 21821 16201 21833 16204
rect 21867 16201 21879 16235
rect 21821 16195 21879 16201
rect 22554 16192 22560 16244
rect 22612 16232 22618 16244
rect 24397 16235 24455 16241
rect 24397 16232 24409 16235
rect 22612 16204 24409 16232
rect 22612 16192 22618 16204
rect 24397 16201 24409 16204
rect 24443 16201 24455 16235
rect 24397 16195 24455 16201
rect 24578 16192 24584 16244
rect 24636 16232 24642 16244
rect 25590 16232 25596 16244
rect 24636 16204 25596 16232
rect 24636 16192 24642 16204
rect 25590 16192 25596 16204
rect 25648 16192 25654 16244
rect 26234 16192 26240 16244
rect 26292 16232 26298 16244
rect 30377 16235 30435 16241
rect 30377 16232 30389 16235
rect 26292 16204 30389 16232
rect 26292 16192 26298 16204
rect 30377 16201 30389 16204
rect 30423 16232 30435 16235
rect 30742 16232 30748 16244
rect 30423 16204 30748 16232
rect 30423 16201 30435 16204
rect 30377 16195 30435 16201
rect 30742 16192 30748 16204
rect 30800 16192 30806 16244
rect 31481 16235 31539 16241
rect 31481 16201 31493 16235
rect 31527 16232 31539 16235
rect 34698 16232 34704 16244
rect 31527 16204 33272 16232
rect 34659 16204 34704 16232
rect 31527 16201 31539 16204
rect 31481 16195 31539 16201
rect 12897 16167 12955 16173
rect 12897 16164 12909 16167
rect 6886 16136 12909 16164
rect 3145 16099 3203 16105
rect 3145 16065 3157 16099
rect 3191 16096 3203 16099
rect 6886 16096 6914 16136
rect 12897 16133 12909 16136
rect 12943 16133 12955 16167
rect 12897 16127 12955 16133
rect 21358 16124 21364 16176
rect 21416 16164 21422 16176
rect 25314 16173 25320 16176
rect 25308 16164 25320 16173
rect 21416 16136 25176 16164
rect 25275 16136 25320 16164
rect 21416 16124 21422 16136
rect 12710 16096 12716 16108
rect 3191 16068 6914 16096
rect 12671 16068 12716 16096
rect 3191 16065 3203 16068
rect 3145 16059 3203 16065
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21968 16068 22017 16096
rect 21968 16056 21974 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22186 16096 22192 16108
rect 22147 16068 22192 16096
rect 22005 16059 22063 16065
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 22281 16099 22339 16105
rect 22281 16065 22293 16099
rect 22327 16096 22339 16099
rect 22738 16096 22744 16108
rect 22327 16068 22744 16096
rect 22327 16065 22339 16068
rect 22281 16059 22339 16065
rect 22738 16056 22744 16068
rect 22796 16056 22802 16108
rect 24305 16099 24363 16105
rect 24305 16065 24317 16099
rect 24351 16096 24363 16099
rect 24762 16096 24768 16108
rect 24351 16068 24768 16096
rect 24351 16065 24363 16068
rect 24305 16059 24363 16065
rect 24762 16056 24768 16068
rect 24820 16056 24826 16108
rect 25038 16096 25044 16108
rect 24999 16068 25044 16096
rect 25038 16056 25044 16068
rect 25096 16056 25102 16108
rect 25148 16096 25176 16136
rect 25308 16127 25320 16136
rect 25314 16124 25320 16127
rect 25372 16124 25378 16176
rect 30466 16164 30472 16176
rect 26804 16136 30472 16164
rect 26804 16096 26832 16136
rect 30466 16124 30472 16136
rect 30524 16124 30530 16176
rect 30834 16124 30840 16176
rect 30892 16164 30898 16176
rect 31570 16164 31576 16176
rect 30892 16136 31576 16164
rect 30892 16124 30898 16136
rect 31570 16124 31576 16136
rect 31628 16124 31634 16176
rect 33134 16164 33140 16176
rect 31680 16136 33140 16164
rect 25148 16068 26832 16096
rect 26878 16056 26884 16108
rect 26936 16096 26942 16108
rect 27229 16099 27287 16105
rect 27229 16096 27241 16099
rect 26936 16068 27241 16096
rect 26936 16056 26942 16068
rect 27229 16065 27241 16068
rect 27275 16065 27287 16099
rect 27229 16059 27287 16065
rect 27706 16056 27712 16108
rect 27764 16096 27770 16108
rect 28997 16099 29055 16105
rect 28997 16096 29009 16099
rect 27764 16068 29009 16096
rect 27764 16056 27770 16068
rect 28997 16065 29009 16068
rect 29043 16065 29055 16099
rect 28997 16059 29055 16065
rect 30098 16056 30104 16108
rect 30156 16096 30162 16108
rect 31680 16105 31708 16136
rect 33134 16124 33140 16136
rect 33192 16124 33198 16176
rect 33244 16164 33272 16204
rect 34698 16192 34704 16204
rect 34756 16192 34762 16244
rect 35621 16235 35679 16241
rect 35621 16201 35633 16235
rect 35667 16201 35679 16235
rect 35621 16195 35679 16201
rect 36081 16235 36139 16241
rect 36081 16201 36093 16235
rect 36127 16232 36139 16235
rect 36538 16232 36544 16244
rect 36127 16204 36544 16232
rect 36127 16201 36139 16204
rect 36081 16195 36139 16201
rect 33566 16167 33624 16173
rect 33566 16164 33578 16167
rect 33244 16136 33578 16164
rect 33566 16133 33578 16136
rect 33612 16133 33624 16167
rect 33566 16127 33624 16133
rect 30285 16099 30343 16105
rect 30285 16096 30297 16099
rect 30156 16068 30297 16096
rect 30156 16056 30162 16068
rect 30285 16065 30297 16068
rect 30331 16065 30343 16099
rect 30285 16059 30343 16065
rect 31113 16099 31171 16105
rect 31113 16065 31125 16099
rect 31159 16065 31171 16099
rect 31113 16059 31171 16065
rect 31665 16099 31723 16105
rect 31665 16065 31677 16099
rect 31711 16065 31723 16099
rect 31665 16059 31723 16065
rect 12529 16031 12587 16037
rect 12529 15997 12541 16031
rect 12575 16028 12587 16031
rect 23290 16028 23296 16040
rect 12575 16000 23296 16028
rect 12575 15997 12587 16000
rect 12529 15991 12587 15997
rect 23290 15988 23296 16000
rect 23348 15988 23354 16040
rect 24578 16028 24584 16040
rect 24539 16000 24584 16028
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 26970 16028 26976 16040
rect 26931 16000 26976 16028
rect 26970 15988 26976 16000
rect 27028 15988 27034 16040
rect 28813 16031 28871 16037
rect 28813 15997 28825 16031
rect 28859 15997 28871 16031
rect 29178 16028 29184 16040
rect 29139 16000 29184 16028
rect 28813 15991 28871 15997
rect 28828 15960 28856 15991
rect 29178 15988 29184 16000
rect 29236 15988 29242 16040
rect 31128 16028 31156 16059
rect 32398 16056 32404 16108
rect 32456 16096 32462 16108
rect 32677 16099 32735 16105
rect 32677 16096 32689 16099
rect 32456 16068 32689 16096
rect 32456 16056 32462 16068
rect 32677 16065 32689 16068
rect 32723 16065 32735 16099
rect 32858 16096 32864 16108
rect 32819 16068 32864 16096
rect 32677 16059 32735 16065
rect 32858 16056 32864 16068
rect 32916 16056 32922 16108
rect 32953 16099 33011 16105
rect 32953 16065 32965 16099
rect 32999 16065 33011 16099
rect 32953 16059 33011 16065
rect 32122 16028 32128 16040
rect 31128 16000 32128 16028
rect 32122 15988 32128 16000
rect 32180 15988 32186 16040
rect 32214 15988 32220 16040
rect 32272 16028 32278 16040
rect 32968 16028 32996 16059
rect 33042 16056 33048 16108
rect 33100 16096 33106 16108
rect 33321 16099 33379 16105
rect 33321 16096 33333 16099
rect 33100 16068 33333 16096
rect 33100 16056 33106 16068
rect 33321 16065 33333 16068
rect 33367 16065 33379 16099
rect 35253 16099 35311 16105
rect 33321 16059 33379 16065
rect 33428 16068 34376 16096
rect 32272 16000 32996 16028
rect 32272 15988 32278 16000
rect 33134 15988 33140 16040
rect 33192 16028 33198 16040
rect 33428 16028 33456 16068
rect 33192 16000 33456 16028
rect 34348 16028 34376 16068
rect 35253 16065 35265 16099
rect 35299 16096 35311 16099
rect 35636 16096 35664 16195
rect 36538 16192 36544 16204
rect 36596 16192 36602 16244
rect 37826 16232 37832 16244
rect 37476 16204 37832 16232
rect 35299 16068 35664 16096
rect 35299 16065 35311 16068
rect 35253 16059 35311 16065
rect 35710 16056 35716 16108
rect 35768 16096 35774 16108
rect 37476 16105 37504 16204
rect 37826 16192 37832 16204
rect 37884 16192 37890 16244
rect 38654 16192 38660 16244
rect 38712 16232 38718 16244
rect 43070 16232 43076 16244
rect 38712 16204 43076 16232
rect 38712 16192 38718 16204
rect 43070 16192 43076 16204
rect 43128 16192 43134 16244
rect 43162 16192 43168 16244
rect 43220 16241 43226 16244
rect 43220 16232 43231 16241
rect 51350 16232 51356 16244
rect 43220 16204 43265 16232
rect 43456 16204 51356 16232
rect 43220 16195 43231 16204
rect 43220 16192 43226 16195
rect 42797 16167 42855 16173
rect 42797 16133 42809 16167
rect 42843 16164 42855 16167
rect 43346 16164 43352 16176
rect 42843 16136 43352 16164
rect 42843 16133 42855 16136
rect 42797 16127 42855 16133
rect 43346 16124 43352 16136
rect 43404 16124 43410 16176
rect 35989 16099 36047 16105
rect 35989 16096 36001 16099
rect 35768 16068 36001 16096
rect 35768 16056 35774 16068
rect 35989 16065 36001 16068
rect 36035 16065 36047 16099
rect 35989 16059 36047 16065
rect 37461 16099 37519 16105
rect 37461 16065 37473 16099
rect 37507 16065 37519 16099
rect 37461 16059 37519 16065
rect 37550 16056 37556 16108
rect 37608 16096 37614 16108
rect 37645 16099 37703 16105
rect 37645 16096 37657 16099
rect 37608 16068 37657 16096
rect 37608 16056 37614 16068
rect 37645 16065 37657 16068
rect 37691 16065 37703 16099
rect 37645 16059 37703 16065
rect 37734 16056 37740 16108
rect 37792 16096 37798 16108
rect 37792 16068 37837 16096
rect 37792 16056 37798 16068
rect 41414 16056 41420 16108
rect 41472 16096 41478 16108
rect 41509 16099 41567 16105
rect 41509 16096 41521 16099
rect 41472 16068 41521 16096
rect 41472 16056 41478 16068
rect 41509 16065 41521 16068
rect 41555 16065 41567 16099
rect 42610 16096 42616 16108
rect 42571 16068 42616 16096
rect 41509 16059 41567 16065
rect 42610 16056 42616 16068
rect 42668 16056 42674 16108
rect 42886 16096 42892 16108
rect 42847 16068 42892 16096
rect 42886 16056 42892 16068
rect 42944 16056 42950 16108
rect 42978 16056 42984 16108
rect 43036 16105 43042 16108
rect 43036 16096 43044 16105
rect 43036 16068 43081 16096
rect 43036 16059 43044 16068
rect 43036 16056 43042 16059
rect 36173 16031 36231 16037
rect 36173 16028 36185 16031
rect 34348 16000 36185 16028
rect 33192 15988 33198 16000
rect 36173 15997 36185 16000
rect 36219 15997 36231 16031
rect 36173 15991 36231 15997
rect 37826 15988 37832 16040
rect 37884 16028 37890 16040
rect 43456 16028 43484 16204
rect 51350 16192 51356 16204
rect 51408 16192 51414 16244
rect 51629 16235 51687 16241
rect 51629 16201 51641 16235
rect 51675 16232 51687 16235
rect 51994 16232 52000 16244
rect 51675 16204 52000 16232
rect 51675 16201 51687 16204
rect 51629 16195 51687 16201
rect 51994 16192 52000 16204
rect 52052 16192 52058 16244
rect 52454 16192 52460 16244
rect 52512 16232 52518 16244
rect 53098 16232 53104 16244
rect 52512 16204 53104 16232
rect 52512 16192 52518 16204
rect 53098 16192 53104 16204
rect 53156 16192 53162 16244
rect 53190 16192 53196 16244
rect 53248 16232 53254 16244
rect 60734 16232 60740 16244
rect 53248 16204 60740 16232
rect 53248 16192 53254 16204
rect 60734 16192 60740 16204
rect 60792 16192 60798 16244
rect 65797 16235 65855 16241
rect 65797 16201 65809 16235
rect 65843 16232 65855 16235
rect 65978 16232 65984 16244
rect 65843 16204 65984 16232
rect 65843 16201 65855 16204
rect 65797 16195 65855 16201
rect 65978 16192 65984 16204
rect 66036 16192 66042 16244
rect 66070 16192 66076 16244
rect 66128 16232 66134 16244
rect 69385 16235 69443 16241
rect 69385 16232 69397 16235
rect 66128 16204 69397 16232
rect 66128 16192 66134 16204
rect 69385 16201 69397 16204
rect 69431 16201 69443 16235
rect 69385 16195 69443 16201
rect 71225 16235 71283 16241
rect 71225 16201 71237 16235
rect 71271 16232 71283 16235
rect 71961 16235 72019 16241
rect 71961 16232 71973 16235
rect 71271 16204 71973 16232
rect 71271 16201 71283 16204
rect 71225 16195 71283 16201
rect 71961 16201 71973 16204
rect 72007 16232 72019 16235
rect 72418 16232 72424 16244
rect 72007 16204 72424 16232
rect 72007 16201 72019 16204
rect 71961 16195 72019 16201
rect 72418 16192 72424 16204
rect 72476 16192 72482 16244
rect 43809 16167 43867 16173
rect 43809 16133 43821 16167
rect 43855 16164 43867 16167
rect 44637 16167 44695 16173
rect 44637 16164 44649 16167
rect 43855 16136 44649 16164
rect 43855 16133 43867 16136
rect 43809 16127 43867 16133
rect 44637 16133 44649 16136
rect 44683 16133 44695 16167
rect 45922 16164 45928 16176
rect 44637 16127 44695 16133
rect 45112 16136 45928 16164
rect 43622 16096 43628 16108
rect 43583 16068 43628 16096
rect 43622 16056 43628 16068
rect 43680 16056 43686 16108
rect 43898 16096 43904 16108
rect 43859 16068 43904 16096
rect 43898 16056 43904 16068
rect 43956 16056 43962 16108
rect 43990 16056 43996 16108
rect 44048 16105 44054 16108
rect 44048 16096 44056 16105
rect 44048 16068 44093 16096
rect 44048 16059 44056 16068
rect 44048 16056 44054 16059
rect 44726 16056 44732 16108
rect 44784 16096 44790 16108
rect 44821 16099 44879 16105
rect 44821 16096 44833 16099
rect 44784 16068 44833 16096
rect 44784 16056 44790 16068
rect 44821 16065 44833 16068
rect 44867 16065 44879 16099
rect 45002 16096 45008 16108
rect 44963 16068 45008 16096
rect 44821 16059 44879 16065
rect 45002 16056 45008 16068
rect 45060 16056 45066 16108
rect 45112 16105 45140 16136
rect 45922 16124 45928 16136
rect 45980 16124 45986 16176
rect 46474 16164 46480 16176
rect 46435 16136 46480 16164
rect 46474 16124 46480 16136
rect 46532 16124 46538 16176
rect 46569 16167 46627 16173
rect 46569 16133 46581 16167
rect 46615 16164 46627 16167
rect 46842 16164 46848 16176
rect 46615 16136 46848 16164
rect 46615 16133 46627 16136
rect 46569 16127 46627 16133
rect 46842 16124 46848 16136
rect 46900 16124 46906 16176
rect 47394 16124 47400 16176
rect 47452 16164 47458 16176
rect 50798 16164 50804 16176
rect 47452 16136 47900 16164
rect 47452 16124 47458 16136
rect 45097 16099 45155 16105
rect 45097 16065 45109 16099
rect 45143 16065 45155 16099
rect 45097 16059 45155 16065
rect 45370 16056 45376 16108
rect 45428 16096 45434 16108
rect 45833 16099 45891 16105
rect 45833 16096 45845 16099
rect 45428 16068 45845 16096
rect 45428 16056 45434 16068
rect 45833 16065 45845 16068
rect 45879 16065 45891 16099
rect 45833 16059 45891 16065
rect 46198 16056 46204 16108
rect 46256 16096 46262 16108
rect 46293 16099 46351 16105
rect 46293 16096 46305 16099
rect 46256 16068 46305 16096
rect 46256 16056 46262 16068
rect 46293 16065 46305 16068
rect 46339 16065 46351 16099
rect 46293 16059 46351 16065
rect 46382 16056 46388 16108
rect 46440 16096 46446 16108
rect 46666 16099 46724 16105
rect 46666 16096 46678 16099
rect 46440 16068 46678 16096
rect 46440 16056 46446 16068
rect 46666 16065 46678 16068
rect 46712 16096 46724 16099
rect 46712 16068 46934 16096
rect 46712 16065 46724 16068
rect 46666 16059 46724 16065
rect 37884 16000 43484 16028
rect 46906 16028 46934 16068
rect 47118 16056 47124 16108
rect 47176 16096 47182 16108
rect 47581 16099 47639 16105
rect 47581 16096 47593 16099
rect 47176 16068 47593 16096
rect 47176 16056 47182 16068
rect 47581 16065 47593 16068
rect 47627 16065 47639 16099
rect 47762 16096 47768 16108
rect 47723 16068 47768 16096
rect 47581 16059 47639 16065
rect 47486 16028 47492 16040
rect 46906 16000 47492 16028
rect 37884 15988 37890 16000
rect 47486 15988 47492 16000
rect 47544 15988 47550 16040
rect 47596 16028 47624 16059
rect 47762 16056 47768 16068
rect 47820 16056 47826 16108
rect 47872 16105 47900 16136
rect 47964 16136 50804 16164
rect 47857 16099 47915 16105
rect 47857 16065 47869 16099
rect 47903 16065 47915 16099
rect 47857 16059 47915 16065
rect 47670 16028 47676 16040
rect 47596 16000 47676 16028
rect 47670 15988 47676 16000
rect 47728 15988 47734 16040
rect 47780 16028 47808 16056
rect 47964 16028 47992 16136
rect 50798 16124 50804 16136
rect 50856 16124 50862 16176
rect 50890 16124 50896 16176
rect 50948 16164 50954 16176
rect 51166 16164 51172 16176
rect 50948 16136 51172 16164
rect 50948 16124 50954 16136
rect 51166 16124 51172 16136
rect 51224 16124 51230 16176
rect 51261 16167 51319 16173
rect 51261 16133 51273 16167
rect 51307 16164 51319 16167
rect 52917 16167 52975 16173
rect 52917 16164 52929 16167
rect 51307 16136 52929 16164
rect 51307 16133 51319 16136
rect 51261 16127 51319 16133
rect 52917 16133 52929 16136
rect 52963 16133 52975 16167
rect 53742 16164 53748 16176
rect 52917 16127 52975 16133
rect 53024 16136 53748 16164
rect 48222 16056 48228 16108
rect 48280 16096 48286 16108
rect 48406 16096 48412 16108
rect 48280 16068 48325 16096
rect 48367 16068 48412 16096
rect 48280 16056 48286 16068
rect 48406 16056 48412 16068
rect 48464 16056 48470 16108
rect 48501 16099 48559 16105
rect 48501 16065 48513 16099
rect 48547 16065 48559 16099
rect 48501 16059 48559 16065
rect 47780 16000 47992 16028
rect 48038 15988 48044 16040
rect 48096 16028 48102 16040
rect 48516 16028 48544 16059
rect 48590 16056 48596 16108
rect 48648 16096 48654 16108
rect 49970 16096 49976 16108
rect 48648 16068 49976 16096
rect 48648 16056 48654 16068
rect 49970 16056 49976 16068
rect 50028 16056 50034 16108
rect 50065 16099 50123 16105
rect 50065 16065 50077 16099
rect 50111 16096 50123 16099
rect 50154 16096 50160 16108
rect 50111 16068 50160 16096
rect 50111 16065 50123 16068
rect 50065 16059 50123 16065
rect 50154 16056 50160 16068
rect 50212 16056 50218 16108
rect 50249 16099 50307 16105
rect 50249 16065 50261 16099
rect 50295 16065 50307 16099
rect 50249 16059 50307 16065
rect 49602 16028 49608 16040
rect 48096 16000 48268 16028
rect 48516 16000 49608 16028
rect 48096 15988 48102 16000
rect 29086 15960 29092 15972
rect 28828 15932 29092 15960
rect 29086 15920 29092 15932
rect 29144 15920 29150 15972
rect 30929 15963 30987 15969
rect 30929 15929 30941 15963
rect 30975 15960 30987 15963
rect 31938 15960 31944 15972
rect 30975 15932 31944 15960
rect 30975 15929 30987 15932
rect 30929 15923 30987 15929
rect 31938 15920 31944 15932
rect 31996 15920 32002 15972
rect 32858 15920 32864 15972
rect 32916 15960 32922 15972
rect 33318 15960 33324 15972
rect 32916 15932 33324 15960
rect 32916 15920 32922 15932
rect 33318 15920 33324 15932
rect 33376 15920 33382 15972
rect 35342 15920 35348 15972
rect 35400 15960 35406 15972
rect 40678 15960 40684 15972
rect 35400 15932 40684 15960
rect 35400 15920 35406 15932
rect 40678 15920 40684 15932
rect 40736 15960 40742 15972
rect 42978 15960 42984 15972
rect 40736 15932 42984 15960
rect 40736 15920 40742 15932
rect 42978 15920 42984 15932
rect 43036 15920 43042 15972
rect 44100 15932 47164 15960
rect 23937 15895 23995 15901
rect 23937 15861 23949 15895
rect 23983 15892 23995 15895
rect 25222 15892 25228 15904
rect 23983 15864 25228 15892
rect 23983 15861 23995 15864
rect 23937 15855 23995 15861
rect 25222 15852 25228 15864
rect 25280 15852 25286 15904
rect 26421 15895 26479 15901
rect 26421 15861 26433 15895
rect 26467 15892 26479 15895
rect 26970 15892 26976 15904
rect 26467 15864 26976 15892
rect 26467 15861 26479 15864
rect 26421 15855 26479 15861
rect 26970 15852 26976 15864
rect 27028 15852 27034 15904
rect 27706 15852 27712 15904
rect 27764 15892 27770 15904
rect 28353 15895 28411 15901
rect 28353 15892 28365 15895
rect 27764 15864 28365 15892
rect 27764 15852 27770 15864
rect 28353 15861 28365 15864
rect 28399 15861 28411 15895
rect 28353 15855 28411 15861
rect 32493 15895 32551 15901
rect 32493 15861 32505 15895
rect 32539 15892 32551 15895
rect 34238 15892 34244 15904
rect 32539 15864 34244 15892
rect 32539 15861 32551 15864
rect 32493 15855 32551 15861
rect 34238 15852 34244 15864
rect 34296 15852 34302 15904
rect 35069 15895 35127 15901
rect 35069 15861 35081 15895
rect 35115 15892 35127 15895
rect 36354 15892 36360 15904
rect 35115 15864 36360 15892
rect 35115 15861 35127 15864
rect 35069 15855 35127 15861
rect 36354 15852 36360 15864
rect 36412 15852 36418 15904
rect 37277 15895 37335 15901
rect 37277 15861 37289 15895
rect 37323 15892 37335 15895
rect 37458 15892 37464 15904
rect 37323 15864 37464 15892
rect 37323 15861 37335 15864
rect 37277 15855 37335 15861
rect 37458 15852 37464 15864
rect 37516 15852 37522 15904
rect 41601 15895 41659 15901
rect 41601 15861 41613 15895
rect 41647 15892 41659 15895
rect 44100 15892 44128 15932
rect 41647 15864 44128 15892
rect 44177 15895 44235 15901
rect 41647 15861 41659 15864
rect 41601 15855 41659 15861
rect 44177 15861 44189 15895
rect 44223 15892 44235 15895
rect 44450 15892 44456 15904
rect 44223 15864 44456 15892
rect 44223 15861 44235 15864
rect 44177 15855 44235 15861
rect 44450 15852 44456 15864
rect 44508 15852 44514 15904
rect 45646 15892 45652 15904
rect 45607 15864 45652 15892
rect 45646 15852 45652 15864
rect 45704 15852 45710 15904
rect 46658 15852 46664 15904
rect 46716 15892 46722 15904
rect 46845 15895 46903 15901
rect 46845 15892 46857 15895
rect 46716 15864 46857 15892
rect 46716 15852 46722 15864
rect 46845 15861 46857 15864
rect 46891 15861 46903 15895
rect 47136 15892 47164 15932
rect 47210 15920 47216 15972
rect 47268 15960 47274 15972
rect 47581 15963 47639 15969
rect 47581 15960 47593 15963
rect 47268 15932 47593 15960
rect 47268 15920 47274 15932
rect 47581 15929 47593 15932
rect 47627 15929 47639 15963
rect 48130 15960 48136 15972
rect 47581 15923 47639 15929
rect 47688 15932 48136 15960
rect 47688 15892 47716 15932
rect 48130 15920 48136 15932
rect 48188 15920 48194 15972
rect 48240 15969 48268 16000
rect 49602 15988 49608 16000
rect 49660 15988 49666 16040
rect 49694 15988 49700 16040
rect 49752 16028 49758 16040
rect 49878 16028 49884 16040
rect 49752 16000 49884 16028
rect 49752 15988 49758 16000
rect 49878 15988 49884 16000
rect 49936 16028 49942 16040
rect 50264 16028 50292 16059
rect 50338 16056 50344 16108
rect 50396 16096 50402 16108
rect 50396 16068 50441 16096
rect 50396 16056 50402 16068
rect 50614 16056 50620 16108
rect 50672 16096 50678 16108
rect 51445 16099 51503 16105
rect 51445 16096 51457 16099
rect 50672 16068 51457 16096
rect 50672 16056 50678 16068
rect 51445 16065 51457 16068
rect 51491 16096 51503 16099
rect 51534 16096 51540 16108
rect 51491 16068 51540 16096
rect 51491 16065 51503 16068
rect 51445 16059 51503 16065
rect 51534 16056 51540 16068
rect 51592 16056 51598 16108
rect 51721 16099 51779 16105
rect 51721 16065 51733 16099
rect 51767 16096 51779 16099
rect 51902 16096 51908 16108
rect 51767 16068 51908 16096
rect 51767 16065 51779 16068
rect 51721 16059 51779 16065
rect 51902 16056 51908 16068
rect 51960 16096 51966 16108
rect 52454 16096 52460 16108
rect 51960 16068 52460 16096
rect 51960 16056 51966 16068
rect 52454 16056 52460 16068
rect 52512 16056 52518 16108
rect 52733 16099 52791 16105
rect 52733 16065 52745 16099
rect 52779 16065 52791 16099
rect 52733 16059 52791 16065
rect 49936 16000 50292 16028
rect 49936 15988 49942 16000
rect 50522 15988 50528 16040
rect 50580 16028 50586 16040
rect 52638 16028 52644 16040
rect 50580 16000 52644 16028
rect 50580 15988 50586 16000
rect 52638 15988 52644 16000
rect 52696 15988 52702 16040
rect 52748 16028 52776 16059
rect 52822 16056 52828 16108
rect 52880 16096 52886 16108
rect 53024 16105 53052 16136
rect 53742 16124 53748 16136
rect 53800 16124 53806 16176
rect 54938 16124 54944 16176
rect 54996 16164 55002 16176
rect 57149 16167 57207 16173
rect 57149 16164 57161 16167
rect 54996 16136 57161 16164
rect 54996 16124 55002 16136
rect 57149 16133 57161 16136
rect 57195 16164 57207 16167
rect 58434 16164 58440 16176
rect 57195 16136 58440 16164
rect 57195 16133 57207 16136
rect 57149 16127 57207 16133
rect 58434 16124 58440 16136
rect 58492 16124 58498 16176
rect 58618 16124 58624 16176
rect 58676 16164 58682 16176
rect 58897 16167 58955 16173
rect 58676 16136 58848 16164
rect 58676 16124 58682 16136
rect 53190 16105 53196 16108
rect 53009 16099 53067 16105
rect 53009 16096 53021 16099
rect 52880 16068 53021 16096
rect 52880 16056 52886 16068
rect 53009 16065 53021 16068
rect 53055 16065 53067 16099
rect 53009 16059 53067 16065
rect 53153 16099 53196 16105
rect 53153 16065 53165 16099
rect 53153 16059 53196 16065
rect 53190 16056 53196 16059
rect 53248 16056 53254 16108
rect 53837 16099 53895 16105
rect 53837 16065 53849 16099
rect 53883 16065 53895 16099
rect 53837 16059 53895 16065
rect 53852 16028 53880 16059
rect 53926 16056 53932 16108
rect 53984 16096 53990 16108
rect 54113 16099 54171 16105
rect 54113 16096 54125 16099
rect 53984 16068 54125 16096
rect 53984 16056 53990 16068
rect 54113 16065 54125 16068
rect 54159 16065 54171 16099
rect 54113 16059 54171 16065
rect 54570 16056 54576 16108
rect 54628 16096 54634 16108
rect 55125 16099 55183 16105
rect 55125 16096 55137 16099
rect 54628 16068 55137 16096
rect 54628 16056 54634 16068
rect 55125 16065 55137 16068
rect 55171 16096 55183 16099
rect 55214 16096 55220 16108
rect 55171 16068 55220 16096
rect 55171 16065 55183 16068
rect 55125 16059 55183 16065
rect 55214 16056 55220 16068
rect 55272 16056 55278 16108
rect 55392 16099 55450 16105
rect 55392 16065 55404 16099
rect 55438 16096 55450 16099
rect 56778 16096 56784 16108
rect 55438 16068 56784 16096
rect 55438 16065 55450 16068
rect 55392 16059 55450 16065
rect 56778 16056 56784 16068
rect 56836 16056 56842 16108
rect 56965 16099 57023 16105
rect 56965 16065 56977 16099
rect 57011 16065 57023 16099
rect 56965 16059 57023 16065
rect 54202 16028 54208 16040
rect 52748 16000 53788 16028
rect 53852 16000 54208 16028
rect 48225 15963 48283 15969
rect 48225 15929 48237 15963
rect 48271 15929 48283 15963
rect 50154 15960 50160 15972
rect 48225 15923 48283 15929
rect 48424 15932 50160 15960
rect 47136 15864 47716 15892
rect 46845 15855 46903 15861
rect 47762 15852 47768 15904
rect 47820 15892 47826 15904
rect 48424 15892 48452 15932
rect 50154 15920 50160 15932
rect 50212 15920 50218 15972
rect 53285 15963 53343 15969
rect 53285 15960 53297 15963
rect 51184 15932 53297 15960
rect 49878 15892 49884 15904
rect 47820 15864 48452 15892
rect 49839 15864 49884 15892
rect 47820 15852 47826 15864
rect 49878 15852 49884 15864
rect 49936 15852 49942 15904
rect 50706 15852 50712 15904
rect 50764 15892 50770 15904
rect 51184 15892 51212 15932
rect 53285 15929 53297 15932
rect 53331 15929 53343 15963
rect 53760 15960 53788 16000
rect 54202 15988 54208 16000
rect 54260 15988 54266 16040
rect 56318 15988 56324 16040
rect 56376 16028 56382 16040
rect 56980 16028 57008 16059
rect 57882 16056 57888 16108
rect 57940 16096 57946 16108
rect 58069 16099 58127 16105
rect 58069 16096 58081 16099
rect 57940 16068 58081 16096
rect 57940 16056 57946 16068
rect 58069 16065 58081 16068
rect 58115 16065 58127 16099
rect 58250 16096 58256 16108
rect 58211 16068 58256 16096
rect 58069 16059 58127 16065
rect 58250 16056 58256 16068
rect 58308 16056 58314 16108
rect 58342 16056 58348 16108
rect 58400 16096 58406 16108
rect 58400 16068 58445 16096
rect 58400 16056 58406 16068
rect 58526 16056 58532 16108
rect 58584 16096 58590 16108
rect 58713 16099 58771 16105
rect 58713 16096 58725 16099
rect 58584 16068 58725 16096
rect 58584 16056 58590 16068
rect 58713 16065 58725 16068
rect 58759 16065 58771 16099
rect 58820 16096 58848 16136
rect 58897 16133 58909 16167
rect 58943 16164 58955 16167
rect 59725 16167 59783 16173
rect 59725 16164 59737 16167
rect 58943 16136 59737 16164
rect 58943 16133 58955 16136
rect 58897 16127 58955 16133
rect 59725 16133 59737 16136
rect 59771 16133 59783 16167
rect 64693 16167 64751 16173
rect 59725 16127 59783 16133
rect 59832 16136 64552 16164
rect 58986 16096 58992 16108
rect 58820 16068 58992 16096
rect 58713 16059 58771 16065
rect 58986 16056 58992 16068
rect 59044 16056 59050 16108
rect 59170 16105 59176 16108
rect 59133 16099 59176 16105
rect 59133 16065 59145 16099
rect 59133 16059 59176 16065
rect 59170 16056 59176 16059
rect 59228 16056 59234 16108
rect 59832 16096 59860 16136
rect 59372 16068 59860 16096
rect 59909 16099 59967 16105
rect 57974 16028 57980 16040
rect 56376 16000 57980 16028
rect 56376 15988 56382 16000
rect 57974 15988 57980 16000
rect 58032 15988 58038 16040
rect 59372 16028 59400 16068
rect 59909 16065 59921 16099
rect 59955 16065 59967 16099
rect 59909 16059 59967 16065
rect 58084 16000 59400 16028
rect 59924 16028 59952 16059
rect 59998 16056 60004 16108
rect 60056 16096 60062 16108
rect 60093 16099 60151 16105
rect 60093 16096 60105 16099
rect 60056 16068 60105 16096
rect 60056 16056 60062 16068
rect 60093 16065 60105 16068
rect 60139 16065 60151 16099
rect 60093 16059 60151 16065
rect 60185 16099 60243 16105
rect 60185 16065 60197 16099
rect 60231 16096 60243 16099
rect 60458 16096 60464 16108
rect 60231 16068 60464 16096
rect 60231 16065 60243 16068
rect 60185 16059 60243 16065
rect 60458 16056 60464 16068
rect 60516 16056 60522 16108
rect 60829 16099 60887 16105
rect 60829 16096 60841 16099
rect 60706 16068 60841 16096
rect 60274 16028 60280 16040
rect 59924 16000 60280 16028
rect 55030 15960 55036 15972
rect 53760 15932 55036 15960
rect 53285 15923 53343 15929
rect 55030 15920 55036 15932
rect 55088 15920 55094 15972
rect 58084 15969 58112 16000
rect 60274 15988 60280 16000
rect 60332 15988 60338 16040
rect 60366 15988 60372 16040
rect 60424 16028 60430 16040
rect 60706 16028 60734 16068
rect 60829 16065 60841 16068
rect 60875 16096 60887 16099
rect 62114 16096 62120 16108
rect 60875 16068 62120 16096
rect 60875 16065 60887 16068
rect 60829 16059 60887 16065
rect 62114 16056 62120 16068
rect 62172 16056 62178 16108
rect 62301 16099 62359 16105
rect 62301 16065 62313 16099
rect 62347 16096 62359 16099
rect 62390 16096 62396 16108
rect 62347 16068 62396 16096
rect 62347 16065 62359 16068
rect 62301 16059 62359 16065
rect 62390 16056 62396 16068
rect 62448 16056 62454 16108
rect 62758 16056 62764 16108
rect 62816 16096 62822 16108
rect 62816 16068 62988 16096
rect 62816 16056 62822 16068
rect 60424 16000 60734 16028
rect 61105 16031 61163 16037
rect 60424 15988 60430 16000
rect 61105 15997 61117 16031
rect 61151 16028 61163 16031
rect 62206 16028 62212 16040
rect 61151 16000 62212 16028
rect 61151 15997 61163 16000
rect 61105 15991 61163 15997
rect 62206 15988 62212 16000
rect 62264 15988 62270 16040
rect 62960 16028 62988 16068
rect 63034 16056 63040 16108
rect 63092 16096 63098 16108
rect 63092 16068 63137 16096
rect 63092 16056 63098 16068
rect 63218 16056 63224 16108
rect 63276 16096 63282 16108
rect 64524 16105 64552 16136
rect 64693 16133 64705 16167
rect 64739 16164 64751 16167
rect 65429 16167 65487 16173
rect 65429 16164 65441 16167
rect 64739 16136 65441 16164
rect 64739 16133 64751 16136
rect 64693 16127 64751 16133
rect 65429 16133 65441 16136
rect 65475 16133 65487 16167
rect 69750 16164 69756 16176
rect 65429 16127 65487 16133
rect 68480 16136 69756 16164
rect 63405 16099 63463 16105
rect 63276 16068 63321 16096
rect 63276 16056 63282 16068
rect 63405 16065 63417 16099
rect 63451 16096 63463 16099
rect 63957 16099 64015 16105
rect 63957 16096 63969 16099
rect 63451 16068 63969 16096
rect 63451 16065 63463 16068
rect 63405 16059 63463 16065
rect 63957 16065 63969 16068
rect 64003 16065 64015 16099
rect 63957 16059 64015 16065
rect 64509 16099 64567 16105
rect 64509 16065 64521 16099
rect 64555 16065 64567 16099
rect 64509 16059 64567 16065
rect 64598 16056 64604 16108
rect 64656 16096 64662 16108
rect 64785 16099 64843 16105
rect 64785 16096 64797 16099
rect 64656 16068 64797 16096
rect 64656 16056 64662 16068
rect 64785 16065 64797 16068
rect 64831 16065 64843 16099
rect 64785 16059 64843 16065
rect 64874 16056 64880 16108
rect 64932 16096 64938 16108
rect 65613 16099 65671 16105
rect 64932 16068 64977 16096
rect 64932 16056 64938 16068
rect 65613 16065 65625 16099
rect 65659 16096 65671 16099
rect 65702 16096 65708 16108
rect 65659 16068 65708 16096
rect 65659 16065 65671 16068
rect 65613 16059 65671 16065
rect 65702 16056 65708 16068
rect 65760 16056 65766 16108
rect 68480 16105 68508 16136
rect 69750 16124 69756 16136
rect 69808 16124 69814 16176
rect 73062 16124 73068 16176
rect 73120 16164 73126 16176
rect 73120 16136 73844 16164
rect 73120 16124 73126 16136
rect 65889 16099 65947 16105
rect 65889 16065 65901 16099
rect 65935 16065 65947 16099
rect 65889 16059 65947 16065
rect 68465 16099 68523 16105
rect 68465 16065 68477 16099
rect 68511 16065 68523 16099
rect 69201 16099 69259 16105
rect 69201 16096 69213 16099
rect 68465 16059 68523 16065
rect 68572 16068 69213 16096
rect 65904 16028 65932 16059
rect 66438 16028 66444 16040
rect 62960 16000 66444 16028
rect 66438 15988 66444 16000
rect 66496 15988 66502 16040
rect 68094 15988 68100 16040
rect 68152 16028 68158 16040
rect 68572 16028 68600 16068
rect 69201 16065 69213 16068
rect 69247 16065 69259 16099
rect 69201 16059 69259 16065
rect 69477 16099 69535 16105
rect 69477 16065 69489 16099
rect 69523 16096 69535 16099
rect 69934 16096 69940 16108
rect 69523 16068 69940 16096
rect 69523 16065 69535 16068
rect 69477 16059 69535 16065
rect 69934 16056 69940 16068
rect 69992 16056 69998 16108
rect 70112 16099 70170 16105
rect 70112 16065 70124 16099
rect 70158 16096 70170 16099
rect 71866 16096 71872 16108
rect 70158 16068 71872 16096
rect 70158 16065 70170 16068
rect 70112 16059 70170 16065
rect 71866 16056 71872 16068
rect 71924 16056 71930 16108
rect 73816 16105 73844 16136
rect 72053 16099 72111 16105
rect 72053 16065 72065 16099
rect 72099 16096 72111 16099
rect 73801 16099 73859 16105
rect 72099 16068 73752 16096
rect 72099 16065 72111 16068
rect 72053 16059 72111 16065
rect 68152 16000 68600 16028
rect 68152 15988 68158 16000
rect 68922 15988 68928 16040
rect 68980 16028 68986 16040
rect 69845 16031 69903 16037
rect 69845 16028 69857 16031
rect 68980 16000 69857 16028
rect 68980 15988 68986 16000
rect 69845 15997 69857 16000
rect 69891 15997 69903 16031
rect 69845 15991 69903 15997
rect 71498 15988 71504 16040
rect 71556 16028 71562 16040
rect 72145 16031 72203 16037
rect 72145 16028 72157 16031
rect 71556 16000 72157 16028
rect 71556 15988 71562 16000
rect 72145 15997 72157 16000
rect 72191 15997 72203 16031
rect 73724 16028 73752 16068
rect 73801 16065 73813 16099
rect 73847 16065 73859 16099
rect 73801 16059 73859 16065
rect 88245 16099 88303 16105
rect 88245 16065 88257 16099
rect 88291 16065 88303 16099
rect 88245 16059 88303 16065
rect 86586 16028 86592 16040
rect 73724 16000 86592 16028
rect 72145 15991 72203 15997
rect 86586 15988 86592 16000
rect 86644 15988 86650 16040
rect 58069 15963 58127 15969
rect 58069 15929 58081 15963
rect 58115 15929 58127 15963
rect 58069 15923 58127 15929
rect 58158 15920 58164 15972
rect 58216 15960 58222 15972
rect 68557 15963 68615 15969
rect 68557 15960 68569 15963
rect 58216 15932 68569 15960
rect 58216 15920 58222 15932
rect 68557 15929 68569 15932
rect 68603 15929 68615 15963
rect 69474 15960 69480 15972
rect 68557 15923 68615 15929
rect 68664 15932 69480 15960
rect 50764 15864 51212 15892
rect 50764 15852 50770 15864
rect 53834 15852 53840 15904
rect 53892 15892 53898 15904
rect 56505 15895 56563 15901
rect 56505 15892 56517 15895
rect 53892 15864 56517 15892
rect 53892 15852 53898 15864
rect 56505 15861 56517 15864
rect 56551 15861 56563 15895
rect 56505 15855 56563 15861
rect 56594 15852 56600 15904
rect 56652 15892 56658 15904
rect 58710 15892 58716 15904
rect 56652 15864 58716 15892
rect 56652 15852 56658 15864
rect 58710 15852 58716 15864
rect 58768 15852 58774 15904
rect 58986 15852 58992 15904
rect 59044 15892 59050 15904
rect 59265 15895 59323 15901
rect 59265 15892 59277 15895
rect 59044 15864 59277 15892
rect 59044 15852 59050 15864
rect 59265 15861 59277 15864
rect 59311 15861 59323 15895
rect 63770 15892 63776 15904
rect 63731 15864 63776 15892
rect 59265 15855 59323 15861
rect 63770 15852 63776 15864
rect 63828 15852 63834 15904
rect 64966 15852 64972 15904
rect 65024 15892 65030 15904
rect 65061 15895 65119 15901
rect 65061 15892 65073 15895
rect 65024 15864 65073 15892
rect 65024 15852 65030 15864
rect 65061 15861 65073 15864
rect 65107 15861 65119 15895
rect 65061 15855 65119 15861
rect 65610 15852 65616 15904
rect 65668 15892 65674 15904
rect 68664 15892 68692 15932
rect 69474 15920 69480 15932
rect 69532 15920 69538 15972
rect 73617 15963 73675 15969
rect 73617 15929 73629 15963
rect 73663 15960 73675 15963
rect 88260 15960 88288 16059
rect 73663 15932 88288 15960
rect 73663 15929 73675 15932
rect 73617 15923 73675 15929
rect 65668 15864 68692 15892
rect 65668 15852 65674 15864
rect 68738 15852 68744 15904
rect 68796 15892 68802 15904
rect 69201 15895 69259 15901
rect 69201 15892 69213 15895
rect 68796 15864 69213 15892
rect 68796 15852 68802 15864
rect 69201 15861 69213 15864
rect 69247 15861 69259 15895
rect 69201 15855 69259 15861
rect 71593 15895 71651 15901
rect 71593 15861 71605 15895
rect 71639 15892 71651 15895
rect 72050 15892 72056 15904
rect 71639 15864 72056 15892
rect 71639 15861 71651 15864
rect 71593 15855 71651 15861
rect 72050 15852 72056 15864
rect 72108 15852 72114 15904
rect 88058 15892 88064 15904
rect 88019 15864 88064 15892
rect 88058 15852 88064 15864
rect 88116 15852 88122 15904
rect 1104 15802 88872 15824
rect 1104 15750 11924 15802
rect 11976 15750 11988 15802
rect 12040 15750 12052 15802
rect 12104 15750 12116 15802
rect 12168 15750 12180 15802
rect 12232 15750 33872 15802
rect 33924 15750 33936 15802
rect 33988 15750 34000 15802
rect 34052 15750 34064 15802
rect 34116 15750 34128 15802
rect 34180 15750 55820 15802
rect 55872 15750 55884 15802
rect 55936 15750 55948 15802
rect 56000 15750 56012 15802
rect 56064 15750 56076 15802
rect 56128 15750 77768 15802
rect 77820 15750 77832 15802
rect 77884 15750 77896 15802
rect 77948 15750 77960 15802
rect 78012 15750 78024 15802
rect 78076 15750 88872 15802
rect 1104 15728 88872 15750
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 25590 15688 25596 15700
rect 22244 15660 25596 15688
rect 22244 15648 22250 15660
rect 25590 15648 25596 15660
rect 25648 15648 25654 15700
rect 25958 15648 25964 15700
rect 26016 15688 26022 15700
rect 27433 15691 27491 15697
rect 27433 15688 27445 15691
rect 26016 15660 27445 15688
rect 26016 15648 26022 15660
rect 27433 15657 27445 15660
rect 27479 15657 27491 15691
rect 27433 15651 27491 15657
rect 27798 15648 27804 15700
rect 27856 15688 27862 15700
rect 32214 15688 32220 15700
rect 27856 15660 32220 15688
rect 27856 15648 27862 15660
rect 32214 15648 32220 15660
rect 32272 15648 32278 15700
rect 32401 15691 32459 15697
rect 32401 15657 32413 15691
rect 32447 15688 32459 15691
rect 32490 15688 32496 15700
rect 32447 15660 32496 15688
rect 32447 15657 32459 15660
rect 32401 15651 32459 15657
rect 32490 15648 32496 15660
rect 32548 15648 32554 15700
rect 33042 15688 33048 15700
rect 32784 15660 33048 15688
rect 27614 15580 27620 15632
rect 27672 15620 27678 15632
rect 30558 15620 30564 15632
rect 27672 15592 30564 15620
rect 27672 15580 27678 15592
rect 20898 15552 20904 15564
rect 20548 15524 20904 15552
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 20548 15493 20576 15524
rect 20898 15512 20904 15524
rect 20956 15552 20962 15564
rect 21910 15552 21916 15564
rect 20956 15524 21916 15552
rect 20956 15512 20962 15524
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 25406 15552 25412 15564
rect 23124 15524 25412 15552
rect 20533 15487 20591 15493
rect 20533 15453 20545 15487
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15484 20867 15487
rect 21082 15484 21088 15496
rect 20855 15456 21088 15484
rect 20855 15453 20867 15456
rect 20809 15447 20867 15453
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 22646 15444 22652 15496
rect 22704 15484 22710 15496
rect 23124 15493 23152 15524
rect 25406 15512 25412 15524
rect 25464 15512 25470 15564
rect 27890 15552 27896 15564
rect 27851 15524 27896 15552
rect 27890 15512 27896 15524
rect 27948 15512 27954 15564
rect 28092 15561 28120 15592
rect 30558 15580 30564 15592
rect 30616 15580 30622 15632
rect 28077 15555 28135 15561
rect 28077 15521 28089 15555
rect 28123 15521 28135 15555
rect 28077 15515 28135 15521
rect 28994 15512 29000 15564
rect 29052 15552 29058 15564
rect 32784 15561 32812 15660
rect 33042 15648 33048 15660
rect 33100 15648 33106 15700
rect 34422 15648 34428 15700
rect 34480 15688 34486 15700
rect 43990 15688 43996 15700
rect 34480 15660 37136 15688
rect 34480 15648 34486 15660
rect 35434 15580 35440 15632
rect 35492 15620 35498 15632
rect 37108 15620 37136 15660
rect 37568 15660 43996 15688
rect 37568 15620 37596 15660
rect 43990 15648 43996 15660
rect 44048 15648 44054 15700
rect 44085 15691 44143 15697
rect 44085 15657 44097 15691
rect 44131 15688 44143 15691
rect 45002 15688 45008 15700
rect 44131 15660 45008 15688
rect 44131 15657 44143 15660
rect 44085 15651 44143 15657
rect 45002 15648 45008 15660
rect 45060 15648 45066 15700
rect 45370 15688 45376 15700
rect 45331 15660 45376 15688
rect 45370 15648 45376 15660
rect 45428 15648 45434 15700
rect 46658 15688 46664 15700
rect 45756 15660 46664 15688
rect 45756 15620 45784 15660
rect 46658 15648 46664 15660
rect 46716 15648 46722 15700
rect 46750 15648 46756 15700
rect 46808 15688 46814 15700
rect 47489 15691 47547 15697
rect 47489 15688 47501 15691
rect 46808 15660 47501 15688
rect 46808 15648 46814 15660
rect 47489 15657 47501 15660
rect 47535 15657 47547 15691
rect 47489 15651 47547 15657
rect 48222 15648 48228 15700
rect 48280 15688 48286 15700
rect 50157 15691 50215 15697
rect 50157 15688 50169 15691
rect 48280 15660 50169 15688
rect 48280 15648 48286 15660
rect 50157 15657 50169 15660
rect 50203 15657 50215 15691
rect 50157 15651 50215 15657
rect 50246 15648 50252 15700
rect 50304 15688 50310 15700
rect 51442 15688 51448 15700
rect 50304 15660 51448 15688
rect 50304 15648 50310 15660
rect 51442 15648 51448 15660
rect 51500 15648 51506 15700
rect 51629 15691 51687 15697
rect 51629 15657 51641 15691
rect 51675 15688 51687 15691
rect 52362 15688 52368 15700
rect 51675 15660 52368 15688
rect 51675 15657 51687 15660
rect 51629 15651 51687 15657
rect 52362 15648 52368 15660
rect 52420 15648 52426 15700
rect 53374 15648 53380 15700
rect 53432 15688 53438 15700
rect 55309 15691 55367 15697
rect 55309 15688 55321 15691
rect 53432 15660 55321 15688
rect 53432 15648 53438 15660
rect 55309 15657 55321 15660
rect 55355 15657 55367 15691
rect 55309 15651 55367 15657
rect 57238 15648 57244 15700
rect 57296 15688 57302 15700
rect 58250 15688 58256 15700
rect 57296 15660 58256 15688
rect 57296 15648 57302 15660
rect 58250 15648 58256 15660
rect 58308 15648 58314 15700
rect 58986 15688 58992 15700
rect 58452 15660 58992 15688
rect 35492 15592 36124 15620
rect 37108 15592 37596 15620
rect 37712 15592 42564 15620
rect 35492 15580 35498 15592
rect 30377 15555 30435 15561
rect 30377 15552 30389 15555
rect 29052 15524 30389 15552
rect 29052 15512 29058 15524
rect 30377 15521 30389 15524
rect 30423 15521 30435 15555
rect 32769 15555 32827 15561
rect 32769 15552 32781 15555
rect 30377 15515 30435 15521
rect 32048 15524 32781 15552
rect 32048 15496 32076 15524
rect 32769 15521 32781 15524
rect 32815 15521 32827 15555
rect 35894 15552 35900 15564
rect 32769 15515 32827 15521
rect 35268 15524 35900 15552
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 22704 15456 23121 15484
rect 22704 15444 22710 15456
rect 23109 15453 23121 15456
rect 23155 15453 23167 15487
rect 25222 15484 25228 15496
rect 25183 15456 25228 15484
rect 23109 15447 23167 15453
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 25593 15487 25651 15493
rect 25593 15453 25605 15487
rect 25639 15484 25651 15487
rect 26142 15484 26148 15496
rect 25639 15456 26148 15484
rect 25639 15453 25651 15456
rect 25593 15447 25651 15453
rect 26142 15444 26148 15456
rect 26200 15444 26206 15496
rect 26970 15444 26976 15496
rect 27028 15484 27034 15496
rect 27801 15487 27859 15493
rect 27801 15484 27813 15487
rect 27028 15456 27813 15484
rect 27028 15444 27034 15456
rect 27801 15453 27813 15456
rect 27847 15453 27859 15487
rect 27801 15447 27859 15453
rect 28258 15444 28264 15496
rect 28316 15484 28322 15496
rect 29546 15484 29552 15496
rect 28316 15456 29552 15484
rect 28316 15444 28322 15456
rect 29546 15444 29552 15456
rect 29604 15484 29610 15496
rect 31021 15487 31079 15493
rect 31021 15484 31033 15487
rect 29604 15456 31033 15484
rect 29604 15444 29610 15456
rect 31021 15453 31033 15456
rect 31067 15484 31079 15487
rect 31110 15484 31116 15496
rect 31067 15456 31116 15484
rect 31067 15453 31079 15456
rect 31021 15447 31079 15453
rect 31110 15444 31116 15456
rect 31168 15484 31174 15496
rect 32030 15484 32036 15496
rect 31168 15456 32036 15484
rect 31168 15444 31174 15456
rect 32030 15444 32036 15456
rect 32088 15444 32094 15496
rect 32490 15444 32496 15496
rect 32548 15484 32554 15496
rect 33025 15487 33083 15493
rect 33025 15484 33037 15487
rect 32548 15456 33037 15484
rect 32548 15444 32554 15456
rect 33025 15453 33037 15456
rect 33071 15453 33083 15487
rect 35066 15484 35072 15496
rect 35027 15456 35072 15484
rect 33025 15447 33083 15453
rect 35066 15444 35072 15456
rect 35124 15444 35130 15496
rect 35268 15493 35296 15524
rect 35894 15512 35900 15524
rect 35952 15512 35958 15564
rect 36096 15561 36124 15592
rect 36081 15555 36139 15561
rect 36081 15521 36093 15555
rect 36127 15521 36139 15555
rect 36081 15515 36139 15521
rect 35253 15487 35311 15493
rect 35253 15453 35265 15487
rect 35299 15453 35311 15487
rect 35253 15447 35311 15453
rect 35342 15444 35348 15496
rect 35400 15484 35406 15496
rect 36096 15484 36124 15515
rect 37366 15512 37372 15564
rect 37424 15552 37430 15564
rect 37712 15552 37740 15592
rect 38378 15552 38384 15564
rect 37424 15524 37740 15552
rect 38339 15524 38384 15552
rect 37424 15512 37430 15524
rect 38378 15512 38384 15524
rect 38436 15512 38442 15564
rect 38565 15555 38623 15561
rect 38565 15521 38577 15555
rect 38611 15552 38623 15555
rect 41509 15555 41567 15561
rect 41509 15552 41521 15555
rect 38611 15524 41521 15552
rect 38611 15521 38623 15524
rect 38565 15515 38623 15521
rect 41509 15521 41521 15524
rect 41555 15521 41567 15555
rect 41509 15515 41567 15521
rect 37274 15484 37280 15496
rect 35400 15456 35445 15484
rect 36096 15456 37280 15484
rect 35400 15444 35406 15456
rect 37274 15444 37280 15456
rect 37332 15444 37338 15496
rect 37642 15444 37648 15496
rect 37700 15484 37706 15496
rect 38580 15484 38608 15515
rect 42334 15484 42340 15496
rect 37700 15456 38608 15484
rect 42295 15456 42340 15484
rect 37700 15444 37706 15456
rect 42334 15444 42340 15456
rect 42392 15444 42398 15496
rect 20714 15416 20720 15428
rect 20627 15388 20720 15416
rect 20714 15376 20720 15388
rect 20772 15416 20778 15428
rect 22186 15416 22192 15428
rect 20772 15388 22192 15416
rect 20772 15376 20778 15388
rect 22186 15376 22192 15388
rect 22244 15376 22250 15428
rect 23934 15376 23940 15428
rect 23992 15416 23998 15428
rect 23992 15388 25268 15416
rect 23992 15376 23998 15388
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 12342 15308 12348 15360
rect 12400 15348 12406 15360
rect 20349 15351 20407 15357
rect 20349 15348 20361 15351
rect 12400 15320 20361 15348
rect 12400 15308 12406 15320
rect 20349 15317 20361 15320
rect 20395 15317 20407 15351
rect 20349 15311 20407 15317
rect 22554 15308 22560 15360
rect 22612 15348 22618 15360
rect 23201 15351 23259 15357
rect 23201 15348 23213 15351
rect 22612 15320 23213 15348
rect 22612 15308 22618 15320
rect 23201 15317 23213 15320
rect 23247 15317 23259 15351
rect 23201 15311 23259 15317
rect 25041 15351 25099 15357
rect 25041 15317 25053 15351
rect 25087 15348 25099 15351
rect 25130 15348 25136 15360
rect 25087 15320 25136 15348
rect 25087 15317 25099 15320
rect 25041 15311 25099 15317
rect 25130 15308 25136 15320
rect 25188 15308 25194 15360
rect 25240 15348 25268 15388
rect 25682 15376 25688 15428
rect 25740 15416 25746 15428
rect 25838 15419 25896 15425
rect 25838 15416 25850 15419
rect 25740 15388 25850 15416
rect 25740 15376 25746 15388
rect 25838 15385 25850 15388
rect 25884 15385 25896 15419
rect 25838 15379 25896 15385
rect 28905 15419 28963 15425
rect 28905 15385 28917 15419
rect 28951 15416 28963 15419
rect 29178 15416 29184 15428
rect 28951 15388 29184 15416
rect 28951 15385 28963 15388
rect 28905 15379 28963 15385
rect 29178 15376 29184 15388
rect 29236 15376 29242 15428
rect 30190 15416 30196 15428
rect 30151 15388 30196 15416
rect 30190 15376 30196 15388
rect 30248 15376 30254 15428
rect 30650 15376 30656 15428
rect 30708 15416 30714 15428
rect 36354 15425 36360 15428
rect 31266 15419 31324 15425
rect 31266 15416 31278 15419
rect 30708 15388 31278 15416
rect 30708 15376 30714 15388
rect 31266 15385 31278 15388
rect 31312 15385 31324 15419
rect 31266 15379 31324 15385
rect 34885 15419 34943 15425
rect 34885 15385 34897 15419
rect 34931 15416 34943 15419
rect 36348 15416 36360 15425
rect 34931 15388 35388 15416
rect 36315 15388 36360 15416
rect 34931 15385 34943 15388
rect 34885 15379 34943 15385
rect 35360 15360 35388 15388
rect 36348 15379 36360 15388
rect 36354 15376 36360 15379
rect 36412 15376 36418 15428
rect 37826 15416 37832 15428
rect 37476 15388 37832 15416
rect 26050 15348 26056 15360
rect 25240 15320 26056 15348
rect 26050 15308 26056 15320
rect 26108 15348 26114 15360
rect 26973 15351 27031 15357
rect 26973 15348 26985 15351
rect 26108 15320 26985 15348
rect 26108 15308 26114 15320
rect 26973 15317 26985 15320
rect 27019 15348 27031 15351
rect 27338 15348 27344 15360
rect 27019 15320 27344 15348
rect 27019 15317 27031 15320
rect 26973 15311 27031 15317
rect 27338 15308 27344 15320
rect 27396 15308 27402 15360
rect 28074 15308 28080 15360
rect 28132 15348 28138 15360
rect 28997 15351 29055 15357
rect 28997 15348 29009 15351
rect 28132 15320 29009 15348
rect 28132 15308 28138 15320
rect 28997 15317 29009 15320
rect 29043 15317 29055 15351
rect 28997 15311 29055 15317
rect 32490 15308 32496 15360
rect 32548 15348 32554 15360
rect 34149 15351 34207 15357
rect 34149 15348 34161 15351
rect 32548 15320 34161 15348
rect 32548 15308 32554 15320
rect 34149 15317 34161 15320
rect 34195 15317 34207 15351
rect 34149 15311 34207 15317
rect 35342 15308 35348 15360
rect 35400 15308 35406 15360
rect 35618 15308 35624 15360
rect 35676 15348 35682 15360
rect 37476 15357 37504 15388
rect 37826 15376 37832 15388
rect 37884 15376 37890 15428
rect 38289 15419 38347 15425
rect 38289 15385 38301 15419
rect 38335 15416 38347 15419
rect 38562 15416 38568 15428
rect 38335 15388 38568 15416
rect 38335 15385 38347 15388
rect 38289 15379 38347 15385
rect 38562 15376 38568 15388
rect 38620 15376 38626 15428
rect 41325 15419 41383 15425
rect 41325 15385 41337 15419
rect 41371 15416 41383 15419
rect 41690 15416 41696 15428
rect 41371 15388 41696 15416
rect 41371 15385 41383 15388
rect 41325 15379 41383 15385
rect 41690 15376 41696 15388
rect 41748 15416 41754 15428
rect 41969 15419 42027 15425
rect 41969 15416 41981 15419
rect 41748 15388 41981 15416
rect 41748 15376 41754 15388
rect 41969 15385 41981 15388
rect 42015 15385 42027 15419
rect 41969 15379 42027 15385
rect 37461 15351 37519 15357
rect 37461 15348 37473 15351
rect 35676 15320 37473 15348
rect 35676 15308 35682 15320
rect 37461 15317 37473 15320
rect 37507 15317 37519 15351
rect 37461 15311 37519 15317
rect 37550 15308 37556 15360
rect 37608 15348 37614 15360
rect 37921 15351 37979 15357
rect 37921 15348 37933 15351
rect 37608 15320 37933 15348
rect 37608 15308 37614 15320
rect 37921 15317 37933 15320
rect 37967 15317 37979 15351
rect 37921 15311 37979 15317
rect 41506 15308 41512 15360
rect 41564 15348 41570 15360
rect 42426 15348 42432 15360
rect 41564 15320 42432 15348
rect 41564 15308 41570 15320
rect 42426 15308 42432 15320
rect 42484 15308 42490 15360
rect 42536 15348 42564 15592
rect 45388 15592 45784 15620
rect 47121 15623 47179 15629
rect 45388 15496 45416 15592
rect 47121 15589 47133 15623
rect 47167 15589 47179 15623
rect 49326 15620 49332 15632
rect 47121 15583 47179 15589
rect 48516 15592 49332 15620
rect 45738 15552 45744 15564
rect 45699 15524 45744 15552
rect 45738 15512 45744 15524
rect 45796 15512 45802 15564
rect 42702 15484 42708 15496
rect 42663 15456 42708 15484
rect 42702 15444 42708 15456
rect 42760 15444 42766 15496
rect 45094 15484 45100 15496
rect 45055 15456 45100 15484
rect 45094 15444 45100 15456
rect 45152 15444 45158 15496
rect 45189 15487 45247 15493
rect 45189 15453 45201 15487
rect 45235 15484 45247 15487
rect 45370 15484 45376 15496
rect 45235 15456 45376 15484
rect 45235 15453 45247 15456
rect 45189 15447 45247 15453
rect 45370 15444 45376 15456
rect 45428 15444 45434 15496
rect 45646 15444 45652 15496
rect 45704 15484 45710 15496
rect 45997 15487 46055 15493
rect 45997 15484 46009 15487
rect 45704 15456 46009 15484
rect 45704 15444 45710 15456
rect 45997 15453 46009 15456
rect 46043 15453 46055 15487
rect 45997 15447 46055 15453
rect 42972 15419 43030 15425
rect 42972 15385 42984 15419
rect 43018 15416 43030 15419
rect 44082 15416 44088 15428
rect 43018 15388 44088 15416
rect 43018 15385 43030 15388
rect 42972 15379 43030 15385
rect 44082 15376 44088 15388
rect 44140 15376 44146 15428
rect 47136 15416 47164 15583
rect 47486 15512 47492 15564
rect 47544 15552 47550 15564
rect 48317 15555 48375 15561
rect 47544 15524 48084 15552
rect 47544 15512 47550 15524
rect 47670 15444 47676 15496
rect 47728 15484 47734 15496
rect 47949 15487 48007 15493
rect 47728 15456 47773 15484
rect 47728 15444 47734 15456
rect 47949 15453 47961 15487
rect 47995 15453 48007 15487
rect 48056 15484 48084 15524
rect 48317 15521 48329 15555
rect 48363 15552 48375 15555
rect 48516 15552 48544 15592
rect 49326 15580 49332 15592
rect 49384 15580 49390 15632
rect 49418 15580 49424 15632
rect 49476 15620 49482 15632
rect 53098 15620 53104 15632
rect 49476 15592 53104 15620
rect 49476 15580 49482 15592
rect 53098 15580 53104 15592
rect 53156 15580 53162 15632
rect 54110 15620 54116 15632
rect 53484 15592 54116 15620
rect 53484 15561 53512 15592
rect 54110 15580 54116 15592
rect 54168 15580 54174 15632
rect 55398 15580 55404 15632
rect 55456 15620 55462 15632
rect 58342 15620 58348 15632
rect 55456 15592 58348 15620
rect 55456 15580 55462 15592
rect 58342 15580 58348 15592
rect 58400 15580 58406 15632
rect 48363 15524 48544 15552
rect 53469 15555 53527 15561
rect 48363 15521 48375 15524
rect 48317 15515 48375 15521
rect 53469 15521 53481 15555
rect 53515 15521 53527 15555
rect 53742 15552 53748 15564
rect 53703 15524 53748 15552
rect 53469 15515 53527 15521
rect 53742 15512 53748 15524
rect 53800 15512 53806 15564
rect 58158 15552 58164 15564
rect 55600 15524 58164 15552
rect 48501 15487 48559 15493
rect 48056 15456 48452 15484
rect 47949 15447 48007 15453
rect 47857 15419 47915 15425
rect 47857 15416 47869 15419
rect 47136 15388 47869 15416
rect 47857 15385 47869 15388
rect 47903 15385 47915 15419
rect 47857 15379 47915 15385
rect 47964 15416 47992 15447
rect 48268 15416 48274 15428
rect 47964 15388 48274 15416
rect 44266 15348 44272 15360
rect 42536 15320 44272 15348
rect 44266 15308 44272 15320
rect 44324 15308 44330 15360
rect 44358 15308 44364 15360
rect 44416 15348 44422 15360
rect 45094 15348 45100 15360
rect 44416 15320 45100 15348
rect 44416 15308 44422 15320
rect 45094 15308 45100 15320
rect 45152 15348 45158 15360
rect 45830 15348 45836 15360
rect 45152 15320 45836 15348
rect 45152 15308 45158 15320
rect 45830 15308 45836 15320
rect 45888 15308 45894 15360
rect 45922 15308 45928 15360
rect 45980 15348 45986 15360
rect 47964 15348 47992 15388
rect 48268 15376 48274 15388
rect 48326 15376 48332 15428
rect 48424 15416 48452 15456
rect 48501 15453 48513 15487
rect 48547 15484 48559 15487
rect 48682 15484 48688 15496
rect 48547 15456 48688 15484
rect 48547 15453 48563 15456
rect 48501 15452 48563 15453
rect 48501 15447 48559 15452
rect 48682 15444 48688 15456
rect 48740 15444 48746 15496
rect 48777 15487 48835 15493
rect 48777 15453 48789 15487
rect 48823 15453 48835 15487
rect 48777 15447 48835 15453
rect 49237 15487 49295 15493
rect 49237 15453 49249 15487
rect 49283 15484 49295 15487
rect 50246 15484 50252 15496
rect 49283 15456 50252 15484
rect 49283 15453 49295 15456
rect 49237 15447 49295 15453
rect 48792 15416 48820 15447
rect 50246 15444 50252 15456
rect 50304 15444 50310 15496
rect 50433 15487 50491 15493
rect 50433 15453 50445 15487
rect 50479 15484 50491 15487
rect 51074 15484 51080 15496
rect 50479 15456 51080 15484
rect 50479 15453 50491 15456
rect 50433 15447 50491 15453
rect 51074 15444 51080 15456
rect 51132 15444 51138 15496
rect 51258 15484 51264 15496
rect 51219 15456 51264 15484
rect 51258 15444 51264 15456
rect 51316 15444 51322 15496
rect 51442 15444 51448 15496
rect 51500 15484 51506 15496
rect 51629 15487 51687 15493
rect 51629 15484 51641 15487
rect 51500 15456 51641 15484
rect 51500 15444 51506 15456
rect 51629 15453 51641 15456
rect 51675 15453 51687 15487
rect 51902 15484 51908 15496
rect 51863 15456 51908 15484
rect 51629 15447 51687 15453
rect 51902 15444 51908 15456
rect 51960 15444 51966 15496
rect 52270 15484 52276 15496
rect 52231 15456 52276 15484
rect 52270 15444 52276 15456
rect 52328 15444 52334 15496
rect 52546 15484 52552 15496
rect 52507 15456 52552 15484
rect 52546 15444 52552 15456
rect 52604 15484 52610 15496
rect 53282 15484 53288 15496
rect 52604 15456 53288 15484
rect 52604 15444 52610 15456
rect 53282 15444 53288 15456
rect 53340 15484 53346 15496
rect 55600 15493 55628 15524
rect 58158 15512 58164 15524
rect 58216 15512 58222 15564
rect 58250 15512 58256 15564
rect 58308 15552 58314 15564
rect 58308 15524 58353 15552
rect 58308 15512 58314 15524
rect 55309 15487 55367 15493
rect 55309 15484 55321 15487
rect 53340 15456 55321 15484
rect 53340 15444 53346 15456
rect 55309 15453 55321 15456
rect 55355 15453 55367 15487
rect 55309 15447 55367 15453
rect 55585 15487 55643 15493
rect 55585 15453 55597 15487
rect 55631 15453 55643 15487
rect 55585 15447 55643 15453
rect 55674 15444 55680 15496
rect 55732 15484 55738 15496
rect 55953 15487 56011 15493
rect 55953 15484 55965 15487
rect 55732 15456 55965 15484
rect 55732 15444 55738 15456
rect 55953 15453 55965 15456
rect 55999 15453 56011 15487
rect 56226 15484 56232 15496
rect 56139 15456 56232 15484
rect 55953 15447 56011 15453
rect 56226 15444 56232 15456
rect 56284 15484 56290 15496
rect 56502 15484 56508 15496
rect 56284 15456 56508 15484
rect 56284 15444 56290 15456
rect 56502 15444 56508 15456
rect 56560 15444 56566 15496
rect 57514 15444 57520 15496
rect 57572 15484 57578 15496
rect 57885 15487 57943 15493
rect 57885 15484 57897 15487
rect 57572 15456 57897 15484
rect 57572 15444 57578 15456
rect 57885 15453 57897 15456
rect 57931 15453 57943 15487
rect 57885 15447 57943 15453
rect 58069 15487 58127 15493
rect 58069 15453 58081 15487
rect 58115 15484 58127 15487
rect 58452 15484 58480 15660
rect 58986 15648 58992 15660
rect 59044 15648 59050 15700
rect 59998 15688 60004 15700
rect 59959 15660 60004 15688
rect 59998 15648 60004 15660
rect 60056 15648 60062 15700
rect 60274 15648 60280 15700
rect 60332 15648 60338 15700
rect 60826 15648 60832 15700
rect 60884 15688 60890 15700
rect 65610 15688 65616 15700
rect 60884 15660 64644 15688
rect 65571 15660 65616 15688
rect 60884 15648 60890 15660
rect 60292 15620 60320 15648
rect 60292 15592 60872 15620
rect 58618 15552 58624 15564
rect 58579 15524 58624 15552
rect 58618 15512 58624 15524
rect 58676 15512 58682 15564
rect 60274 15512 60280 15564
rect 60332 15552 60338 15564
rect 60844 15561 60872 15592
rect 62390 15580 62396 15632
rect 62448 15620 62454 15632
rect 62850 15620 62856 15632
rect 62448 15592 62856 15620
rect 62448 15580 62454 15592
rect 62850 15580 62856 15592
rect 62908 15580 62914 15632
rect 64616 15620 64644 15660
rect 65610 15648 65616 15660
rect 65668 15648 65674 15700
rect 70765 15691 70823 15697
rect 70765 15688 70777 15691
rect 68940 15660 70777 15688
rect 68465 15623 68523 15629
rect 68465 15620 68477 15623
rect 64616 15592 68477 15620
rect 68465 15589 68477 15592
rect 68511 15589 68523 15623
rect 68465 15583 68523 15589
rect 60553 15555 60611 15561
rect 60553 15552 60565 15555
rect 60332 15524 60565 15552
rect 60332 15512 60338 15524
rect 60553 15521 60565 15524
rect 60599 15521 60611 15555
rect 60553 15515 60611 15521
rect 60829 15555 60887 15561
rect 60829 15521 60841 15555
rect 60875 15552 60887 15555
rect 62574 15552 62580 15564
rect 60875 15524 62580 15552
rect 60875 15521 60887 15524
rect 60829 15515 60887 15521
rect 62574 15512 62580 15524
rect 62632 15512 62638 15564
rect 62666 15512 62672 15564
rect 62724 15552 62730 15564
rect 62945 15555 63003 15561
rect 62945 15552 62957 15555
rect 62724 15524 62957 15552
rect 62724 15512 62730 15524
rect 62945 15521 62957 15524
rect 62991 15521 63003 15555
rect 62945 15515 63003 15521
rect 64138 15512 64144 15564
rect 64196 15552 64202 15564
rect 65334 15552 65340 15564
rect 64196 15524 65340 15552
rect 64196 15512 64202 15524
rect 65334 15512 65340 15524
rect 65392 15552 65398 15564
rect 67266 15552 67272 15564
rect 65392 15524 67272 15552
rect 65392 15512 65398 15524
rect 58115 15456 58480 15484
rect 58115 15453 58127 15456
rect 58069 15447 58127 15453
rect 58710 15444 58716 15496
rect 58768 15484 58774 15496
rect 60366 15484 60372 15496
rect 58768 15456 60372 15484
rect 58768 15444 58774 15456
rect 60366 15444 60372 15456
rect 60424 15444 60430 15496
rect 62025 15487 62083 15493
rect 62025 15453 62037 15487
rect 62071 15484 62083 15487
rect 63034 15484 63040 15496
rect 62071 15456 63040 15484
rect 62071 15453 62083 15456
rect 62025 15447 62083 15453
rect 63034 15444 63040 15456
rect 63092 15444 63098 15496
rect 63212 15487 63270 15493
rect 63212 15453 63224 15487
rect 63258 15484 63270 15487
rect 63770 15484 63776 15496
rect 63258 15456 63776 15484
rect 63258 15453 63270 15456
rect 63212 15447 63270 15453
rect 63770 15444 63776 15456
rect 63828 15444 63834 15496
rect 64874 15484 64880 15496
rect 64835 15456 64880 15484
rect 64874 15444 64880 15456
rect 64932 15444 64938 15496
rect 65242 15444 65248 15496
rect 65300 15484 65306 15496
rect 65794 15484 65800 15496
rect 65300 15456 65800 15484
rect 65300 15444 65306 15456
rect 65794 15444 65800 15456
rect 65852 15444 65858 15496
rect 65996 15493 66024 15524
rect 67266 15512 67272 15524
rect 67324 15512 67330 15564
rect 68940 15552 68968 15660
rect 70765 15657 70777 15660
rect 70811 15657 70823 15691
rect 71866 15688 71872 15700
rect 71827 15660 71872 15688
rect 70765 15651 70823 15657
rect 71866 15648 71872 15660
rect 71924 15648 71930 15700
rect 69934 15580 69940 15632
rect 69992 15620 69998 15632
rect 72513 15623 72571 15629
rect 72513 15620 72525 15623
rect 69992 15592 72525 15620
rect 69992 15580 69998 15592
rect 72513 15589 72525 15592
rect 72559 15589 72571 15623
rect 72513 15583 72571 15589
rect 71222 15552 71228 15564
rect 68020 15524 68968 15552
rect 71183 15524 71228 15552
rect 68020 15493 68048 15524
rect 71222 15512 71228 15524
rect 71280 15512 71286 15564
rect 71409 15555 71467 15561
rect 71409 15521 71421 15555
rect 71455 15552 71467 15555
rect 71498 15552 71504 15564
rect 71455 15524 71504 15552
rect 71455 15521 71467 15524
rect 71409 15515 71467 15521
rect 71498 15512 71504 15524
rect 71556 15512 71562 15564
rect 65981 15487 66039 15493
rect 65981 15453 65993 15487
rect 66027 15453 66039 15487
rect 65981 15447 66039 15453
rect 66073 15487 66131 15493
rect 66073 15453 66085 15487
rect 66119 15453 66131 15487
rect 66073 15447 66131 15453
rect 68005 15487 68063 15493
rect 68005 15453 68017 15487
rect 68051 15453 68063 15487
rect 68005 15447 68063 15453
rect 68373 15487 68431 15493
rect 68373 15453 68385 15487
rect 68419 15480 68431 15487
rect 68922 15484 68928 15496
rect 68419 15453 68508 15480
rect 68883 15456 68928 15484
rect 68373 15452 68508 15453
rect 68373 15447 68431 15452
rect 48424 15388 48820 15416
rect 50154 15376 50160 15428
rect 50212 15416 50218 15428
rect 50212 15388 50257 15416
rect 50212 15376 50218 15388
rect 50798 15376 50804 15428
rect 50856 15416 50862 15428
rect 51813 15419 51871 15425
rect 50856 15388 51764 15416
rect 50856 15376 50862 15388
rect 45980 15320 47992 15348
rect 45980 15308 45986 15320
rect 48038 15308 48044 15360
rect 48096 15348 48102 15360
rect 48685 15351 48743 15357
rect 48685 15348 48697 15351
rect 48096 15320 48697 15348
rect 48096 15308 48102 15320
rect 48685 15317 48697 15320
rect 48731 15348 48743 15351
rect 49694 15348 49700 15360
rect 48731 15320 49700 15348
rect 48731 15317 48743 15320
rect 48685 15311 48743 15317
rect 49694 15308 49700 15320
rect 49752 15308 49758 15360
rect 49970 15308 49976 15360
rect 50028 15348 50034 15360
rect 50341 15351 50399 15357
rect 50341 15348 50353 15351
rect 50028 15320 50353 15348
rect 50028 15308 50034 15320
rect 50341 15317 50353 15320
rect 50387 15317 50399 15351
rect 50341 15311 50399 15317
rect 50430 15308 50436 15360
rect 50488 15348 50494 15360
rect 51077 15351 51135 15357
rect 51077 15348 51089 15351
rect 50488 15320 51089 15348
rect 50488 15308 50494 15320
rect 51077 15317 51089 15320
rect 51123 15317 51135 15351
rect 51736 15348 51764 15388
rect 51813 15385 51825 15419
rect 51859 15416 51871 15419
rect 51994 15416 52000 15428
rect 51859 15388 52000 15416
rect 51859 15385 51871 15388
rect 51813 15379 51871 15385
rect 51994 15376 52000 15388
rect 52052 15416 52058 15428
rect 53558 15416 53564 15428
rect 52052 15388 53564 15416
rect 52052 15376 52058 15388
rect 53558 15376 53564 15388
rect 53616 15416 53622 15428
rect 53742 15416 53748 15428
rect 53616 15388 53748 15416
rect 53616 15376 53622 15388
rect 53742 15376 53748 15388
rect 53800 15376 53806 15428
rect 55122 15416 55128 15428
rect 54680 15388 55128 15416
rect 54680 15348 54708 15388
rect 55122 15376 55128 15388
rect 55180 15376 55186 15428
rect 55493 15419 55551 15425
rect 55493 15416 55505 15419
rect 55324 15388 55505 15416
rect 51736 15320 54708 15348
rect 51077 15311 51135 15317
rect 54754 15308 54760 15360
rect 54812 15348 54818 15360
rect 55324 15348 55352 15388
rect 55493 15385 55505 15388
rect 55539 15385 55551 15419
rect 55493 15379 55551 15385
rect 56778 15376 56784 15428
rect 56836 15416 56842 15428
rect 57241 15419 57299 15425
rect 57241 15416 57253 15419
rect 56836 15388 57253 15416
rect 56836 15376 56842 15388
rect 57241 15385 57253 15388
rect 57287 15385 57299 15419
rect 57241 15379 57299 15385
rect 57974 15376 57980 15428
rect 58032 15416 58038 15428
rect 58866 15419 58924 15425
rect 58866 15416 58878 15419
rect 58032 15388 58878 15416
rect 58032 15376 58038 15388
rect 58866 15385 58878 15388
rect 58912 15385 58924 15419
rect 61838 15416 61844 15428
rect 61799 15388 61844 15416
rect 58866 15379 58924 15385
rect 61838 15376 61844 15388
rect 61896 15376 61902 15428
rect 62301 15419 62359 15425
rect 62301 15416 62313 15419
rect 61948 15388 62313 15416
rect 54812 15320 55352 15348
rect 54812 15308 54818 15320
rect 55398 15308 55404 15360
rect 55456 15348 55462 15360
rect 57330 15348 57336 15360
rect 55456 15320 57336 15348
rect 55456 15308 55462 15320
rect 57330 15308 57336 15320
rect 57388 15308 57394 15360
rect 57422 15308 57428 15360
rect 57480 15348 57486 15360
rect 60550 15348 60556 15360
rect 57480 15320 60556 15348
rect 57480 15308 57486 15320
rect 60550 15308 60556 15320
rect 60608 15308 60614 15360
rect 60918 15308 60924 15360
rect 60976 15348 60982 15360
rect 61948 15348 61976 15388
rect 62301 15385 62313 15388
rect 62347 15385 62359 15419
rect 62301 15379 62359 15385
rect 62390 15376 62396 15428
rect 62448 15416 62454 15428
rect 66088 15416 66116 15447
rect 62448 15388 66116 15416
rect 62448 15376 62454 15388
rect 60976 15320 61976 15348
rect 60976 15308 60982 15320
rect 62114 15308 62120 15360
rect 62172 15348 62178 15360
rect 62209 15351 62267 15357
rect 62209 15348 62221 15351
rect 62172 15320 62221 15348
rect 62172 15308 62178 15320
rect 62209 15317 62221 15320
rect 62255 15348 62267 15351
rect 62666 15348 62672 15360
rect 62255 15320 62672 15348
rect 62255 15317 62267 15320
rect 62209 15311 62267 15317
rect 62666 15308 62672 15320
rect 62724 15348 62730 15360
rect 64138 15348 64144 15360
rect 62724 15320 64144 15348
rect 62724 15308 62730 15320
rect 64138 15308 64144 15320
rect 64196 15308 64202 15360
rect 64322 15348 64328 15360
rect 64283 15320 64328 15348
rect 64322 15308 64328 15320
rect 64380 15308 64386 15360
rect 64598 15308 64604 15360
rect 64656 15348 64662 15360
rect 64693 15351 64751 15357
rect 64693 15348 64705 15351
rect 64656 15320 64705 15348
rect 64656 15308 64662 15320
rect 64693 15317 64705 15320
rect 64739 15317 64751 15351
rect 67818 15348 67824 15360
rect 67779 15320 67824 15348
rect 64693 15311 64751 15317
rect 67818 15308 67824 15320
rect 67876 15308 67882 15360
rect 68480 15348 68508 15452
rect 68922 15444 68928 15456
rect 68980 15444 68986 15496
rect 69192 15487 69250 15493
rect 69192 15453 69204 15487
rect 69238 15484 69250 15487
rect 70118 15484 70124 15496
rect 69238 15456 70124 15484
rect 69238 15453 69250 15456
rect 69192 15447 69250 15453
rect 70118 15444 70124 15456
rect 70176 15444 70182 15496
rect 72050 15484 72056 15496
rect 72011 15456 72056 15484
rect 72050 15444 72056 15456
rect 72108 15444 72114 15496
rect 72418 15484 72424 15496
rect 72379 15456 72424 15484
rect 72418 15444 72424 15456
rect 72476 15444 72482 15496
rect 88058 15416 88064 15428
rect 88019 15388 88064 15416
rect 88058 15376 88064 15388
rect 88116 15376 88122 15428
rect 70302 15348 70308 15360
rect 68480 15320 70308 15348
rect 70302 15308 70308 15320
rect 70360 15308 70366 15360
rect 70394 15308 70400 15360
rect 70452 15348 70458 15360
rect 71133 15351 71191 15357
rect 71133 15348 71145 15351
rect 70452 15320 71145 15348
rect 70452 15308 70458 15320
rect 71133 15317 71145 15320
rect 71179 15317 71191 15351
rect 88150 15348 88156 15360
rect 88111 15320 88156 15348
rect 71133 15311 71191 15317
rect 88150 15308 88156 15320
rect 88208 15308 88214 15360
rect 1104 15258 88872 15280
rect 1104 15206 22898 15258
rect 22950 15206 22962 15258
rect 23014 15206 23026 15258
rect 23078 15206 23090 15258
rect 23142 15206 23154 15258
rect 23206 15206 44846 15258
rect 44898 15206 44910 15258
rect 44962 15206 44974 15258
rect 45026 15206 45038 15258
rect 45090 15206 45102 15258
rect 45154 15206 66794 15258
rect 66846 15206 66858 15258
rect 66910 15206 66922 15258
rect 66974 15206 66986 15258
rect 67038 15206 67050 15258
rect 67102 15206 88872 15258
rect 1104 15184 88872 15206
rect 11698 15104 11704 15156
rect 11756 15144 11762 15156
rect 11756 15116 12434 15144
rect 11756 15104 11762 15116
rect 12406 15076 12434 15116
rect 16482 15104 16488 15156
rect 16540 15144 16546 15156
rect 18601 15147 18659 15153
rect 18601 15144 18613 15147
rect 16540 15116 18613 15144
rect 16540 15104 16546 15116
rect 18601 15113 18613 15116
rect 18647 15113 18659 15147
rect 18601 15107 18659 15113
rect 19886 15104 19892 15156
rect 19944 15144 19950 15156
rect 20073 15147 20131 15153
rect 20073 15144 20085 15147
rect 19944 15116 20085 15144
rect 19944 15104 19950 15116
rect 20073 15113 20085 15116
rect 20119 15113 20131 15147
rect 20073 15107 20131 15113
rect 20441 15147 20499 15153
rect 20441 15113 20453 15147
rect 20487 15144 20499 15147
rect 20714 15144 20720 15156
rect 20487 15116 20720 15144
rect 20487 15113 20499 15116
rect 20441 15107 20499 15113
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 20898 15144 20904 15156
rect 20824 15116 20904 15144
rect 12710 15076 12716 15088
rect 12406 15048 12716 15076
rect 12710 15036 12716 15048
rect 12768 15076 12774 15088
rect 20824 15076 20852 15116
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 22094 15144 22100 15156
rect 22066 15104 22100 15144
rect 22152 15104 22158 15156
rect 22281 15147 22339 15153
rect 22281 15113 22293 15147
rect 22327 15144 22339 15147
rect 22462 15144 22468 15156
rect 22327 15116 22468 15144
rect 22327 15113 22339 15116
rect 22281 15107 22339 15113
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 22572 15116 24072 15144
rect 22066 15076 22094 15104
rect 12768 15048 19104 15076
rect 12768 15036 12774 15048
rect 19076 15020 19104 15048
rect 20272 15048 20852 15076
rect 20916 15048 22094 15076
rect 18782 15008 18788 15020
rect 18743 14980 18788 15008
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 18966 15008 18972 15020
rect 18927 14980 18972 15008
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 19058 14968 19064 15020
rect 19116 15008 19122 15020
rect 20272 15017 20300 15048
rect 20916 15017 20944 15048
rect 20257 15011 20315 15017
rect 19116 14980 19161 15008
rect 19116 14968 19122 14980
rect 20257 14977 20269 15011
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20533 15011 20591 15017
rect 20533 14977 20545 15011
rect 20579 14977 20591 15011
rect 20533 14971 20591 14977
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 20548 14872 20576 14971
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22097 15011 22155 15017
rect 22097 15008 22109 15011
rect 22060 14980 22109 15008
rect 22060 14968 22066 14980
rect 22097 14977 22109 14980
rect 22143 14977 22155 15011
rect 22370 15008 22376 15020
rect 22283 14980 22376 15008
rect 22097 14971 22155 14977
rect 22370 14968 22376 14980
rect 22428 15008 22434 15020
rect 22572 15008 22600 15116
rect 23382 15036 23388 15088
rect 23440 15076 23446 15088
rect 23937 15079 23995 15085
rect 23937 15076 23949 15079
rect 23440 15048 23949 15076
rect 23440 15036 23446 15048
rect 23937 15045 23949 15048
rect 23983 15045 23995 15079
rect 24044 15076 24072 15116
rect 24302 15104 24308 15156
rect 24360 15144 24366 15156
rect 24854 15144 24860 15156
rect 24360 15116 24860 15144
rect 24360 15104 24366 15116
rect 24854 15104 24860 15116
rect 24912 15144 24918 15156
rect 25498 15144 25504 15156
rect 24912 15116 25504 15144
rect 24912 15104 24918 15116
rect 25498 15104 25504 15116
rect 25556 15104 25562 15156
rect 25590 15104 25596 15156
rect 25648 15144 25654 15156
rect 25648 15116 27272 15144
rect 25648 15104 25654 15116
rect 24670 15076 24676 15088
rect 24044 15048 24676 15076
rect 23937 15039 23995 15045
rect 24670 15036 24676 15048
rect 24728 15036 24734 15088
rect 27244 15076 27272 15116
rect 27338 15104 27344 15156
rect 27396 15144 27402 15156
rect 27433 15147 27491 15153
rect 27433 15144 27445 15147
rect 27396 15116 27445 15144
rect 27396 15104 27402 15116
rect 27433 15113 27445 15116
rect 27479 15113 27491 15147
rect 27433 15107 27491 15113
rect 27522 15104 27528 15156
rect 27580 15144 27586 15156
rect 30469 15147 30527 15153
rect 27580 15116 28856 15144
rect 27580 15104 27586 15116
rect 28828 15085 28856 15116
rect 30469 15113 30481 15147
rect 30515 15144 30527 15147
rect 31938 15144 31944 15156
rect 30515 15116 31944 15144
rect 30515 15113 30527 15116
rect 30469 15107 30527 15113
rect 31938 15104 31944 15116
rect 31996 15104 32002 15156
rect 32122 15144 32128 15156
rect 32083 15116 32128 15144
rect 32122 15104 32128 15116
rect 32180 15104 32186 15156
rect 32306 15104 32312 15156
rect 32364 15144 32370 15156
rect 32585 15147 32643 15153
rect 32585 15144 32597 15147
rect 32364 15116 32597 15144
rect 32364 15104 32370 15116
rect 32585 15113 32597 15116
rect 32631 15113 32643 15147
rect 33226 15144 33232 15156
rect 33187 15116 33232 15144
rect 32585 15107 32643 15113
rect 33226 15104 33232 15116
rect 33284 15104 33290 15156
rect 33318 15104 33324 15156
rect 33376 15144 33382 15156
rect 33597 15147 33655 15153
rect 33597 15144 33609 15147
rect 33376 15116 33609 15144
rect 33376 15104 33382 15116
rect 33597 15113 33609 15116
rect 33643 15144 33655 15147
rect 41506 15144 41512 15156
rect 33643 15116 35664 15144
rect 33643 15113 33655 15116
rect 33597 15107 33655 15113
rect 28721 15079 28779 15085
rect 28721 15076 28733 15079
rect 27244 15048 28733 15076
rect 22738 15008 22744 15020
rect 22428 14980 22600 15008
rect 22699 14980 22744 15008
rect 22428 14968 22434 14980
rect 22738 14968 22744 14980
rect 22796 14968 22802 15020
rect 23290 14968 23296 15020
rect 23348 15006 23354 15020
rect 23661 15011 23719 15017
rect 23661 15008 23673 15011
rect 23400 15006 23673 15008
rect 23348 14980 23673 15006
rect 23348 14978 23428 14980
rect 23348 14968 23354 14978
rect 23661 14977 23673 14980
rect 23707 14977 23719 15011
rect 23661 14971 23719 14977
rect 23753 15011 23811 15017
rect 23753 14977 23765 15011
rect 23799 15008 23811 15011
rect 24210 15008 24216 15020
rect 23799 14980 24216 15008
rect 23799 14977 23811 14980
rect 23753 14971 23811 14977
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 21913 14943 21971 14949
rect 21913 14940 21925 14943
rect 20680 14912 21925 14940
rect 20680 14900 20686 14912
rect 21913 14909 21925 14912
rect 21959 14909 21971 14943
rect 23676 14940 23704 14971
rect 24210 14968 24216 14980
rect 24268 14968 24274 15020
rect 24302 14968 24308 15020
rect 24360 15008 24366 15020
rect 24489 15011 24547 15017
rect 24360 14980 24405 15008
rect 24360 14968 24366 14980
rect 24489 14977 24501 15011
rect 24535 14977 24547 15011
rect 25038 15008 25044 15020
rect 24999 14980 25044 15008
rect 24489 14971 24547 14977
rect 24118 14940 24124 14952
rect 23676 14912 24124 14940
rect 21913 14903 21971 14909
rect 24118 14900 24124 14912
rect 24176 14900 24182 14952
rect 24394 14900 24400 14952
rect 24452 14940 24458 14952
rect 24504 14940 24532 14971
rect 25038 14968 25044 14980
rect 25096 14968 25102 15020
rect 25130 14968 25136 15020
rect 25188 15008 25194 15020
rect 25297 15011 25355 15017
rect 25297 15008 25309 15011
rect 25188 14980 25309 15008
rect 25188 14968 25194 14980
rect 25297 14977 25309 14980
rect 25343 14977 25355 15011
rect 25297 14971 25355 14977
rect 26510 14968 26516 15020
rect 26568 15008 26574 15020
rect 27246 15008 27252 15020
rect 26568 14980 27252 15008
rect 26568 14968 26574 14980
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 15008 27399 15011
rect 27706 15008 27712 15020
rect 27387 14980 27712 15008
rect 27387 14977 27399 14980
rect 27341 14971 27399 14977
rect 24452 14912 24532 14940
rect 24452 14900 24458 14912
rect 26234 14900 26240 14952
rect 26292 14940 26298 14952
rect 26786 14940 26792 14952
rect 26292 14912 26792 14940
rect 26292 14900 26298 14912
rect 26786 14900 26792 14912
rect 26844 14900 26850 14952
rect 27356 14940 27384 14971
rect 27706 14968 27712 14980
rect 27764 14968 27770 15020
rect 27430 14940 27436 14952
rect 27356 14912 27436 14940
rect 27430 14900 27436 14912
rect 27488 14900 27494 14952
rect 27522 14900 27528 14952
rect 27580 14940 27586 14952
rect 28368 14940 28396 15048
rect 28721 15045 28733 15048
rect 28767 15045 28779 15079
rect 28721 15039 28779 15045
rect 28813 15079 28871 15085
rect 28813 15045 28825 15079
rect 28859 15045 28871 15079
rect 28813 15039 28871 15045
rect 28902 15036 28908 15088
rect 28960 15076 28966 15088
rect 32490 15076 32496 15088
rect 28960 15048 30236 15076
rect 28960 15036 28966 15048
rect 28534 15008 28540 15020
rect 28495 14980 28540 15008
rect 28534 14968 28540 14980
rect 28592 15008 28598 15020
rect 28994 15008 29000 15020
rect 28592 15006 28672 15008
rect 28736 15006 29000 15008
rect 28592 14980 29000 15006
rect 28592 14968 28598 14980
rect 28644 14978 28764 14980
rect 28994 14968 29000 14980
rect 29052 14968 29058 15020
rect 29178 15008 29184 15020
rect 29091 14980 29184 15008
rect 29178 14968 29184 14980
rect 29236 15008 29242 15020
rect 30098 15008 30104 15020
rect 29236 14980 30104 15008
rect 29236 14968 29242 14980
rect 30098 14968 30104 14980
rect 30156 14968 30162 15020
rect 28902 14940 28908 14952
rect 27580 14912 27625 14940
rect 28368 14912 28908 14940
rect 27580 14900 27586 14912
rect 28902 14900 28908 14912
rect 28960 14940 28966 14952
rect 29457 14943 29515 14949
rect 29457 14940 29469 14943
rect 28960 14912 29469 14940
rect 28960 14900 28966 14912
rect 29457 14909 29469 14912
rect 29503 14909 29515 14943
rect 30208 14940 30236 15048
rect 30392 15048 31432 15076
rect 32451 15048 32496 15076
rect 30392 15017 30420 15048
rect 30377 15011 30435 15017
rect 30377 14977 30389 15011
rect 30423 14977 30435 15011
rect 31294 15008 31300 15020
rect 31255 14980 31300 15008
rect 30377 14971 30435 14977
rect 31294 14968 31300 14980
rect 31352 14968 31358 15020
rect 31404 15008 31432 15048
rect 32490 15036 32496 15048
rect 32548 15036 32554 15088
rect 32674 15036 32680 15088
rect 32732 15076 32738 15088
rect 32732 15048 34100 15076
rect 32732 15036 32738 15048
rect 32508 15008 32536 15036
rect 31404 14980 32536 15008
rect 32582 14968 32588 15020
rect 32640 15008 32646 15020
rect 33413 15011 33471 15017
rect 32640 14980 33180 15008
rect 32640 14968 32646 14980
rect 31389 14943 31447 14949
rect 31389 14940 31401 14943
rect 30208 14912 31401 14940
rect 29457 14903 29515 14909
rect 31389 14909 31401 14912
rect 31435 14909 31447 14943
rect 31389 14903 31447 14909
rect 31573 14943 31631 14949
rect 31573 14909 31585 14943
rect 31619 14940 31631 14943
rect 32769 14943 32827 14949
rect 32769 14940 32781 14943
rect 31619 14912 32781 14940
rect 31619 14909 31631 14912
rect 31573 14903 31631 14909
rect 32769 14909 32781 14912
rect 32815 14909 32827 14943
rect 33152 14940 33180 14980
rect 33413 14977 33425 15011
rect 33459 15008 33471 15011
rect 33502 15008 33508 15020
rect 33459 14980 33508 15008
rect 33459 14977 33471 14980
rect 33413 14971 33471 14977
rect 33502 14968 33508 14980
rect 33560 14968 33566 15020
rect 33594 14968 33600 15020
rect 33652 15008 33658 15020
rect 33689 15011 33747 15017
rect 33689 15008 33701 15011
rect 33652 14980 33701 15008
rect 33652 14968 33658 14980
rect 33689 14977 33701 14980
rect 33735 15008 33747 15011
rect 33962 15008 33968 15020
rect 33735 14980 33968 15008
rect 33735 14977 33747 14980
rect 33689 14971 33747 14977
rect 33962 14968 33968 14980
rect 34020 14968 34026 15020
rect 34072 15017 34100 15048
rect 34238 15036 34244 15088
rect 34296 15076 34302 15088
rect 34296 15048 35480 15076
rect 34296 15036 34302 15048
rect 35452 15020 35480 15048
rect 34057 15011 34115 15017
rect 34057 14977 34069 15011
rect 34103 14977 34115 15011
rect 34609 15011 34667 15017
rect 34609 15008 34621 15011
rect 34057 14971 34115 14977
rect 34164 14980 34621 15008
rect 34164 14940 34192 14980
rect 34609 14977 34621 14980
rect 34655 14977 34667 15011
rect 35250 15008 35256 15020
rect 35211 14980 35256 15008
rect 34609 14971 34667 14977
rect 35250 14968 35256 14980
rect 35308 14968 35314 15020
rect 35434 15008 35440 15020
rect 35395 14980 35440 15008
rect 35434 14968 35440 14980
rect 35492 14968 35498 15020
rect 35529 15011 35587 15017
rect 35529 14977 35541 15011
rect 35575 14977 35587 15011
rect 35636 15008 35664 15116
rect 36004 15116 41512 15144
rect 36004 15085 36032 15116
rect 41506 15104 41512 15116
rect 41564 15104 41570 15156
rect 42426 15104 42432 15156
rect 42484 15144 42490 15156
rect 53098 15144 53104 15156
rect 42484 15116 53104 15144
rect 42484 15104 42490 15116
rect 53098 15104 53104 15116
rect 53156 15104 53162 15156
rect 53469 15147 53527 15153
rect 53469 15113 53481 15147
rect 53515 15144 53527 15147
rect 53515 15116 53696 15144
rect 53515 15113 53527 15116
rect 53469 15107 53527 15113
rect 35989 15079 36047 15085
rect 35989 15045 36001 15079
rect 36035 15045 36047 15079
rect 49688 15079 49746 15085
rect 35989 15039 36047 15045
rect 36096 15048 48820 15076
rect 36096 15008 36124 15048
rect 35636 14980 36124 15008
rect 35529 14971 35587 14977
rect 33152 14912 34192 14940
rect 32769 14903 32827 14909
rect 32784 14872 32812 14903
rect 34514 14900 34520 14952
rect 34572 14940 34578 14952
rect 35544 14940 35572 14971
rect 36170 14968 36176 15020
rect 36228 15008 36234 15020
rect 36357 15011 36415 15017
rect 36228 14980 36273 15008
rect 36228 14968 36234 14980
rect 36357 14977 36369 15011
rect 36403 14977 36415 15011
rect 36357 14971 36415 14977
rect 34572 14912 35572 14940
rect 34572 14900 34578 14912
rect 36262 14900 36268 14952
rect 36320 14940 36326 14952
rect 36372 14940 36400 14971
rect 36446 14968 36452 15020
rect 36504 15008 36510 15020
rect 36504 14980 36549 15008
rect 36504 14968 36510 14980
rect 37090 14968 37096 15020
rect 37148 15008 37154 15020
rect 37533 15011 37591 15017
rect 37533 15008 37545 15011
rect 37148 14980 37545 15008
rect 37148 14968 37154 14980
rect 37533 14977 37545 14980
rect 37579 14977 37591 15011
rect 37533 14971 37591 14977
rect 37826 14968 37832 15020
rect 37884 15008 37890 15020
rect 39649 15011 39707 15017
rect 39649 15008 39661 15011
rect 37884 14980 39661 15008
rect 37884 14968 37890 14980
rect 39649 14977 39661 14980
rect 39695 14977 39707 15011
rect 39649 14971 39707 14977
rect 39942 14968 39948 15020
rect 40000 15008 40006 15020
rect 41141 15011 41199 15017
rect 41141 15008 41153 15011
rect 40000 14980 41153 15008
rect 40000 14968 40006 14980
rect 41141 14977 41153 14980
rect 41187 14977 41199 15011
rect 41690 15008 41696 15020
rect 41603 14980 41696 15008
rect 41141 14971 41199 14977
rect 41690 14968 41696 14980
rect 41748 15008 41754 15020
rect 42429 15011 42487 15017
rect 42429 15008 42441 15011
rect 41748 14980 42441 15008
rect 41748 14968 41754 14980
rect 42429 14977 42441 14980
rect 42475 15008 42487 15011
rect 42475 14980 43300 15008
rect 42475 14977 42487 14980
rect 42429 14971 42487 14977
rect 37274 14940 37280 14952
rect 36320 14912 36400 14940
rect 37235 14912 37280 14940
rect 36320 14900 36326 14912
rect 37274 14900 37280 14912
rect 37332 14900 37338 14952
rect 39390 14940 39396 14952
rect 39351 14912 39396 14940
rect 39390 14900 39396 14912
rect 39448 14900 39454 14952
rect 41233 14943 41291 14949
rect 41233 14909 41245 14943
rect 41279 14940 41291 14943
rect 41279 14912 43024 14940
rect 41279 14909 41291 14912
rect 41233 14903 41291 14909
rect 20548 14844 25084 14872
rect 21174 14804 21180 14816
rect 21135 14776 21180 14804
rect 21174 14764 21180 14776
rect 21232 14764 21238 14816
rect 21358 14804 21364 14816
rect 21319 14776 21364 14804
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 22094 14764 22100 14816
rect 22152 14804 22158 14816
rect 23017 14807 23075 14813
rect 23017 14804 23029 14807
rect 22152 14776 23029 14804
rect 22152 14764 22158 14776
rect 23017 14773 23029 14776
rect 23063 14804 23075 14807
rect 23106 14804 23112 14816
rect 23063 14776 23112 14804
rect 23063 14773 23075 14776
rect 23017 14767 23075 14773
rect 23106 14764 23112 14776
rect 23164 14764 23170 14816
rect 23201 14807 23259 14813
rect 23201 14773 23213 14807
rect 23247 14804 23259 14807
rect 23842 14804 23848 14816
rect 23247 14776 23848 14804
rect 23247 14773 23259 14776
rect 23201 14767 23259 14773
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 24302 14804 24308 14816
rect 24263 14776 24308 14804
rect 24302 14764 24308 14776
rect 24360 14764 24366 14816
rect 25056 14804 25084 14844
rect 25976 14844 32444 14872
rect 32784 14844 36032 14872
rect 25976 14804 26004 14844
rect 26418 14804 26424 14816
rect 25056 14776 26004 14804
rect 26379 14776 26424 14804
rect 26418 14764 26424 14776
rect 26476 14764 26482 14816
rect 26510 14764 26516 14816
rect 26568 14804 26574 14816
rect 26973 14807 27031 14813
rect 26973 14804 26985 14807
rect 26568 14776 26985 14804
rect 26568 14764 26574 14776
rect 26973 14773 26985 14776
rect 27019 14773 27031 14807
rect 26973 14767 27031 14773
rect 27062 14764 27068 14816
rect 27120 14804 27126 14816
rect 27522 14804 27528 14816
rect 27120 14776 27528 14804
rect 27120 14764 27126 14776
rect 27522 14764 27528 14776
rect 27580 14764 27586 14816
rect 27982 14764 27988 14816
rect 28040 14804 28046 14816
rect 28353 14807 28411 14813
rect 28353 14804 28365 14807
rect 28040 14776 28365 14804
rect 28040 14764 28046 14776
rect 28353 14773 28365 14776
rect 28399 14773 28411 14807
rect 28353 14767 28411 14773
rect 28534 14764 28540 14816
rect 28592 14804 28598 14816
rect 30834 14804 30840 14816
rect 28592 14776 30840 14804
rect 28592 14764 28598 14776
rect 30834 14764 30840 14776
rect 30892 14764 30898 14816
rect 30929 14807 30987 14813
rect 30929 14773 30941 14807
rect 30975 14804 30987 14807
rect 31754 14804 31760 14816
rect 30975 14776 31760 14804
rect 30975 14773 30987 14776
rect 30929 14767 30987 14773
rect 31754 14764 31760 14776
rect 31812 14764 31818 14816
rect 31846 14764 31852 14816
rect 31904 14804 31910 14816
rect 32122 14804 32128 14816
rect 31904 14776 32128 14804
rect 31904 14764 31910 14776
rect 32122 14764 32128 14776
rect 32180 14764 32186 14816
rect 32416 14804 32444 14844
rect 33226 14804 33232 14816
rect 32416 14776 33232 14804
rect 33226 14764 33232 14776
rect 33284 14764 33290 14816
rect 34149 14807 34207 14813
rect 34149 14773 34161 14807
rect 34195 14804 34207 14807
rect 34514 14804 34520 14816
rect 34195 14776 34520 14804
rect 34195 14773 34207 14776
rect 34149 14767 34207 14773
rect 34514 14764 34520 14776
rect 34572 14764 34578 14816
rect 34698 14804 34704 14816
rect 34659 14776 34704 14804
rect 34698 14764 34704 14776
rect 34756 14764 34762 14816
rect 35253 14807 35311 14813
rect 35253 14773 35265 14807
rect 35299 14804 35311 14807
rect 35894 14804 35900 14816
rect 35299 14776 35900 14804
rect 35299 14773 35311 14776
rect 35253 14767 35311 14773
rect 35894 14764 35900 14776
rect 35952 14764 35958 14816
rect 36004 14804 36032 14844
rect 38203 14844 39436 14872
rect 38203 14804 38231 14844
rect 36004 14776 38231 14804
rect 38562 14764 38568 14816
rect 38620 14804 38626 14816
rect 38657 14807 38715 14813
rect 38657 14804 38669 14807
rect 38620 14776 38669 14804
rect 38620 14764 38626 14776
rect 38657 14773 38669 14776
rect 38703 14773 38715 14807
rect 39408 14804 39436 14844
rect 40328 14844 40908 14872
rect 40328 14804 40356 14844
rect 40770 14804 40776 14816
rect 39408 14776 40356 14804
rect 40731 14776 40776 14804
rect 38657 14767 38715 14773
rect 40770 14764 40776 14776
rect 40828 14764 40834 14816
rect 40880 14804 40908 14844
rect 41782 14832 41788 14884
rect 41840 14872 41846 14884
rect 41877 14875 41935 14881
rect 41877 14872 41889 14875
rect 41840 14844 41889 14872
rect 41840 14832 41846 14844
rect 41877 14841 41889 14844
rect 41923 14872 41935 14875
rect 41966 14872 41972 14884
rect 41923 14844 41972 14872
rect 41923 14841 41935 14844
rect 41877 14835 41935 14841
rect 41966 14832 41972 14844
rect 42024 14832 42030 14884
rect 42613 14807 42671 14813
rect 42613 14804 42625 14807
rect 40880 14776 42625 14804
rect 42613 14773 42625 14776
rect 42659 14804 42671 14807
rect 42886 14804 42892 14816
rect 42659 14776 42892 14804
rect 42659 14773 42671 14776
rect 42613 14767 42671 14773
rect 42886 14764 42892 14776
rect 42944 14764 42950 14816
rect 42996 14804 43024 14912
rect 43070 14900 43076 14952
rect 43128 14940 43134 14952
rect 43128 14912 43173 14940
rect 43128 14900 43134 14912
rect 43272 14872 43300 14980
rect 44358 14968 44364 15020
rect 44416 15008 44422 15020
rect 44416 14980 44461 15008
rect 44416 14968 44422 14980
rect 44542 14968 44548 15020
rect 44600 15008 44606 15020
rect 44729 15011 44787 15017
rect 44600 14980 44645 15008
rect 44600 14968 44606 14980
rect 44729 14977 44741 15011
rect 44775 15008 44787 15011
rect 45281 15011 45339 15017
rect 45281 15008 45293 15011
rect 44775 14980 45293 15008
rect 44775 14977 44787 14980
rect 44729 14971 44787 14977
rect 45281 14977 45293 14980
rect 45327 14977 45339 15011
rect 45281 14971 45339 14977
rect 48225 15011 48283 15017
rect 48225 14977 48237 15011
rect 48271 15008 48283 15011
rect 48314 15008 48320 15020
rect 48271 14980 48320 15008
rect 48271 14977 48283 14980
rect 48225 14971 48283 14977
rect 48314 14968 48320 14980
rect 48372 14968 48378 15020
rect 48590 14968 48596 15020
rect 48648 15008 48654 15020
rect 48685 15011 48743 15017
rect 48685 15008 48697 15011
rect 48648 14980 48697 15008
rect 48648 14968 48654 14980
rect 48685 14977 48697 14980
rect 48731 14977 48743 15011
rect 48792 15008 48820 15048
rect 49688 15045 49700 15079
rect 49734 15076 49746 15079
rect 50430 15076 50436 15088
rect 49734 15048 50436 15076
rect 49734 15045 49746 15048
rect 49688 15039 49746 15045
rect 50430 15036 50436 15048
rect 50488 15036 50494 15088
rect 51074 15036 51080 15088
rect 51132 15076 51138 15088
rect 51445 15079 51503 15085
rect 51445 15076 51457 15079
rect 51132 15048 51457 15076
rect 51132 15036 51138 15048
rect 51445 15045 51457 15048
rect 51491 15045 51503 15079
rect 51445 15039 51503 15045
rect 51534 15036 51540 15088
rect 51592 15076 51598 15088
rect 52181 15079 52239 15085
rect 52181 15076 52193 15079
rect 51592 15048 52193 15076
rect 51592 15036 51598 15048
rect 52181 15045 52193 15048
rect 52227 15045 52239 15079
rect 52914 15076 52920 15088
rect 52181 15039 52239 15045
rect 52288 15048 52920 15076
rect 51169 15011 51227 15017
rect 51169 15008 51181 15011
rect 48792 14980 50476 15008
rect 48685 14971 48743 14977
rect 43349 14943 43407 14949
rect 43349 14909 43361 14943
rect 43395 14940 43407 14943
rect 43438 14940 43444 14952
rect 43395 14912 43444 14940
rect 43395 14909 43407 14912
rect 43349 14903 43407 14909
rect 43438 14900 43444 14912
rect 43496 14900 43502 14952
rect 44082 14900 44088 14952
rect 44140 14940 44146 14952
rect 45646 14940 45652 14952
rect 44140 14912 45140 14940
rect 45607 14912 45652 14940
rect 44140 14900 44146 14912
rect 45112 14881 45140 14912
rect 45646 14900 45652 14912
rect 45704 14900 45710 14952
rect 45830 14900 45836 14952
rect 45888 14940 45894 14952
rect 45925 14943 45983 14949
rect 45925 14940 45937 14943
rect 45888 14912 45937 14940
rect 45888 14900 45894 14912
rect 45925 14909 45937 14912
rect 45971 14940 45983 14943
rect 46842 14940 46848 14952
rect 45971 14912 46848 14940
rect 45971 14909 45983 14912
rect 45925 14903 45983 14909
rect 46842 14900 46848 14912
rect 46900 14900 46906 14952
rect 48866 14940 48872 14952
rect 48827 14912 48872 14940
rect 48866 14900 48872 14912
rect 48924 14900 48930 14952
rect 49421 14943 49479 14949
rect 49421 14909 49433 14943
rect 49467 14909 49479 14943
rect 49421 14903 49479 14909
rect 45097 14875 45155 14881
rect 43272 14844 44216 14872
rect 44082 14804 44088 14816
rect 42996 14776 44088 14804
rect 44082 14764 44088 14776
rect 44140 14764 44146 14816
rect 44188 14804 44216 14844
rect 45097 14841 45109 14875
rect 45143 14841 45155 14875
rect 45097 14835 45155 14841
rect 45738 14832 45744 14884
rect 45796 14872 45802 14884
rect 46750 14872 46756 14884
rect 45796 14844 46756 14872
rect 45796 14832 45802 14844
rect 46750 14832 46756 14844
rect 46808 14832 46814 14884
rect 46934 14832 46940 14884
rect 46992 14872 46998 14884
rect 48884 14872 48912 14900
rect 46992 14844 48912 14872
rect 46992 14832 46998 14844
rect 45554 14804 45560 14816
rect 44188 14776 45560 14804
rect 45554 14764 45560 14776
rect 45612 14764 45618 14816
rect 48041 14807 48099 14813
rect 48041 14773 48053 14807
rect 48087 14804 48099 14807
rect 48590 14804 48596 14816
rect 48087 14776 48596 14804
rect 48087 14773 48099 14776
rect 48041 14767 48099 14773
rect 48590 14764 48596 14776
rect 48648 14764 48654 14816
rect 49436 14804 49464 14903
rect 49786 14804 49792 14816
rect 49436 14776 49792 14804
rect 49786 14764 49792 14776
rect 49844 14764 49850 14816
rect 50448 14804 50476 14980
rect 50816 14980 51181 15008
rect 50816 14881 50844 14980
rect 51169 14977 51181 14980
rect 51215 14977 51227 15011
rect 51169 14971 51227 14977
rect 51997 15011 52055 15017
rect 51997 14977 52009 15011
rect 52043 15008 52055 15011
rect 52288 15008 52316 15048
rect 52914 15036 52920 15048
rect 52972 15036 52978 15088
rect 53668 15076 53696 15116
rect 54294 15104 54300 15156
rect 54352 15144 54358 15156
rect 62942 15144 62948 15156
rect 54352 15116 62948 15144
rect 54352 15104 54358 15116
rect 62942 15104 62948 15116
rect 63000 15104 63006 15156
rect 63773 15147 63831 15153
rect 63773 15113 63785 15147
rect 63819 15144 63831 15147
rect 64322 15144 64328 15156
rect 63819 15116 64328 15144
rect 63819 15113 63831 15116
rect 63773 15107 63831 15113
rect 64322 15104 64328 15116
rect 64380 15104 64386 15156
rect 65518 15144 65524 15156
rect 65168 15116 65524 15144
rect 53834 15076 53840 15088
rect 53668 15048 53840 15076
rect 53834 15036 53840 15048
rect 53892 15036 53898 15088
rect 54938 15036 54944 15088
rect 54996 15076 55002 15088
rect 55033 15079 55091 15085
rect 55033 15076 55045 15079
rect 54996 15048 55045 15076
rect 54996 15036 55002 15048
rect 55033 15045 55045 15048
rect 55079 15045 55091 15079
rect 55033 15039 55091 15045
rect 55122 15036 55128 15088
rect 55180 15076 55186 15088
rect 55217 15079 55275 15085
rect 55217 15076 55229 15079
rect 55180 15048 55229 15076
rect 55180 15036 55186 15048
rect 55217 15045 55229 15048
rect 55263 15045 55275 15079
rect 56318 15076 56324 15088
rect 55217 15039 55275 15045
rect 55324 15048 56324 15076
rect 53282 15008 53288 15020
rect 52043 14980 52316 15008
rect 53243 14980 53288 15008
rect 52043 14977 52055 14980
rect 51997 14971 52055 14977
rect 53282 14968 53288 14980
rect 53340 14968 53346 15020
rect 53466 14968 53472 15020
rect 53524 15008 53530 15020
rect 53561 15011 53619 15017
rect 53561 15008 53573 15011
rect 53524 14980 53573 15008
rect 53524 14968 53530 14980
rect 53561 14977 53573 14980
rect 53607 14977 53619 15011
rect 53561 14971 53619 14977
rect 54202 14968 54208 15020
rect 54260 15008 54266 15020
rect 54297 15011 54355 15017
rect 54297 15008 54309 15011
rect 54260 14980 54309 15008
rect 54260 14968 54266 14980
rect 54297 14977 54309 14980
rect 54343 14977 54355 15011
rect 54297 14971 54355 14977
rect 54478 14968 54484 15020
rect 54536 15008 54542 15020
rect 55324 15017 55352 15048
rect 56318 15036 56324 15048
rect 56376 15036 56382 15088
rect 56413 15079 56471 15085
rect 56413 15045 56425 15079
rect 56459 15076 56471 15079
rect 58158 15076 58164 15088
rect 56459 15048 58164 15076
rect 56459 15045 56471 15048
rect 56413 15039 56471 15045
rect 58158 15036 58164 15048
rect 58216 15036 58222 15088
rect 58250 15036 58256 15088
rect 58308 15036 58314 15088
rect 59354 15076 59360 15088
rect 59280 15048 59360 15076
rect 55309 15011 55367 15017
rect 54536 14980 54581 15008
rect 54536 14968 54542 14980
rect 55309 14977 55321 15011
rect 55355 14977 55367 15011
rect 55309 14971 55367 14977
rect 55674 14968 55680 15020
rect 55732 15008 55738 15020
rect 55769 15011 55827 15017
rect 55769 15008 55781 15011
rect 55732 14980 55781 15008
rect 55732 14968 55738 14980
rect 55769 14977 55781 14980
rect 55815 14977 55827 15011
rect 55769 14971 55827 14977
rect 56597 15011 56655 15017
rect 56597 14977 56609 15011
rect 56643 14977 56655 15011
rect 56597 14971 56655 14977
rect 56612 14940 56640 14971
rect 56686 14968 56692 15020
rect 56744 15008 56750 15020
rect 56781 15011 56839 15017
rect 56781 15008 56793 15011
rect 56744 14980 56793 15008
rect 56744 14968 56750 14980
rect 56781 14977 56793 14980
rect 56827 14977 56839 15011
rect 56781 14971 56839 14977
rect 56870 14968 56876 15020
rect 56928 15008 56934 15020
rect 57425 15011 57483 15017
rect 56928 14980 56973 15008
rect 56928 14968 56934 14980
rect 57425 14977 57437 15011
rect 57471 15008 57483 15011
rect 57471 15006 58204 15008
rect 58268 15006 58296 15036
rect 59280 15017 59308 15048
rect 59354 15036 59360 15048
rect 59412 15036 59418 15088
rect 62209 15079 62267 15085
rect 61764 15048 62160 15076
rect 61764 15020 61792 15048
rect 57471 14980 58296 15006
rect 57471 14977 57483 14980
rect 58176 14978 58296 14980
rect 59265 15011 59323 15017
rect 57425 14971 57483 14977
rect 59265 14977 59277 15011
rect 59311 14977 59323 15011
rect 59265 14971 59323 14977
rect 59449 15011 59507 15017
rect 59449 14977 59461 15011
rect 59495 15008 59507 15011
rect 59538 15008 59544 15020
rect 59495 14980 59544 15008
rect 59495 14977 59507 14980
rect 59449 14971 59507 14977
rect 59538 14968 59544 14980
rect 59596 14968 59602 15020
rect 60737 15011 60795 15017
rect 60737 14977 60749 15011
rect 60783 15008 60795 15011
rect 61746 15008 61752 15020
rect 60783 14980 61752 15008
rect 60783 14977 60795 14980
rect 60737 14971 60795 14977
rect 61746 14968 61752 14980
rect 61804 14968 61810 15020
rect 62022 15008 62028 15020
rect 61983 14980 62028 15008
rect 62022 14968 62028 14980
rect 62080 14968 62086 15020
rect 56962 14940 56968 14952
rect 50908 14912 56548 14940
rect 56612 14912 56968 14940
rect 50801 14875 50859 14881
rect 50801 14841 50813 14875
rect 50847 14841 50859 14875
rect 50801 14835 50859 14841
rect 50908 14804 50936 14912
rect 50982 14832 50988 14884
rect 51040 14872 51046 14884
rect 51261 14875 51319 14881
rect 51261 14872 51273 14875
rect 51040 14844 51273 14872
rect 51040 14832 51046 14844
rect 51261 14841 51273 14844
rect 51307 14841 51319 14875
rect 51261 14835 51319 14841
rect 52638 14832 52644 14884
rect 52696 14872 52702 14884
rect 53101 14875 53159 14881
rect 53101 14872 53113 14875
rect 52696 14844 53113 14872
rect 52696 14832 52702 14844
rect 53101 14841 53113 14844
rect 53147 14841 53159 14875
rect 55030 14872 55036 14884
rect 54991 14844 55036 14872
rect 53101 14835 53159 14841
rect 55030 14832 55036 14844
rect 55088 14832 55094 14884
rect 50448 14776 50936 14804
rect 51074 14764 51080 14816
rect 51132 14804 51138 14816
rect 51169 14807 51227 14813
rect 51169 14804 51181 14807
rect 51132 14776 51181 14804
rect 51132 14764 51138 14776
rect 51169 14773 51181 14776
rect 51215 14773 51227 14807
rect 51169 14767 51227 14773
rect 51350 14764 51356 14816
rect 51408 14804 51414 14816
rect 54294 14804 54300 14816
rect 51408 14776 54300 14804
rect 51408 14764 51414 14776
rect 54294 14764 54300 14776
rect 54352 14764 54358 14816
rect 54662 14804 54668 14816
rect 54623 14776 54668 14804
rect 54662 14764 54668 14776
rect 54720 14764 54726 14816
rect 54846 14764 54852 14816
rect 54904 14804 54910 14816
rect 55861 14807 55919 14813
rect 55861 14804 55873 14807
rect 54904 14776 55873 14804
rect 54904 14764 54910 14776
rect 55861 14773 55873 14776
rect 55907 14773 55919 14807
rect 56520 14804 56548 14912
rect 56962 14900 56968 14912
rect 57020 14900 57026 14952
rect 58066 14940 58072 14952
rect 58027 14912 58072 14940
rect 58066 14900 58072 14912
rect 58124 14900 58130 14952
rect 58391 14943 58449 14949
rect 58391 14909 58403 14943
rect 58437 14940 58449 14943
rect 58710 14940 58716 14952
rect 58437 14912 58716 14940
rect 58437 14909 58449 14912
rect 58391 14903 58449 14909
rect 58710 14900 58716 14912
rect 58768 14900 58774 14952
rect 59354 14900 59360 14952
rect 59412 14940 59418 14952
rect 60461 14943 60519 14949
rect 60461 14940 60473 14943
rect 59412 14912 60473 14940
rect 59412 14900 59418 14912
rect 60461 14909 60473 14912
rect 60507 14909 60519 14943
rect 60461 14903 60519 14909
rect 60826 14900 60832 14952
rect 60884 14940 60890 14952
rect 61838 14940 61844 14952
rect 60884 14912 61844 14940
rect 60884 14900 60890 14912
rect 61838 14900 61844 14912
rect 61896 14900 61902 14952
rect 62132 14940 62160 15048
rect 62209 15045 62221 15079
rect 62255 15076 62267 15079
rect 63405 15079 63463 15085
rect 63405 15076 63417 15079
rect 62255 15048 63417 15076
rect 62255 15045 62267 15048
rect 62209 15039 62267 15045
rect 63405 15045 63417 15048
rect 63451 15045 63463 15079
rect 65168 15076 65196 15116
rect 65518 15104 65524 15116
rect 65576 15104 65582 15156
rect 65705 15147 65763 15153
rect 65705 15113 65717 15147
rect 65751 15144 65763 15147
rect 66441 15147 66499 15153
rect 66441 15144 66453 15147
rect 65751 15116 66453 15144
rect 65751 15113 65763 15116
rect 65705 15107 65763 15113
rect 66441 15113 66453 15116
rect 66487 15113 66499 15147
rect 67266 15144 67272 15156
rect 67227 15116 67272 15144
rect 66441 15107 66499 15113
rect 67266 15104 67272 15116
rect 67324 15104 67330 15156
rect 69198 15144 69204 15156
rect 68664 15116 69204 15144
rect 63405 15039 63463 15045
rect 64340 15048 65196 15076
rect 62298 15008 62304 15020
rect 62259 14980 62304 15008
rect 62298 14968 62304 14980
rect 62356 14968 62362 15020
rect 62390 14968 62396 15020
rect 62448 15008 62454 15020
rect 63586 15008 63592 15020
rect 62448 14980 62493 15008
rect 63547 14980 63592 15008
rect 62448 14968 62454 14980
rect 63586 14968 63592 14980
rect 63644 14968 63650 15020
rect 64340 15017 64368 15048
rect 65242 15036 65248 15088
rect 65300 15076 65306 15088
rect 68002 15076 68008 15088
rect 65300 15048 68008 15076
rect 65300 15036 65306 15048
rect 68002 15036 68008 15048
rect 68060 15036 68066 15088
rect 64598 15017 64604 15020
rect 63865 15011 63923 15017
rect 63865 14977 63877 15011
rect 63911 14977 63923 15011
rect 63865 14971 63923 14977
rect 64325 15011 64383 15017
rect 64325 14977 64337 15011
rect 64371 14977 64383 15011
rect 64592 15008 64604 15017
rect 64559 14980 64604 15008
rect 64325 14971 64383 14977
rect 64592 14971 64604 14980
rect 62758 14940 62764 14952
rect 62132 14912 62764 14940
rect 62758 14900 62764 14912
rect 62816 14940 62822 14952
rect 63880 14940 63908 14971
rect 64598 14968 64604 14971
rect 64656 14968 64662 15020
rect 65702 14968 65708 15020
rect 65760 15008 65766 15020
rect 66257 15011 66315 15017
rect 66257 15008 66269 15011
rect 65760 14980 66269 15008
rect 65760 14968 65766 14980
rect 66257 14977 66269 14980
rect 66303 14977 66315 15011
rect 66257 14971 66315 14977
rect 66438 14968 66444 15020
rect 66496 15008 66502 15020
rect 66533 15011 66591 15017
rect 66533 15008 66545 15011
rect 66496 14980 66545 15008
rect 66496 14968 66502 14980
rect 66533 14977 66545 14980
rect 66579 14977 66591 15011
rect 67085 15011 67143 15017
rect 67085 15008 67097 15011
rect 66533 14971 66591 14977
rect 66640 14980 67097 15008
rect 62816 14912 63908 14940
rect 62816 14900 62822 14912
rect 65794 14900 65800 14952
rect 65852 14940 65858 14952
rect 66640 14940 66668 14980
rect 67085 14977 67097 14980
rect 67131 14977 67143 15011
rect 67085 14971 67143 14977
rect 67361 15011 67419 15017
rect 67361 14977 67373 15011
rect 67407 15008 67419 15011
rect 68664 15008 68692 15116
rect 69198 15104 69204 15116
rect 69256 15104 69262 15156
rect 69290 15104 69296 15156
rect 69348 15144 69354 15156
rect 69348 15116 69393 15144
rect 69348 15104 69354 15116
rect 69658 15104 69664 15156
rect 69716 15144 69722 15156
rect 69716 15116 70624 15144
rect 69716 15104 69722 15116
rect 68925 15079 68983 15085
rect 68925 15045 68937 15079
rect 68971 15076 68983 15079
rect 70596 15076 70624 15116
rect 70854 15104 70860 15156
rect 70912 15144 70918 15156
rect 70912 15116 80054 15144
rect 70912 15104 70918 15116
rect 71958 15076 71964 15088
rect 68971 15048 69428 15076
rect 70596 15048 71964 15076
rect 68971 15045 68983 15048
rect 68925 15039 68983 15045
rect 67407 14980 68692 15008
rect 67407 14977 67419 14980
rect 67361 14971 67419 14977
rect 68738 14968 68744 15020
rect 68796 15008 68802 15020
rect 69013 15011 69071 15017
rect 69013 15008 69025 15011
rect 68796 14980 68841 15008
rect 68934 14980 69025 15008
rect 68796 14968 68802 14980
rect 65852 14912 66668 14940
rect 66901 14943 66959 14949
rect 65852 14900 65858 14912
rect 66901 14909 66913 14943
rect 66947 14940 66959 14943
rect 68646 14940 68652 14952
rect 66947 14912 68652 14940
rect 66947 14909 66959 14912
rect 66901 14903 66959 14909
rect 68646 14900 68652 14912
rect 68704 14900 68710 14952
rect 68934 14940 68962 14980
rect 69013 14977 69025 14980
rect 69059 14977 69071 15011
rect 69013 14971 69071 14977
rect 69109 15011 69167 15017
rect 69109 14977 69121 15011
rect 69155 15008 69167 15011
rect 69198 15008 69204 15020
rect 69155 14980 69204 15008
rect 69155 14977 69167 14980
rect 69109 14971 69167 14977
rect 69198 14968 69204 14980
rect 69256 14968 69262 15020
rect 69400 15008 69428 15048
rect 71958 15036 71964 15048
rect 72016 15036 72022 15088
rect 80026 15076 80054 15116
rect 88242 15076 88248 15088
rect 80026 15048 88248 15076
rect 88242 15036 88248 15048
rect 88300 15036 88306 15088
rect 69474 15008 69480 15020
rect 69400 14980 69480 15008
rect 69474 14968 69480 14980
rect 69532 14968 69538 15020
rect 69661 15011 69719 15017
rect 69661 15008 69673 15011
rect 69584 14980 69673 15008
rect 69584 14940 69612 14980
rect 69661 14977 69673 14980
rect 69707 15008 69719 15011
rect 69750 15008 69756 15020
rect 69707 14980 69756 15008
rect 69707 14977 69719 14980
rect 69661 14971 69719 14977
rect 69750 14968 69756 14980
rect 69808 14968 69814 15020
rect 69937 15011 69995 15017
rect 69937 14977 69949 15011
rect 69983 15008 69995 15011
rect 71685 15011 71743 15017
rect 71685 15008 71697 15011
rect 69983 14980 71697 15008
rect 69983 14977 69995 14980
rect 69937 14971 69995 14977
rect 71685 14977 71697 14980
rect 71731 15008 71743 15011
rect 88150 15008 88156 15020
rect 71731 14980 88156 15008
rect 71731 14977 71743 14980
rect 71685 14971 71743 14977
rect 69952 14940 69980 14971
rect 88150 14968 88156 14980
rect 88208 14968 88214 15020
rect 68776 14912 68962 14940
rect 69032 14912 69612 14940
rect 69656 14912 69980 14940
rect 57241 14875 57299 14881
rect 57241 14841 57253 14875
rect 57287 14872 57299 14875
rect 57974 14872 57980 14884
rect 57287 14844 57980 14872
rect 57287 14841 57299 14844
rect 57241 14835 57299 14841
rect 57974 14832 57980 14844
rect 58032 14832 58038 14884
rect 63954 14872 63960 14884
rect 58084 14844 63960 14872
rect 58084 14804 58112 14844
rect 63954 14832 63960 14844
rect 64012 14832 64018 14884
rect 65334 14832 65340 14884
rect 65392 14872 65398 14884
rect 68776 14872 68804 14912
rect 65392 14844 68804 14872
rect 65392 14832 65398 14844
rect 68922 14832 68928 14884
rect 68980 14872 68986 14884
rect 69032 14872 69060 14912
rect 69656 14872 69684 14912
rect 70670 14900 70676 14952
rect 70728 14940 70734 14952
rect 71041 14943 71099 14949
rect 71041 14940 71053 14943
rect 70728 14912 71053 14940
rect 70728 14900 70734 14912
rect 71041 14909 71053 14912
rect 71087 14909 71099 14943
rect 71041 14903 71099 14909
rect 74810 14872 74816 14884
rect 68980 14844 69060 14872
rect 69124 14844 69684 14872
rect 70964 14844 74816 14872
rect 68980 14832 68986 14844
rect 56520 14776 58112 14804
rect 55861 14767 55919 14773
rect 58342 14764 58348 14816
rect 58400 14804 58406 14816
rect 59633 14807 59691 14813
rect 59633 14804 59645 14807
rect 58400 14776 59645 14804
rect 58400 14764 58406 14776
rect 59633 14773 59645 14776
rect 59679 14773 59691 14807
rect 59633 14767 59691 14773
rect 62577 14807 62635 14813
rect 62577 14773 62589 14807
rect 62623 14804 62635 14807
rect 63218 14804 63224 14816
rect 62623 14776 63224 14804
rect 62623 14773 62635 14776
rect 62577 14767 62635 14773
rect 63218 14764 63224 14776
rect 63276 14764 63282 14816
rect 63586 14764 63592 14816
rect 63644 14804 63650 14816
rect 63862 14804 63868 14816
rect 63644 14776 63868 14804
rect 63644 14764 63650 14776
rect 63862 14764 63868 14776
rect 63920 14764 63926 14816
rect 64598 14764 64604 14816
rect 64656 14804 64662 14816
rect 66073 14807 66131 14813
rect 66073 14804 66085 14807
rect 64656 14776 66085 14804
rect 64656 14764 64662 14776
rect 66073 14773 66085 14776
rect 66119 14773 66131 14807
rect 66073 14767 66131 14773
rect 68738 14764 68744 14816
rect 68796 14804 68802 14816
rect 69124 14804 69152 14844
rect 68796 14776 69152 14804
rect 68796 14764 68802 14776
rect 69198 14764 69204 14816
rect 69256 14804 69262 14816
rect 70964 14804 70992 14844
rect 74810 14832 74816 14844
rect 74868 14832 74874 14884
rect 69256 14776 70992 14804
rect 69256 14764 69262 14776
rect 71222 14764 71228 14816
rect 71280 14804 71286 14816
rect 71869 14807 71927 14813
rect 71869 14804 71881 14807
rect 71280 14776 71881 14804
rect 71280 14764 71286 14776
rect 71869 14773 71881 14776
rect 71915 14804 71927 14807
rect 72050 14804 72056 14816
rect 71915 14776 72056 14804
rect 71915 14773 71927 14776
rect 71869 14767 71927 14773
rect 72050 14764 72056 14776
rect 72108 14764 72114 14816
rect 1104 14714 88872 14736
rect 1104 14662 11924 14714
rect 11976 14662 11988 14714
rect 12040 14662 12052 14714
rect 12104 14662 12116 14714
rect 12168 14662 12180 14714
rect 12232 14662 33872 14714
rect 33924 14662 33936 14714
rect 33988 14662 34000 14714
rect 34052 14662 34064 14714
rect 34116 14662 34128 14714
rect 34180 14662 55820 14714
rect 55872 14662 55884 14714
rect 55936 14662 55948 14714
rect 56000 14662 56012 14714
rect 56064 14662 56076 14714
rect 56128 14662 77768 14714
rect 77820 14662 77832 14714
rect 77884 14662 77896 14714
rect 77948 14662 77960 14714
rect 78012 14662 78024 14714
rect 78076 14662 88872 14714
rect 1104 14640 88872 14662
rect 21174 14560 21180 14612
rect 21232 14600 21238 14612
rect 21634 14600 21640 14612
rect 21232 14572 21640 14600
rect 21232 14560 21238 14572
rect 21634 14560 21640 14572
rect 21692 14600 21698 14612
rect 22738 14600 22744 14612
rect 21692 14572 22744 14600
rect 21692 14560 21698 14572
rect 22738 14560 22744 14572
rect 22796 14560 22802 14612
rect 23201 14603 23259 14609
rect 23201 14569 23213 14603
rect 23247 14569 23259 14603
rect 23201 14563 23259 14569
rect 6638 14492 6644 14544
rect 6696 14532 6702 14544
rect 6696 14504 21680 14532
rect 6696 14492 6702 14504
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 21652 14405 21680 14504
rect 22186 14492 22192 14544
rect 22244 14532 22250 14544
rect 22554 14532 22560 14544
rect 22244 14504 22560 14532
rect 22244 14492 22250 14504
rect 22554 14492 22560 14504
rect 22612 14492 22618 14544
rect 23216 14532 23244 14563
rect 23290 14560 23296 14612
rect 23348 14600 23354 14612
rect 26050 14600 26056 14612
rect 23348 14572 26056 14600
rect 23348 14560 23354 14572
rect 26050 14560 26056 14572
rect 26108 14560 26114 14612
rect 26145 14603 26203 14609
rect 26145 14569 26157 14603
rect 26191 14600 26203 14603
rect 26878 14600 26884 14612
rect 26191 14572 26884 14600
rect 26191 14569 26203 14572
rect 26145 14563 26203 14569
rect 26878 14560 26884 14572
rect 26936 14560 26942 14612
rect 27062 14560 27068 14612
rect 27120 14600 27126 14612
rect 28810 14600 28816 14612
rect 27120 14572 28816 14600
rect 27120 14560 27126 14572
rect 28810 14560 28816 14572
rect 28868 14560 28874 14612
rect 31294 14560 31300 14612
rect 31352 14600 31358 14612
rect 31846 14600 31852 14612
rect 31352 14572 31852 14600
rect 31352 14560 31358 14572
rect 31846 14560 31852 14572
rect 31904 14560 31910 14612
rect 31938 14560 31944 14612
rect 31996 14600 32002 14612
rect 37090 14600 37096 14612
rect 31996 14572 36952 14600
rect 37051 14572 37096 14600
rect 31996 14560 32002 14572
rect 24762 14532 24768 14544
rect 23216 14504 24768 14532
rect 24762 14492 24768 14504
rect 24820 14532 24826 14544
rect 24946 14532 24952 14544
rect 24820 14504 24952 14532
rect 24820 14492 24826 14504
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 26602 14532 26608 14544
rect 26252 14504 26608 14532
rect 21726 14424 21732 14476
rect 21784 14464 21790 14476
rect 22649 14467 22707 14473
rect 22649 14464 22661 14467
rect 21784 14436 22661 14464
rect 21784 14424 21790 14436
rect 22649 14433 22661 14436
rect 22695 14433 22707 14467
rect 26252 14464 26280 14504
rect 26602 14492 26608 14504
rect 26660 14492 26666 14544
rect 28077 14535 28135 14541
rect 28077 14532 28089 14535
rect 27724 14504 28089 14532
rect 22649 14427 22707 14433
rect 23124 14436 26280 14464
rect 20533 14399 20591 14405
rect 20533 14396 20545 14399
rect 20404 14368 20545 14396
rect 20404 14356 20410 14368
rect 20533 14365 20545 14368
rect 20579 14365 20591 14399
rect 20533 14359 20591 14365
rect 20625 14399 20683 14405
rect 20625 14365 20637 14399
rect 20671 14396 20683 14399
rect 21269 14399 21327 14405
rect 21269 14396 21281 14399
rect 20671 14368 21281 14396
rect 20671 14365 20683 14368
rect 20625 14359 20683 14365
rect 21269 14365 21281 14368
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 21361 14399 21419 14405
rect 21361 14365 21373 14399
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 21545 14399 21603 14405
rect 21545 14365 21557 14399
rect 21591 14365 21603 14399
rect 21545 14359 21603 14365
rect 21637 14399 21695 14405
rect 21637 14365 21649 14399
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 20898 14288 20904 14340
rect 20956 14328 20962 14340
rect 21376 14328 21404 14359
rect 20956 14300 21404 14328
rect 21560 14328 21588 14359
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 22189 14399 22247 14405
rect 22189 14396 22201 14399
rect 22152 14368 22201 14396
rect 22152 14356 22158 14368
rect 22189 14365 22201 14368
rect 22235 14365 22247 14399
rect 22189 14359 22247 14365
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 23124 14405 23152 14436
rect 23109 14399 23167 14405
rect 22336 14368 22381 14396
rect 22480 14368 23060 14396
rect 22336 14356 22342 14368
rect 22480 14328 22508 14368
rect 21560 14300 22508 14328
rect 20956 14288 20962 14300
rect 22554 14288 22560 14340
rect 22612 14328 22618 14340
rect 23032 14328 23060 14368
rect 23109 14365 23121 14399
rect 23155 14365 23167 14399
rect 24394 14396 24400 14408
rect 24355 14368 24400 14396
rect 23109 14359 23167 14365
rect 24394 14356 24400 14368
rect 24452 14356 24458 14408
rect 24762 14396 24768 14408
rect 24723 14368 24768 14396
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 25590 14396 25596 14408
rect 24872 14368 25596 14396
rect 23934 14328 23940 14340
rect 22612 14300 22657 14328
rect 23032 14300 23940 14328
rect 22612 14288 22618 14300
rect 23934 14288 23940 14300
rect 23992 14288 23998 14340
rect 24581 14331 24639 14337
rect 24581 14297 24593 14331
rect 24627 14297 24639 14331
rect 24581 14291 24639 14297
rect 1397 14263 1455 14269
rect 1397 14229 1409 14263
rect 1443 14260 1455 14263
rect 18230 14260 18236 14272
rect 1443 14232 18236 14260
rect 1443 14229 1455 14232
rect 1397 14223 1455 14229
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 20254 14220 20260 14272
rect 20312 14260 20318 14272
rect 20622 14260 20628 14272
rect 20312 14232 20628 14260
rect 20312 14220 20318 14232
rect 20622 14220 20628 14232
rect 20680 14220 20686 14272
rect 21085 14263 21143 14269
rect 21085 14229 21097 14263
rect 21131 14260 21143 14263
rect 21542 14260 21548 14272
rect 21131 14232 21548 14260
rect 21131 14229 21143 14232
rect 21085 14223 21143 14229
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 22005 14263 22063 14269
rect 22005 14229 22017 14263
rect 22051 14260 22063 14263
rect 22462 14260 22468 14272
rect 22051 14232 22468 14260
rect 22051 14229 22063 14232
rect 22005 14223 22063 14229
rect 22462 14220 22468 14232
rect 22520 14220 22526 14272
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 23569 14263 23627 14269
rect 23569 14260 23581 14263
rect 22796 14232 23581 14260
rect 22796 14220 22802 14232
rect 23569 14229 23581 14232
rect 23615 14229 23627 14263
rect 24596 14260 24624 14291
rect 24670 14288 24676 14340
rect 24728 14328 24734 14340
rect 24872 14328 24900 14368
rect 25590 14356 25596 14368
rect 25648 14356 25654 14408
rect 25774 14396 25780 14408
rect 25735 14368 25780 14396
rect 25774 14356 25780 14368
rect 25832 14356 25838 14408
rect 26329 14399 26387 14405
rect 26329 14365 26341 14399
rect 26375 14395 26387 14399
rect 26510 14396 26516 14408
rect 26436 14395 26516 14396
rect 26375 14368 26516 14395
rect 26375 14367 26464 14368
rect 26375 14365 26387 14367
rect 26329 14359 26387 14365
rect 26510 14356 26516 14368
rect 26568 14356 26574 14408
rect 26694 14396 26700 14408
rect 26655 14368 26700 14396
rect 26694 14356 26700 14368
rect 26752 14356 26758 14408
rect 27246 14356 27252 14408
rect 27304 14396 27310 14408
rect 27724 14396 27752 14504
rect 28077 14501 28089 14504
rect 28123 14501 28135 14535
rect 31478 14532 31484 14544
rect 28077 14495 28135 14501
rect 28736 14504 31484 14532
rect 27890 14424 27896 14476
rect 27948 14464 27954 14476
rect 28736 14464 28764 14504
rect 31478 14492 31484 14504
rect 31536 14492 31542 14544
rect 33689 14535 33747 14541
rect 33689 14501 33701 14535
rect 33735 14532 33747 14535
rect 34514 14532 34520 14544
rect 33735 14504 34520 14532
rect 33735 14501 33747 14504
rect 33689 14495 33747 14501
rect 34514 14492 34520 14504
rect 34572 14492 34578 14544
rect 35066 14492 35072 14544
rect 35124 14532 35130 14544
rect 35805 14535 35863 14541
rect 35805 14532 35817 14535
rect 35124 14504 35817 14532
rect 35124 14492 35130 14504
rect 35805 14501 35817 14504
rect 35851 14501 35863 14535
rect 36924 14532 36952 14572
rect 37090 14560 37096 14572
rect 37148 14560 37154 14612
rect 37737 14603 37795 14609
rect 37737 14569 37749 14603
rect 37783 14600 37795 14603
rect 37826 14600 37832 14612
rect 37783 14572 37832 14600
rect 37783 14569 37795 14572
rect 37737 14563 37795 14569
rect 37826 14560 37832 14572
rect 37884 14560 37890 14612
rect 45002 14600 45008 14612
rect 38626 14572 45008 14600
rect 38626 14532 38654 14572
rect 45002 14560 45008 14572
rect 45060 14560 45066 14612
rect 45186 14560 45192 14612
rect 45244 14600 45250 14612
rect 50890 14600 50896 14612
rect 45244 14572 50896 14600
rect 45244 14560 45250 14572
rect 50890 14560 50896 14572
rect 50948 14560 50954 14612
rect 51626 14560 51632 14612
rect 51684 14600 51690 14612
rect 52181 14603 52239 14609
rect 52181 14600 52193 14603
rect 51684 14572 52193 14600
rect 51684 14560 51690 14572
rect 52181 14569 52193 14572
rect 52227 14600 52239 14603
rect 53282 14600 53288 14612
rect 52227 14572 53288 14600
rect 52227 14569 52239 14572
rect 52181 14563 52239 14569
rect 53282 14560 53288 14572
rect 53340 14600 53346 14612
rect 54386 14600 54392 14612
rect 53340 14572 54392 14600
rect 53340 14560 53346 14572
rect 54386 14560 54392 14572
rect 54444 14560 54450 14612
rect 56060 14572 80054 14600
rect 36924 14504 38654 14532
rect 39209 14535 39267 14541
rect 35805 14495 35863 14501
rect 39209 14501 39221 14535
rect 39255 14501 39267 14535
rect 39209 14495 39267 14501
rect 27948 14436 28764 14464
rect 27948 14424 27954 14436
rect 28736 14405 28764 14436
rect 30466 14424 30472 14476
rect 30524 14464 30530 14476
rect 30837 14467 30895 14473
rect 30837 14464 30849 14467
rect 30524 14436 30849 14464
rect 30524 14424 30530 14436
rect 30837 14433 30849 14436
rect 30883 14464 30895 14467
rect 31662 14464 31668 14476
rect 30883 14436 31668 14464
rect 30883 14433 30895 14436
rect 30837 14427 30895 14433
rect 31662 14424 31668 14436
rect 31720 14424 31726 14476
rect 32030 14464 32036 14476
rect 31991 14436 32036 14464
rect 32030 14424 32036 14436
rect 32088 14424 32094 14476
rect 35618 14464 35624 14476
rect 33612 14436 35624 14464
rect 27304 14368 27752 14396
rect 28721 14399 28779 14405
rect 27304 14356 27310 14368
rect 28721 14365 28733 14399
rect 28767 14365 28779 14399
rect 28902 14396 28908 14408
rect 28863 14368 28908 14396
rect 28721 14359 28779 14365
rect 28902 14356 28908 14368
rect 28960 14356 28966 14408
rect 28997 14399 29055 14405
rect 28997 14365 29009 14399
rect 29043 14396 29055 14399
rect 29270 14396 29276 14408
rect 29043 14368 29276 14396
rect 29043 14365 29055 14368
rect 28997 14359 29055 14365
rect 29270 14356 29276 14368
rect 29328 14396 29334 14408
rect 29638 14396 29644 14408
rect 29328 14368 29644 14396
rect 29328 14356 29334 14368
rect 29638 14356 29644 14368
rect 29696 14356 29702 14408
rect 30009 14399 30067 14405
rect 30009 14365 30021 14399
rect 30055 14396 30067 14399
rect 30190 14396 30196 14408
rect 30055 14368 30196 14396
rect 30055 14365 30067 14368
rect 30009 14359 30067 14365
rect 30190 14356 30196 14368
rect 30248 14396 30254 14408
rect 30653 14399 30711 14405
rect 30653 14396 30665 14399
rect 30248 14368 30665 14396
rect 30248 14356 30254 14368
rect 30653 14365 30665 14368
rect 30699 14396 30711 14399
rect 31110 14396 31116 14408
rect 30699 14368 31116 14396
rect 30699 14365 30711 14368
rect 30653 14359 30711 14365
rect 31110 14356 31116 14368
rect 31168 14396 31174 14408
rect 31297 14399 31355 14405
rect 31297 14396 31309 14399
rect 31168 14368 31309 14396
rect 31168 14356 31174 14368
rect 31297 14365 31309 14368
rect 31343 14396 31355 14399
rect 31846 14396 31852 14408
rect 31343 14368 31852 14396
rect 31343 14365 31355 14368
rect 31297 14359 31355 14365
rect 31846 14356 31852 14368
rect 31904 14356 31910 14408
rect 32766 14356 32772 14408
rect 32824 14396 32830 14408
rect 33612 14396 33640 14436
rect 35618 14424 35624 14436
rect 35676 14424 35682 14476
rect 36541 14467 36599 14473
rect 36541 14464 36553 14467
rect 36096 14436 36553 14464
rect 32824 14368 33640 14396
rect 33689 14399 33747 14405
rect 32824 14356 32830 14368
rect 33689 14365 33701 14399
rect 33735 14396 33747 14399
rect 33870 14396 33876 14408
rect 33735 14368 33876 14396
rect 33735 14365 33747 14368
rect 33689 14359 33747 14365
rect 33870 14356 33876 14368
rect 33928 14356 33934 14408
rect 33965 14399 34023 14405
rect 33965 14365 33977 14399
rect 34011 14396 34023 14399
rect 34698 14396 34704 14408
rect 34011 14368 34704 14396
rect 34011 14365 34023 14368
rect 33965 14359 34023 14365
rect 34698 14356 34704 14368
rect 34756 14356 34762 14408
rect 34974 14396 34980 14408
rect 34935 14368 34980 14396
rect 34974 14356 34980 14368
rect 35032 14356 35038 14408
rect 36096 14405 36124 14436
rect 36541 14433 36553 14436
rect 36587 14433 36599 14467
rect 38562 14464 38568 14476
rect 36541 14427 36599 14433
rect 37200 14436 38568 14464
rect 35161 14399 35219 14405
rect 35161 14365 35173 14399
rect 35207 14396 35219 14399
rect 35713 14399 35771 14405
rect 35713 14396 35725 14399
rect 35207 14368 35725 14396
rect 35207 14365 35219 14368
rect 35161 14359 35219 14365
rect 35713 14365 35725 14368
rect 35759 14396 35771 14399
rect 36081 14399 36139 14405
rect 35759 14368 36032 14396
rect 35759 14365 35771 14368
rect 35713 14359 35771 14365
rect 26942 14331 27000 14337
rect 26942 14328 26954 14331
rect 24728 14300 24900 14328
rect 25608 14300 26954 14328
rect 24728 14288 24734 14300
rect 24854 14260 24860 14272
rect 24596 14232 24860 14260
rect 23569 14223 23627 14229
rect 24854 14220 24860 14232
rect 24912 14220 24918 14272
rect 24949 14263 25007 14269
rect 24949 14229 24961 14263
rect 24995 14260 25007 14263
rect 25222 14260 25228 14272
rect 24995 14232 25228 14260
rect 24995 14229 25007 14232
rect 24949 14223 25007 14229
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 25608 14269 25636 14300
rect 26942 14297 26954 14300
rect 26988 14297 27000 14331
rect 26942 14291 27000 14297
rect 27062 14288 27068 14340
rect 27120 14328 27126 14340
rect 27522 14328 27528 14340
rect 27120 14300 27528 14328
rect 27120 14288 27126 14300
rect 27522 14288 27528 14300
rect 27580 14288 27586 14340
rect 27706 14288 27712 14340
rect 27764 14328 27770 14340
rect 28537 14331 28595 14337
rect 28537 14328 28549 14331
rect 27764 14300 28549 14328
rect 27764 14288 27770 14300
rect 28537 14297 28549 14300
rect 28583 14297 28595 14331
rect 28537 14291 28595 14297
rect 28810 14288 28816 14340
rect 28868 14328 28874 14340
rect 30742 14328 30748 14340
rect 28868 14300 30748 14328
rect 28868 14288 28874 14300
rect 30742 14288 30748 14300
rect 30800 14288 30806 14340
rect 31570 14288 31576 14340
rect 31628 14328 31634 14340
rect 32278 14331 32336 14337
rect 32278 14328 32290 14331
rect 31628 14300 32290 14328
rect 31628 14288 31634 14300
rect 32278 14297 32290 14300
rect 32324 14297 32336 14331
rect 34238 14328 34244 14340
rect 32278 14291 32336 14297
rect 33428 14300 34244 14328
rect 25593 14263 25651 14269
rect 25593 14229 25605 14263
rect 25639 14229 25651 14263
rect 25593 14223 25651 14229
rect 26050 14220 26056 14272
rect 26108 14260 26114 14272
rect 27890 14260 27896 14272
rect 26108 14232 27896 14260
rect 26108 14220 26114 14232
rect 27890 14220 27896 14232
rect 27948 14220 27954 14272
rect 30006 14220 30012 14272
rect 30064 14260 30070 14272
rect 30101 14263 30159 14269
rect 30101 14260 30113 14263
rect 30064 14232 30113 14260
rect 30064 14220 30070 14232
rect 30101 14229 30113 14232
rect 30147 14229 30159 14263
rect 30101 14223 30159 14229
rect 31202 14220 31208 14272
rect 31260 14260 31266 14272
rect 33428 14269 33456 14300
rect 34238 14288 34244 14300
rect 34296 14288 34302 14340
rect 34333 14331 34391 14337
rect 34333 14297 34345 14331
rect 34379 14328 34391 14331
rect 34882 14328 34888 14340
rect 34379 14300 34888 14328
rect 34379 14297 34391 14300
rect 34333 14291 34391 14297
rect 34882 14288 34888 14300
rect 34940 14328 34946 14340
rect 35176 14328 35204 14359
rect 34940 14300 35204 14328
rect 34940 14288 34946 14300
rect 35434 14288 35440 14340
rect 35492 14328 35498 14340
rect 35492 14300 35664 14328
rect 35492 14288 35498 14300
rect 31389 14263 31447 14269
rect 31389 14260 31401 14263
rect 31260 14232 31401 14260
rect 31260 14220 31266 14232
rect 31389 14229 31401 14232
rect 31435 14229 31447 14263
rect 31389 14223 31447 14229
rect 33413 14263 33471 14269
rect 33413 14229 33425 14263
rect 33459 14229 33471 14263
rect 33413 14223 33471 14229
rect 33873 14263 33931 14269
rect 33873 14229 33885 14263
rect 33919 14260 33931 14263
rect 34146 14260 34152 14272
rect 33919 14232 34152 14260
rect 33919 14229 33931 14232
rect 33873 14223 33931 14229
rect 34146 14220 34152 14232
rect 34204 14220 34210 14272
rect 34422 14220 34428 14272
rect 34480 14260 34486 14272
rect 35345 14263 35403 14269
rect 35345 14260 35357 14263
rect 34480 14232 35357 14260
rect 34480 14220 34486 14232
rect 35345 14229 35357 14232
rect 35391 14229 35403 14263
rect 35636 14260 35664 14300
rect 35802 14288 35808 14340
rect 35860 14328 35866 14340
rect 36004 14328 36032 14368
rect 36081 14365 36093 14399
rect 36127 14365 36139 14399
rect 36081 14359 36139 14365
rect 36449 14399 36507 14405
rect 36449 14365 36461 14399
rect 36495 14396 36507 14399
rect 37200 14396 37228 14436
rect 38562 14424 38568 14436
rect 38620 14424 38626 14476
rect 39224 14464 39252 14495
rect 39390 14492 39396 14544
rect 39448 14532 39454 14544
rect 41233 14535 41291 14541
rect 39448 14504 39896 14532
rect 39448 14492 39454 14504
rect 39224 14436 39712 14464
rect 36495 14368 37228 14396
rect 37277 14399 37335 14405
rect 36495 14365 36507 14368
rect 36449 14359 36507 14365
rect 37277 14365 37289 14399
rect 37323 14396 37335 14399
rect 37550 14396 37556 14408
rect 37323 14368 37556 14396
rect 37323 14365 37335 14368
rect 37277 14359 37335 14365
rect 37550 14356 37556 14368
rect 37608 14356 37614 14408
rect 37918 14396 37924 14408
rect 37879 14368 37924 14396
rect 37918 14356 37924 14368
rect 37976 14356 37982 14408
rect 38286 14396 38292 14408
rect 38247 14368 38292 14396
rect 38286 14356 38292 14368
rect 38344 14356 38350 14408
rect 38470 14396 38476 14408
rect 38431 14368 38476 14396
rect 38470 14356 38476 14368
rect 38528 14356 38534 14408
rect 39390 14396 39396 14408
rect 39351 14368 39396 14396
rect 39390 14356 39396 14368
rect 39448 14356 39454 14408
rect 39684 14396 39712 14436
rect 39758 14424 39764 14476
rect 39816 14464 39822 14476
rect 39868 14473 39896 14504
rect 41233 14501 41245 14535
rect 41279 14532 41291 14535
rect 41322 14532 41328 14544
rect 41279 14504 41328 14532
rect 41279 14501 41291 14504
rect 41233 14495 41291 14501
rect 41322 14492 41328 14504
rect 41380 14492 41386 14544
rect 42794 14532 42800 14544
rect 42076 14504 42800 14532
rect 39853 14467 39911 14473
rect 39853 14464 39865 14467
rect 39816 14436 39865 14464
rect 39816 14424 39822 14436
rect 39853 14433 39865 14436
rect 39899 14433 39911 14467
rect 39853 14427 39911 14433
rect 41601 14467 41659 14473
rect 41601 14433 41613 14467
rect 41647 14464 41659 14467
rect 42076 14464 42104 14504
rect 42794 14492 42800 14504
rect 42852 14492 42858 14544
rect 44174 14532 44180 14544
rect 44135 14504 44180 14532
rect 44174 14492 44180 14504
rect 44232 14492 44238 14544
rect 45278 14492 45284 14544
rect 45336 14492 45342 14544
rect 45554 14532 45560 14544
rect 45515 14504 45560 14532
rect 45554 14492 45560 14504
rect 45612 14492 45618 14544
rect 46201 14535 46259 14541
rect 46201 14501 46213 14535
rect 46247 14532 46259 14535
rect 46247 14504 50660 14532
rect 46247 14501 46259 14504
rect 46201 14495 46259 14501
rect 41647 14436 42104 14464
rect 41647 14433 41659 14436
rect 41601 14427 41659 14433
rect 42150 14424 42156 14476
rect 42208 14464 42214 14476
rect 43257 14467 43315 14473
rect 43257 14464 43269 14467
rect 42208 14436 43269 14464
rect 42208 14424 42214 14436
rect 43257 14433 43269 14436
rect 43303 14433 43315 14467
rect 43257 14427 43315 14433
rect 43441 14467 43499 14473
rect 43441 14433 43453 14467
rect 43487 14464 43499 14467
rect 43530 14464 43536 14476
rect 43487 14436 43536 14464
rect 43487 14433 43499 14436
rect 43441 14427 43499 14433
rect 43530 14424 43536 14436
rect 43588 14424 43594 14476
rect 44818 14464 44824 14476
rect 43640 14436 44824 14464
rect 40109 14399 40167 14405
rect 40109 14396 40121 14399
rect 39684 14368 40121 14396
rect 40109 14365 40121 14368
rect 40155 14365 40167 14399
rect 40109 14359 40167 14365
rect 40586 14356 40592 14408
rect 40644 14396 40650 14408
rect 41874 14396 41880 14408
rect 40644 14368 41880 14396
rect 40644 14356 40650 14368
rect 41874 14356 41880 14368
rect 41932 14356 41938 14408
rect 43640 14396 43668 14436
rect 44818 14424 44824 14436
rect 44876 14424 44882 14476
rect 45097 14467 45155 14473
rect 45097 14464 45109 14467
rect 44928 14436 45109 14464
rect 43898 14396 43904 14408
rect 43088 14368 43668 14396
rect 43859 14368 43904 14396
rect 36170 14328 36176 14340
rect 35860 14300 35905 14328
rect 36004 14300 36176 14328
rect 35860 14288 35866 14300
rect 36170 14288 36176 14300
rect 36228 14328 36234 14340
rect 39942 14328 39948 14340
rect 36228 14300 39948 14328
rect 36228 14288 36234 14300
rect 39942 14288 39948 14300
rect 40000 14288 40006 14340
rect 40218 14288 40224 14340
rect 40276 14328 40282 14340
rect 43088 14328 43116 14368
rect 43898 14356 43904 14368
rect 43956 14356 43962 14408
rect 43990 14356 43996 14408
rect 44048 14396 44054 14408
rect 44177 14399 44235 14405
rect 44177 14396 44189 14399
rect 44048 14368 44189 14396
rect 44048 14356 44054 14368
rect 44177 14365 44189 14368
rect 44223 14365 44235 14399
rect 44177 14359 44235 14365
rect 44542 14356 44548 14408
rect 44600 14396 44606 14408
rect 44928 14396 44956 14436
rect 45097 14433 45109 14436
rect 45143 14433 45155 14467
rect 45296 14464 45324 14492
rect 48869 14467 48927 14473
rect 45296 14436 46244 14464
rect 45097 14427 45155 14433
rect 44600 14368 44956 14396
rect 45005 14399 45063 14405
rect 44600 14356 44606 14368
rect 45005 14365 45017 14399
rect 45051 14398 45063 14399
rect 45051 14396 45140 14398
rect 45278 14396 45284 14408
rect 45051 14370 45284 14396
rect 45051 14365 45063 14370
rect 45112 14368 45284 14370
rect 45005 14359 45063 14365
rect 45278 14356 45284 14368
rect 45336 14396 45342 14408
rect 45741 14399 45799 14405
rect 45741 14396 45753 14399
rect 45336 14368 45753 14396
rect 45336 14356 45342 14368
rect 45741 14365 45753 14368
rect 45787 14365 45799 14399
rect 45741 14359 45799 14365
rect 46109 14399 46167 14405
rect 46109 14365 46121 14399
rect 46155 14365 46167 14399
rect 46109 14359 46167 14365
rect 40276 14300 43116 14328
rect 43165 14331 43223 14337
rect 40276 14288 40282 14300
rect 43165 14297 43177 14331
rect 43211 14328 43223 14331
rect 43622 14328 43628 14340
rect 43211 14300 43628 14328
rect 43211 14297 43223 14300
rect 43165 14291 43223 14297
rect 43622 14288 43628 14300
rect 43680 14328 43686 14340
rect 46124 14328 46152 14359
rect 43680 14300 46152 14328
rect 46216 14328 46244 14436
rect 47596 14436 47900 14464
rect 47596 14405 47624 14436
rect 47581 14399 47639 14405
rect 47581 14365 47593 14399
rect 47627 14365 47639 14399
rect 47762 14396 47768 14408
rect 47723 14368 47768 14396
rect 47581 14359 47639 14365
rect 47762 14356 47768 14368
rect 47820 14356 47826 14408
rect 47872 14396 47900 14436
rect 48869 14433 48881 14467
rect 48915 14464 48927 14467
rect 50632 14464 50660 14504
rect 50982 14492 50988 14544
rect 51040 14532 51046 14544
rect 56060 14532 56088 14572
rect 51040 14504 52132 14532
rect 51040 14492 51046 14504
rect 51994 14464 52000 14476
rect 48915 14436 50568 14464
rect 50632 14436 52000 14464
rect 48915 14433 48927 14436
rect 48869 14427 48927 14433
rect 48319 14399 48377 14405
rect 48319 14396 48331 14399
rect 47872 14368 48331 14396
rect 48319 14365 48331 14368
rect 48365 14396 48377 14399
rect 48590 14396 48596 14408
rect 48365 14368 48596 14396
rect 48365 14365 48377 14368
rect 48319 14359 48377 14365
rect 48590 14356 48596 14368
rect 48648 14396 48654 14408
rect 48884 14396 48912 14427
rect 49142 14396 49148 14408
rect 48648 14368 48912 14396
rect 49103 14368 49148 14396
rect 48648 14356 48654 14368
rect 49142 14356 49148 14368
rect 49200 14356 49206 14408
rect 50540 14405 50568 14436
rect 51994 14424 52000 14436
rect 52052 14424 52058 14476
rect 50525 14399 50583 14405
rect 50525 14365 50537 14399
rect 50571 14365 50583 14399
rect 50525 14359 50583 14365
rect 50709 14399 50767 14405
rect 50709 14365 50721 14399
rect 50755 14396 50767 14399
rect 50890 14396 50896 14408
rect 50755 14368 50896 14396
rect 50755 14365 50767 14368
rect 50709 14359 50767 14365
rect 50890 14356 50896 14368
rect 50948 14356 50954 14408
rect 51074 14396 51080 14408
rect 51035 14368 51080 14396
rect 51074 14356 51080 14368
rect 51132 14356 51138 14408
rect 52104 14405 52132 14504
rect 52380 14504 56088 14532
rect 52178 14424 52184 14476
rect 52236 14464 52242 14476
rect 52380 14464 52408 14504
rect 56410 14492 56416 14544
rect 56468 14532 56474 14544
rect 58342 14532 58348 14544
rect 56468 14504 58348 14532
rect 56468 14492 56474 14504
rect 58342 14492 58348 14504
rect 58400 14492 58406 14544
rect 59630 14492 59636 14544
rect 59688 14532 59694 14544
rect 61013 14535 61071 14541
rect 61013 14532 61025 14535
rect 59688 14504 61025 14532
rect 59688 14492 59694 14504
rect 61013 14501 61025 14504
rect 61059 14501 61071 14535
rect 61013 14495 61071 14501
rect 61838 14492 61844 14544
rect 61896 14532 61902 14544
rect 62022 14532 62028 14544
rect 61896 14504 62028 14532
rect 61896 14492 61902 14504
rect 62022 14492 62028 14504
rect 62080 14492 62086 14544
rect 70305 14535 70363 14541
rect 70305 14501 70317 14535
rect 70351 14532 70363 14535
rect 70394 14532 70400 14544
rect 70351 14504 70400 14532
rect 70351 14501 70363 14504
rect 70305 14495 70363 14501
rect 70394 14492 70400 14504
rect 70452 14492 70458 14544
rect 70762 14532 70768 14544
rect 70723 14504 70768 14532
rect 70762 14492 70768 14504
rect 70820 14492 70826 14544
rect 72237 14535 72295 14541
rect 72237 14501 72249 14535
rect 72283 14532 72295 14535
rect 73430 14532 73436 14544
rect 72283 14504 73436 14532
rect 72283 14501 72295 14504
rect 72237 14495 72295 14501
rect 73430 14492 73436 14504
rect 73488 14492 73494 14544
rect 80026 14532 80054 14572
rect 87230 14532 87236 14544
rect 80026 14504 87236 14532
rect 87230 14492 87236 14504
rect 87288 14492 87294 14544
rect 53837 14467 53895 14473
rect 53837 14464 53849 14467
rect 52236 14436 52408 14464
rect 52656 14436 53849 14464
rect 52236 14424 52242 14436
rect 52656 14405 52684 14436
rect 53837 14433 53849 14436
rect 53883 14433 53895 14467
rect 53837 14427 53895 14433
rect 54478 14424 54484 14476
rect 54536 14464 54542 14476
rect 54846 14464 54852 14476
rect 54536 14436 54852 14464
rect 54536 14424 54542 14436
rect 54846 14424 54852 14436
rect 54904 14424 54910 14476
rect 54938 14424 54944 14476
rect 54996 14464 55002 14476
rect 55677 14467 55735 14473
rect 55677 14464 55689 14467
rect 54996 14436 55689 14464
rect 54996 14424 55002 14436
rect 55677 14433 55689 14436
rect 55723 14433 55735 14467
rect 55677 14427 55735 14433
rect 51261 14399 51319 14405
rect 51261 14365 51273 14399
rect 51307 14365 51319 14399
rect 51261 14359 51319 14365
rect 52089 14399 52147 14405
rect 52089 14365 52101 14399
rect 52135 14396 52147 14399
rect 52641 14399 52699 14405
rect 52641 14396 52653 14399
rect 52135 14368 52653 14396
rect 52135 14365 52147 14368
rect 52089 14359 52147 14365
rect 52641 14365 52653 14368
rect 52687 14365 52699 14399
rect 52914 14396 52920 14408
rect 52827 14368 52920 14396
rect 52641 14359 52699 14365
rect 50430 14328 50436 14340
rect 46216 14300 50436 14328
rect 43680 14288 43686 14300
rect 50430 14288 50436 14300
rect 50488 14288 50494 14340
rect 51276 14328 51304 14359
rect 52914 14356 52920 14368
rect 52972 14356 52978 14408
rect 54110 14396 54116 14408
rect 54071 14368 54116 14396
rect 54110 14356 54116 14368
rect 54168 14356 54174 14408
rect 54662 14356 54668 14408
rect 54720 14396 54726 14408
rect 55309 14399 55367 14405
rect 55309 14396 55321 14399
rect 54720 14368 55321 14396
rect 54720 14356 54726 14368
rect 55309 14365 55321 14368
rect 55355 14365 55367 14399
rect 55692 14396 55720 14427
rect 56502 14424 56508 14476
rect 56560 14464 56566 14476
rect 58158 14464 58164 14476
rect 56560 14436 58164 14464
rect 56560 14424 56566 14436
rect 58158 14424 58164 14436
rect 58216 14424 58222 14476
rect 58253 14467 58311 14473
rect 58253 14433 58265 14467
rect 58299 14464 58311 14467
rect 58434 14464 58440 14476
rect 58299 14436 58440 14464
rect 58299 14433 58311 14436
rect 58253 14427 58311 14433
rect 58434 14424 58440 14436
rect 58492 14424 58498 14476
rect 58618 14464 58624 14476
rect 58579 14436 58624 14464
rect 58618 14424 58624 14436
rect 58676 14424 58682 14476
rect 59906 14424 59912 14476
rect 59964 14464 59970 14476
rect 61473 14467 61531 14473
rect 61473 14464 61485 14467
rect 59964 14436 60596 14464
rect 59964 14424 59970 14436
rect 57974 14396 57980 14408
rect 55692 14368 57980 14396
rect 55309 14359 55367 14365
rect 57974 14356 57980 14368
rect 58032 14356 58038 14408
rect 58066 14356 58072 14408
rect 58124 14396 58130 14408
rect 60458 14396 60464 14408
rect 58124 14368 59124 14396
rect 60419 14368 60464 14396
rect 58124 14356 58130 14368
rect 50540 14300 51304 14328
rect 52932 14328 52960 14356
rect 59096 14340 59124 14368
rect 60458 14356 60464 14368
rect 60516 14356 60522 14408
rect 53926 14328 53932 14340
rect 52932 14300 53932 14328
rect 35989 14263 36047 14269
rect 35989 14260 36001 14263
rect 35636 14232 36001 14260
rect 35345 14223 35403 14229
rect 35989 14229 36001 14232
rect 36035 14260 36047 14263
rect 36998 14260 37004 14272
rect 36035 14232 37004 14260
rect 36035 14229 36047 14232
rect 35989 14223 36047 14229
rect 36998 14220 37004 14232
rect 37056 14220 37062 14272
rect 37090 14220 37096 14272
rect 37148 14260 37154 14272
rect 38657 14263 38715 14269
rect 38657 14260 38669 14263
rect 37148 14232 38669 14260
rect 37148 14220 37154 14232
rect 38657 14229 38669 14232
rect 38703 14229 38715 14263
rect 38657 14223 38715 14229
rect 40770 14220 40776 14272
rect 40828 14260 40834 14272
rect 42797 14263 42855 14269
rect 42797 14260 42809 14263
rect 40828 14232 42809 14260
rect 40828 14220 40834 14232
rect 42797 14229 42809 14232
rect 42843 14229 42855 14263
rect 42797 14223 42855 14229
rect 42978 14220 42984 14272
rect 43036 14260 43042 14272
rect 47486 14260 47492 14272
rect 43036 14232 47492 14260
rect 43036 14220 43042 14232
rect 47486 14220 47492 14232
rect 47544 14220 47550 14272
rect 47670 14260 47676 14272
rect 47631 14232 47676 14260
rect 47670 14220 47676 14232
rect 47728 14220 47734 14272
rect 48406 14260 48412 14272
rect 48367 14232 48412 14260
rect 48406 14220 48412 14232
rect 48464 14220 48470 14272
rect 48498 14220 48504 14272
rect 48556 14260 48562 14272
rect 49050 14260 49056 14272
rect 48556 14232 49056 14260
rect 48556 14220 48562 14232
rect 49050 14220 49056 14232
rect 49108 14220 49114 14272
rect 49510 14220 49516 14272
rect 49568 14260 49574 14272
rect 50540 14260 50568 14300
rect 53926 14288 53932 14300
rect 53984 14288 53990 14340
rect 55214 14288 55220 14340
rect 55272 14328 55278 14340
rect 56594 14328 56600 14340
rect 55272 14300 56600 14328
rect 55272 14288 55278 14300
rect 56594 14288 56600 14300
rect 56652 14288 56658 14340
rect 56778 14328 56784 14340
rect 56739 14300 56784 14328
rect 56778 14288 56784 14300
rect 56836 14288 56842 14340
rect 56962 14288 56968 14340
rect 57020 14328 57026 14340
rect 57425 14331 57483 14337
rect 57425 14328 57437 14331
rect 57020 14300 57437 14328
rect 57020 14288 57026 14300
rect 57425 14297 57437 14300
rect 57471 14297 57483 14331
rect 57425 14291 57483 14297
rect 57609 14331 57667 14337
rect 57609 14297 57621 14331
rect 57655 14328 57667 14331
rect 57790 14328 57796 14340
rect 57655 14300 57796 14328
rect 57655 14297 57667 14300
rect 57609 14291 57667 14297
rect 57790 14288 57796 14300
rect 57848 14288 57854 14340
rect 58158 14288 58164 14340
rect 58216 14328 58222 14340
rect 58866 14331 58924 14337
rect 58866 14328 58878 14331
rect 58216 14300 58878 14328
rect 58216 14288 58222 14300
rect 58866 14297 58878 14300
rect 58912 14297 58924 14331
rect 58866 14291 58924 14297
rect 59078 14288 59084 14340
rect 59136 14288 59142 14340
rect 60366 14328 60372 14340
rect 59556 14300 60372 14328
rect 49568 14232 50568 14260
rect 49568 14220 49574 14232
rect 50614 14220 50620 14272
rect 50672 14260 50678 14272
rect 51169 14263 51227 14269
rect 51169 14260 51181 14263
rect 50672 14232 51181 14260
rect 50672 14220 50678 14232
rect 51169 14229 51181 14232
rect 51215 14260 51227 14263
rect 55674 14260 55680 14272
rect 51215 14232 55680 14260
rect 51215 14229 51227 14232
rect 51169 14223 51227 14229
rect 55674 14220 55680 14232
rect 55732 14220 55738 14272
rect 56873 14263 56931 14269
rect 56873 14229 56885 14263
rect 56919 14260 56931 14263
rect 57238 14260 57244 14272
rect 56919 14232 57244 14260
rect 56919 14229 56931 14232
rect 56873 14223 56931 14229
rect 57238 14220 57244 14232
rect 57296 14220 57302 14272
rect 57808 14260 57836 14288
rect 59556 14260 59584 14300
rect 60366 14288 60372 14300
rect 60424 14288 60430 14340
rect 60568 14328 60596 14436
rect 60660 14436 61485 14464
rect 60660 14405 60688 14436
rect 61473 14433 61485 14436
rect 61519 14433 61531 14467
rect 62114 14464 62120 14476
rect 61473 14427 61531 14433
rect 61672 14436 62120 14464
rect 60918 14405 60924 14408
rect 60645 14399 60703 14405
rect 60645 14365 60657 14399
rect 60691 14365 60703 14399
rect 60645 14359 60703 14365
rect 60881 14399 60924 14405
rect 60881 14365 60893 14399
rect 60976 14396 60982 14408
rect 61286 14396 61292 14408
rect 60976 14368 61292 14396
rect 60881 14359 60924 14365
rect 60918 14356 60924 14359
rect 60976 14356 60982 14368
rect 61286 14356 61292 14368
rect 61344 14356 61350 14408
rect 61672 14405 61700 14436
rect 62114 14424 62120 14436
rect 62172 14424 62178 14476
rect 64598 14424 64604 14476
rect 64656 14424 64662 14476
rect 64966 14464 64972 14476
rect 64708 14436 64972 14464
rect 61657 14399 61715 14405
rect 61657 14365 61669 14399
rect 61703 14365 61715 14399
rect 61657 14359 61715 14365
rect 61746 14356 61752 14408
rect 61804 14396 61810 14408
rect 61933 14399 61991 14405
rect 61933 14396 61945 14399
rect 61804 14368 61945 14396
rect 61804 14356 61810 14368
rect 61933 14365 61945 14368
rect 61979 14365 61991 14399
rect 61933 14359 61991 14365
rect 62022 14356 62028 14408
rect 62080 14396 62086 14408
rect 62485 14399 62543 14405
rect 62485 14396 62497 14399
rect 62080 14368 62497 14396
rect 62080 14356 62086 14368
rect 62485 14365 62497 14368
rect 62531 14365 62543 14399
rect 62666 14396 62672 14408
rect 62627 14368 62672 14396
rect 62485 14359 62543 14365
rect 62666 14356 62672 14368
rect 62724 14356 62730 14408
rect 62761 14399 62819 14405
rect 62761 14365 62773 14399
rect 62807 14365 62819 14399
rect 62761 14359 62819 14365
rect 60737 14331 60795 14337
rect 60737 14328 60749 14331
rect 60568 14300 60749 14328
rect 60737 14297 60749 14300
rect 60783 14297 60795 14331
rect 61841 14331 61899 14337
rect 61841 14328 61853 14331
rect 60737 14291 60795 14297
rect 61304 14300 61853 14328
rect 57808 14232 59584 14260
rect 60001 14263 60059 14269
rect 60001 14229 60013 14263
rect 60047 14260 60059 14263
rect 61304 14260 61332 14300
rect 61841 14297 61853 14300
rect 61887 14297 61899 14331
rect 62776 14328 62804 14359
rect 63770 14356 63776 14408
rect 63828 14396 63834 14408
rect 63954 14396 63960 14408
rect 63828 14368 63873 14396
rect 63915 14368 63960 14396
rect 63828 14356 63834 14368
rect 63954 14356 63960 14368
rect 64012 14356 64018 14408
rect 64046 14356 64052 14408
rect 64104 14396 64110 14408
rect 64414 14396 64420 14408
rect 64104 14368 64149 14396
rect 64375 14368 64420 14396
rect 64104 14356 64110 14368
rect 64414 14356 64420 14368
rect 64472 14356 64478 14408
rect 64616 14337 64644 14424
rect 64708 14405 64736 14436
rect 64966 14424 64972 14436
rect 65024 14464 65030 14476
rect 65334 14464 65340 14476
rect 65024 14436 65340 14464
rect 65024 14424 65030 14436
rect 65334 14424 65340 14436
rect 65392 14424 65398 14476
rect 67450 14424 67456 14476
rect 67508 14464 67514 14476
rect 68922 14464 68928 14476
rect 67508 14436 68804 14464
rect 68883 14436 68928 14464
rect 67508 14424 67514 14436
rect 64689 14399 64747 14405
rect 64689 14365 64701 14399
rect 64735 14365 64747 14399
rect 64689 14359 64747 14365
rect 64785 14399 64843 14405
rect 64785 14365 64797 14399
rect 64831 14365 64843 14399
rect 64785 14359 64843 14365
rect 66441 14399 66499 14405
rect 66441 14365 66453 14399
rect 66487 14396 66499 14399
rect 66530 14396 66536 14408
rect 66487 14368 66536 14396
rect 66487 14365 66499 14368
rect 66441 14359 66499 14365
rect 64601 14331 64659 14337
rect 62776 14300 64184 14328
rect 61841 14291 61899 14297
rect 64156 14272 64184 14300
rect 64601 14297 64613 14331
rect 64647 14297 64659 14331
rect 64800 14328 64828 14359
rect 66530 14356 66536 14368
rect 66588 14356 66594 14408
rect 66714 14405 66720 14408
rect 66708 14359 66720 14405
rect 66772 14396 66778 14408
rect 68373 14399 68431 14405
rect 66772 14368 66808 14396
rect 66714 14356 66720 14359
rect 66772 14356 66778 14368
rect 68373 14365 68385 14399
rect 68419 14365 68431 14399
rect 68776 14396 68804 14436
rect 68922 14424 68928 14436
rect 68980 14424 68986 14476
rect 70026 14424 70032 14476
rect 70084 14464 70090 14476
rect 71317 14467 71375 14473
rect 71317 14464 71329 14467
rect 70084 14436 71329 14464
rect 70084 14424 70090 14436
rect 71317 14433 71329 14436
rect 71363 14433 71375 14467
rect 82814 14464 82820 14476
rect 71317 14427 71375 14433
rect 74736 14436 82820 14464
rect 68776 14368 69428 14396
rect 68373 14359 68431 14365
rect 64601 14291 64659 14297
rect 64717 14300 64828 14328
rect 68388 14328 68416 14359
rect 68646 14328 68652 14340
rect 68388 14300 68652 14328
rect 60047 14232 61332 14260
rect 60047 14229 60059 14232
rect 60001 14223 60059 14229
rect 61378 14220 61384 14272
rect 61436 14260 61442 14272
rect 62301 14263 62359 14269
rect 62301 14260 62313 14263
rect 61436 14232 62313 14260
rect 61436 14220 61442 14232
rect 62301 14229 62313 14232
rect 62347 14229 62359 14263
rect 63586 14260 63592 14272
rect 63547 14232 63592 14260
rect 62301 14223 62359 14229
rect 63586 14220 63592 14232
rect 63644 14220 63650 14272
rect 64138 14220 64144 14272
rect 64196 14260 64202 14272
rect 64717 14260 64745 14300
rect 68646 14288 68652 14300
rect 68704 14288 68710 14340
rect 69198 14337 69204 14340
rect 69192 14291 69204 14337
rect 69256 14328 69262 14340
rect 69256 14300 69292 14328
rect 69198 14288 69204 14291
rect 69256 14288 69262 14300
rect 64966 14260 64972 14272
rect 64196 14232 64745 14260
rect 64927 14232 64972 14260
rect 64196 14220 64202 14232
rect 64966 14220 64972 14232
rect 65024 14220 65030 14272
rect 67821 14263 67879 14269
rect 67821 14229 67833 14263
rect 67867 14260 67879 14263
rect 68370 14260 68376 14272
rect 67867 14232 68376 14260
rect 67867 14229 67879 14232
rect 67821 14223 67879 14229
rect 68370 14220 68376 14232
rect 68428 14220 68434 14272
rect 68462 14220 68468 14272
rect 68520 14260 68526 14272
rect 69400 14260 69428 14368
rect 70302 14356 70308 14408
rect 70360 14396 70366 14408
rect 71133 14399 71191 14405
rect 71133 14396 71145 14399
rect 70360 14368 71145 14396
rect 70360 14356 70366 14368
rect 71133 14365 71145 14368
rect 71179 14365 71191 14399
rect 71133 14359 71191 14365
rect 71225 14399 71283 14405
rect 71225 14365 71237 14399
rect 71271 14396 71283 14399
rect 74736 14396 74764 14436
rect 82814 14424 82820 14436
rect 82872 14424 82878 14476
rect 71271 14368 74764 14396
rect 71271 14365 71283 14368
rect 71225 14359 71283 14365
rect 74810 14356 74816 14408
rect 74868 14396 74874 14408
rect 84838 14396 84844 14408
rect 74868 14368 84844 14396
rect 74868 14356 74874 14368
rect 84838 14356 84844 14368
rect 84896 14356 84902 14408
rect 69474 14288 69480 14340
rect 69532 14328 69538 14340
rect 71869 14331 71927 14337
rect 71869 14328 71881 14331
rect 69532 14300 71881 14328
rect 69532 14288 69538 14300
rect 71869 14297 71881 14300
rect 71915 14297 71927 14331
rect 72050 14328 72056 14340
rect 72011 14300 72056 14328
rect 71869 14291 71927 14297
rect 72050 14288 72056 14300
rect 72108 14288 72114 14340
rect 88058 14328 88064 14340
rect 88019 14300 88064 14328
rect 88058 14288 88064 14300
rect 88116 14288 88122 14340
rect 73706 14260 73712 14272
rect 68520 14232 68565 14260
rect 69400 14232 73712 14260
rect 68520 14220 68526 14232
rect 73706 14220 73712 14232
rect 73764 14220 73770 14272
rect 88150 14260 88156 14272
rect 88111 14232 88156 14260
rect 88150 14220 88156 14232
rect 88208 14220 88214 14272
rect 1104 14170 88872 14192
rect 1104 14118 22898 14170
rect 22950 14118 22962 14170
rect 23014 14118 23026 14170
rect 23078 14118 23090 14170
rect 23142 14118 23154 14170
rect 23206 14118 44846 14170
rect 44898 14118 44910 14170
rect 44962 14118 44974 14170
rect 45026 14118 45038 14170
rect 45090 14118 45102 14170
rect 45154 14118 66794 14170
rect 66846 14118 66858 14170
rect 66910 14118 66922 14170
rect 66974 14118 66986 14170
rect 67038 14118 67050 14170
rect 67102 14118 88872 14170
rect 1104 14096 88872 14118
rect 2869 14059 2927 14065
rect 2869 14025 2881 14059
rect 2915 14025 2927 14059
rect 2869 14019 2927 14025
rect 19429 14059 19487 14065
rect 19429 14025 19441 14059
rect 19475 14056 19487 14059
rect 20993 14059 21051 14065
rect 20993 14056 21005 14059
rect 19475 14028 21005 14056
rect 19475 14025 19487 14028
rect 19429 14019 19487 14025
rect 20993 14025 21005 14028
rect 21039 14025 21051 14059
rect 20993 14019 21051 14025
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 2884 13920 2912 14019
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 23474 14056 23480 14068
rect 21232 14028 23480 14056
rect 21232 14016 21238 14028
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 23658 14016 23664 14068
rect 23716 14056 23722 14068
rect 24302 14056 24308 14068
rect 23716 14028 24308 14056
rect 23716 14016 23722 14028
rect 24302 14016 24308 14028
rect 24360 14016 24366 14068
rect 24394 14016 24400 14068
rect 24452 14056 24458 14068
rect 24765 14059 24823 14065
rect 24765 14056 24777 14059
rect 24452 14028 24777 14056
rect 24452 14016 24458 14028
rect 24765 14025 24777 14028
rect 24811 14025 24823 14059
rect 24765 14019 24823 14025
rect 24946 14016 24952 14068
rect 25004 14056 25010 14068
rect 26418 14056 26424 14068
rect 25004 14028 26424 14056
rect 25004 14016 25010 14028
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 26510 14016 26516 14068
rect 26568 14056 26574 14068
rect 28537 14059 28595 14065
rect 28537 14056 28549 14059
rect 26568 14028 28549 14056
rect 26568 14016 26574 14028
rect 28537 14025 28549 14028
rect 28583 14025 28595 14059
rect 29086 14056 29092 14068
rect 29047 14028 29092 14056
rect 28537 14019 28595 14025
rect 29086 14016 29092 14028
rect 29144 14056 29150 14068
rect 29362 14056 29368 14068
rect 29144 14028 29368 14056
rect 29144 14016 29150 14028
rect 29362 14016 29368 14028
rect 29420 14016 29426 14068
rect 29638 14016 29644 14068
rect 29696 14056 29702 14068
rect 34241 14059 34299 14065
rect 29696 14028 33824 14056
rect 29696 14016 29702 14028
rect 20438 13988 20444 14000
rect 6886 13960 20444 13988
rect 1627 13892 2912 13920
rect 3053 13923 3111 13929
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 3053 13889 3065 13923
rect 3099 13920 3111 13923
rect 6886 13920 6914 13960
rect 20438 13948 20444 13960
rect 20496 13948 20502 14000
rect 21358 13988 21364 14000
rect 20916 13960 21364 13988
rect 3099 13892 6914 13920
rect 18141 13923 18199 13929
rect 3099 13889 3111 13892
rect 3053 13883 3111 13889
rect 18141 13889 18153 13923
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 18156 13784 18184 13883
rect 18230 13880 18236 13932
rect 18288 13920 18294 13932
rect 18969 13923 19027 13929
rect 18969 13920 18981 13923
rect 18288 13892 18981 13920
rect 18288 13880 18294 13892
rect 18969 13889 18981 13892
rect 19015 13889 19027 13923
rect 19794 13920 19800 13932
rect 19755 13892 19800 13920
rect 18969 13883 19027 13889
rect 19794 13880 19800 13892
rect 19852 13880 19858 13932
rect 20916 13929 20944 13960
rect 21358 13948 21364 13960
rect 21416 13948 21422 14000
rect 21542 13948 21548 14000
rect 21600 13988 21606 14000
rect 26145 13991 26203 13997
rect 21600 13960 25360 13988
rect 21600 13948 21606 13960
rect 20901 13923 20959 13929
rect 20901 13889 20913 13923
rect 20947 13889 20959 13923
rect 20901 13883 20959 13889
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13920 21143 13923
rect 22738 13920 22744 13932
rect 21131 13892 22744 13920
rect 21131 13889 21143 13892
rect 21085 13883 21143 13889
rect 22738 13880 22744 13892
rect 22796 13880 22802 13932
rect 22830 13880 22836 13932
rect 22888 13920 22894 13932
rect 23017 13923 23075 13929
rect 23017 13920 23029 13923
rect 22888 13892 23029 13920
rect 22888 13880 22894 13892
rect 23017 13889 23029 13892
rect 23063 13889 23075 13923
rect 23017 13883 23075 13889
rect 23201 13923 23259 13929
rect 23201 13889 23213 13923
rect 23247 13889 23259 13923
rect 23842 13920 23848 13932
rect 23803 13892 23848 13920
rect 23201 13883 23259 13889
rect 18601 13855 18659 13861
rect 18601 13821 18613 13855
rect 18647 13852 18659 13855
rect 19610 13852 19616 13864
rect 18647 13824 19616 13852
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 20257 13855 20315 13861
rect 20257 13821 20269 13855
rect 20303 13852 20315 13855
rect 21174 13852 21180 13864
rect 20303 13824 21180 13852
rect 20303 13821 20315 13824
rect 20257 13815 20315 13821
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 21361 13855 21419 13861
rect 21361 13821 21373 13855
rect 21407 13852 21419 13855
rect 22186 13852 22192 13864
rect 21407 13824 22192 13852
rect 21407 13821 21419 13824
rect 21361 13815 21419 13821
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 22278 13812 22284 13864
rect 22336 13852 22342 13864
rect 23216 13852 23244 13883
rect 23842 13880 23848 13892
rect 23900 13880 23906 13932
rect 24670 13920 24676 13932
rect 24631 13892 24676 13920
rect 24670 13880 24676 13892
rect 24728 13880 24734 13932
rect 25222 13920 25228 13932
rect 25183 13892 25228 13920
rect 25222 13880 25228 13892
rect 25280 13880 25286 13932
rect 25332 13929 25360 13960
rect 26145 13957 26157 13991
rect 26191 13988 26203 13991
rect 26191 13960 26556 13988
rect 26191 13957 26203 13960
rect 26145 13951 26203 13957
rect 25317 13923 25375 13929
rect 25317 13889 25329 13923
rect 25363 13889 25375 13923
rect 25961 13923 26019 13929
rect 25961 13920 25973 13923
rect 25317 13883 25375 13889
rect 25424 13892 25973 13920
rect 22336 13824 23244 13852
rect 22336 13812 22342 13824
rect 23290 13812 23296 13864
rect 23348 13852 23354 13864
rect 23661 13855 23719 13861
rect 23661 13852 23673 13855
rect 23348 13824 23673 13852
rect 23348 13812 23354 13824
rect 23661 13821 23673 13824
rect 23707 13821 23719 13855
rect 23661 13815 23719 13821
rect 23753 13855 23811 13861
rect 23753 13821 23765 13855
rect 23799 13821 23811 13855
rect 23753 13815 23811 13821
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 24578 13852 24584 13864
rect 24167 13824 24584 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 20806 13784 20812 13796
rect 18156 13756 19196 13784
rect 20767 13756 20812 13784
rect 19168 13728 19196 13756
rect 20806 13744 20812 13756
rect 20864 13744 20870 13796
rect 22094 13784 22100 13796
rect 20916 13756 22100 13784
rect 1394 13716 1400 13728
rect 1355 13688 1400 13716
rect 1394 13676 1400 13688
rect 1452 13676 1458 13728
rect 18230 13716 18236 13728
rect 18191 13688 18236 13716
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 19150 13716 19156 13728
rect 19111 13688 19156 13716
rect 19150 13676 19156 13688
rect 19208 13676 19214 13728
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 19889 13719 19947 13725
rect 19889 13716 19901 13719
rect 19576 13688 19901 13716
rect 19576 13676 19582 13688
rect 19889 13685 19901 13688
rect 19935 13716 19947 13719
rect 20916 13716 20944 13756
rect 22094 13744 22100 13756
rect 22152 13744 22158 13796
rect 22554 13744 22560 13796
rect 22612 13784 22618 13796
rect 22833 13787 22891 13793
rect 22833 13784 22845 13787
rect 22612 13756 22845 13784
rect 22612 13744 22618 13756
rect 22833 13753 22845 13756
rect 22879 13753 22891 13787
rect 23566 13784 23572 13796
rect 23527 13756 23572 13784
rect 22833 13747 22891 13753
rect 23566 13744 23572 13756
rect 23624 13744 23630 13796
rect 23768 13728 23796 13815
rect 24578 13812 24584 13824
rect 24636 13812 24642 13864
rect 25424 13852 25452 13892
rect 25961 13889 25973 13892
rect 26007 13889 26019 13923
rect 26234 13920 26240 13932
rect 26195 13892 26240 13920
rect 25961 13883 26019 13889
rect 26234 13880 26240 13892
rect 26292 13880 26298 13932
rect 26326 13880 26332 13932
rect 26384 13920 26390 13932
rect 26528 13920 26556 13960
rect 26602 13948 26608 14000
rect 26660 13988 26666 14000
rect 28074 13988 28080 14000
rect 26660 13960 28080 13988
rect 26660 13948 26666 13960
rect 28074 13948 28080 13960
rect 28132 13948 28138 14000
rect 28997 13991 29055 13997
rect 28997 13957 29009 13991
rect 29043 13988 29055 13991
rect 29178 13988 29184 14000
rect 29043 13960 29184 13988
rect 29043 13957 29055 13960
rect 28997 13951 29055 13957
rect 29178 13948 29184 13960
rect 29236 13988 29242 14000
rect 30834 13988 30840 14000
rect 29236 13960 30840 13988
rect 29236 13948 29242 13960
rect 30834 13948 30840 13960
rect 30892 13948 30898 14000
rect 31478 13988 31484 14000
rect 31439 13960 31484 13988
rect 31478 13948 31484 13960
rect 31536 13948 31542 14000
rect 31662 13948 31668 14000
rect 31720 13988 31726 14000
rect 32306 13988 32312 14000
rect 31720 13960 32312 13988
rect 31720 13948 31726 13960
rect 32306 13948 32312 13960
rect 32364 13948 32370 14000
rect 33410 13948 33416 14000
rect 33468 13988 33474 14000
rect 33505 13991 33563 13997
rect 33505 13988 33517 13991
rect 33468 13960 33517 13988
rect 33468 13948 33474 13960
rect 33505 13957 33517 13960
rect 33551 13988 33563 13991
rect 33686 13988 33692 14000
rect 33551 13960 33692 13988
rect 33551 13957 33563 13960
rect 33505 13951 33563 13957
rect 33686 13948 33692 13960
rect 33744 13948 33750 14000
rect 33796 13988 33824 14028
rect 34241 14025 34253 14059
rect 34287 14056 34299 14059
rect 34790 14056 34796 14068
rect 34287 14028 34796 14056
rect 34287 14025 34299 14028
rect 34241 14019 34299 14025
rect 34790 14016 34796 14028
rect 34848 14016 34854 14068
rect 35434 14056 35440 14068
rect 34900 14028 35440 14056
rect 34900 13988 34928 14028
rect 35434 14016 35440 14028
rect 35492 14016 35498 14068
rect 35638 14059 35696 14065
rect 35638 14025 35650 14059
rect 35684 14056 35696 14059
rect 36081 14059 36139 14065
rect 36081 14056 36093 14059
rect 35684 14028 36093 14056
rect 35684 14025 35696 14028
rect 35638 14019 35696 14025
rect 36081 14025 36093 14028
rect 36127 14056 36139 14059
rect 36170 14056 36176 14068
rect 36127 14028 36176 14056
rect 36127 14025 36139 14028
rect 36081 14019 36139 14025
rect 36170 14016 36176 14028
rect 36228 14016 36234 14068
rect 37918 14016 37924 14068
rect 37976 14056 37982 14068
rect 38746 14056 38752 14068
rect 37976 14028 38752 14056
rect 37976 14016 37982 14028
rect 38746 14016 38752 14028
rect 38804 14016 38810 14068
rect 39298 14056 39304 14068
rect 39151 14028 39304 14056
rect 33796 13960 34928 13988
rect 37461 13991 37519 13997
rect 37461 13957 37473 13991
rect 37507 13988 37519 13991
rect 38838 13988 38844 14000
rect 37507 13960 38844 13988
rect 37507 13957 37519 13960
rect 37461 13951 37519 13957
rect 38838 13948 38844 13960
rect 38896 13948 38902 14000
rect 26694 13920 26700 13932
rect 26384 13892 26429 13920
rect 26528 13892 26700 13920
rect 26384 13880 26390 13892
rect 26694 13880 26700 13892
rect 26752 13880 26758 13932
rect 26878 13880 26884 13932
rect 26936 13920 26942 13932
rect 27246 13920 27252 13932
rect 26936 13892 27252 13920
rect 26936 13880 26942 13892
rect 27246 13880 27252 13892
rect 27304 13920 27310 13932
rect 27341 13923 27399 13929
rect 27341 13920 27353 13923
rect 27304 13892 27353 13920
rect 27304 13880 27310 13892
rect 27341 13889 27353 13892
rect 27387 13920 27399 13923
rect 27387 13892 28994 13920
rect 27387 13889 27399 13892
rect 27341 13883 27399 13889
rect 28092 13864 28120 13892
rect 24688 13824 25452 13852
rect 24486 13744 24492 13796
rect 24544 13784 24550 13796
rect 24688 13784 24716 13824
rect 25774 13812 25780 13864
rect 25832 13852 25838 13864
rect 27430 13852 27436 13864
rect 25832 13824 27016 13852
rect 27391 13824 27436 13852
rect 25832 13812 25838 13824
rect 26513 13787 26571 13793
rect 26513 13784 26525 13787
rect 24544 13756 24716 13784
rect 25424 13756 26525 13784
rect 24544 13744 24550 13756
rect 21266 13716 21272 13728
rect 19935 13688 20944 13716
rect 21227 13688 21272 13716
rect 19935 13685 19947 13688
rect 19889 13679 19947 13685
rect 21266 13676 21272 13688
rect 21324 13716 21330 13728
rect 21726 13716 21732 13728
rect 21324 13688 21732 13716
rect 21324 13676 21330 13688
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 22462 13716 22468 13728
rect 22423 13688 22468 13716
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 22738 13716 22744 13728
rect 22699 13688 22744 13716
rect 22738 13676 22744 13688
rect 22796 13676 22802 13728
rect 22925 13719 22983 13725
rect 22925 13685 22937 13719
rect 22971 13716 22983 13719
rect 23658 13716 23664 13728
rect 22971 13688 23664 13716
rect 22971 13685 22983 13688
rect 22925 13679 22983 13685
rect 23658 13676 23664 13688
rect 23716 13676 23722 13728
rect 23750 13676 23756 13728
rect 23808 13676 23814 13728
rect 24026 13716 24032 13728
rect 23987 13688 24032 13716
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 25424 13725 25452 13756
rect 26513 13753 26525 13756
rect 26559 13753 26571 13787
rect 26513 13747 26571 13753
rect 26602 13744 26608 13796
rect 26660 13784 26666 13796
rect 26878 13784 26884 13796
rect 26660 13756 26884 13784
rect 26660 13744 26666 13756
rect 26878 13744 26884 13756
rect 26936 13744 26942 13796
rect 26988 13793 27016 13824
rect 27430 13812 27436 13824
rect 27488 13812 27494 13864
rect 27525 13855 27583 13861
rect 27525 13821 27537 13855
rect 27571 13821 27583 13855
rect 27525 13815 27583 13821
rect 26973 13787 27031 13793
rect 26973 13753 26985 13787
rect 27019 13753 27031 13787
rect 27540 13784 27568 13815
rect 28074 13812 28080 13864
rect 28132 13812 28138 13864
rect 27614 13784 27620 13796
rect 27540 13756 27620 13784
rect 26973 13747 27031 13753
rect 27614 13744 27620 13756
rect 27672 13744 27678 13796
rect 28445 13787 28503 13793
rect 28445 13753 28457 13787
rect 28491 13784 28503 13787
rect 28718 13784 28724 13796
rect 28491 13756 28724 13784
rect 28491 13753 28503 13756
rect 28445 13747 28503 13753
rect 25409 13719 25467 13725
rect 25409 13685 25421 13719
rect 25455 13685 25467 13719
rect 25409 13679 25467 13685
rect 25593 13719 25651 13725
rect 25593 13685 25605 13719
rect 25639 13716 25651 13719
rect 25682 13716 25688 13728
rect 25639 13688 25688 13716
rect 25639 13685 25651 13688
rect 25593 13679 25651 13685
rect 25682 13676 25688 13688
rect 25740 13676 25746 13728
rect 26418 13676 26424 13728
rect 26476 13716 26482 13728
rect 28460 13716 28488 13747
rect 28718 13744 28724 13756
rect 28776 13744 28782 13796
rect 28966 13784 28994 13892
rect 30098 13880 30104 13932
rect 30156 13920 30162 13932
rect 30193 13923 30251 13929
rect 30193 13920 30205 13923
rect 30156 13892 30205 13920
rect 30156 13880 30162 13892
rect 30193 13889 30205 13892
rect 30239 13889 30251 13923
rect 30193 13883 30251 13889
rect 31110 13880 31116 13932
rect 31168 13920 31174 13932
rect 31297 13923 31355 13929
rect 31297 13920 31309 13923
rect 31168 13892 31309 13920
rect 31168 13880 31174 13892
rect 31297 13889 31309 13892
rect 31343 13889 31355 13923
rect 32490 13920 32496 13932
rect 32451 13892 32496 13920
rect 31297 13883 31355 13889
rect 32490 13880 32496 13892
rect 32548 13880 32554 13932
rect 32677 13923 32735 13929
rect 32677 13889 32689 13923
rect 32723 13920 32735 13923
rect 33134 13920 33140 13932
rect 32723 13892 33140 13920
rect 32723 13889 32735 13892
rect 32677 13883 32735 13889
rect 33134 13880 33140 13892
rect 33192 13880 33198 13932
rect 33229 13923 33287 13929
rect 33229 13889 33241 13923
rect 33275 13889 33287 13923
rect 34422 13920 34428 13932
rect 34383 13892 34428 13920
rect 33229 13883 33287 13889
rect 29822 13784 29828 13796
rect 28966 13756 29828 13784
rect 29822 13744 29828 13756
rect 29880 13744 29886 13796
rect 30377 13787 30435 13793
rect 30377 13753 30389 13787
rect 30423 13784 30435 13787
rect 31110 13784 31116 13796
rect 30423 13756 31116 13784
rect 30423 13753 30435 13756
rect 30377 13747 30435 13753
rect 31110 13744 31116 13756
rect 31168 13744 31174 13796
rect 33244 13784 33272 13883
rect 34422 13880 34428 13892
rect 34480 13880 34486 13932
rect 34793 13923 34851 13929
rect 34793 13889 34805 13923
rect 34839 13920 34851 13923
rect 34882 13920 34888 13932
rect 34839 13892 34888 13920
rect 34839 13889 34851 13892
rect 34793 13883 34851 13889
rect 34882 13880 34888 13892
rect 34940 13880 34946 13932
rect 35066 13920 35072 13932
rect 35027 13892 35072 13920
rect 35066 13880 35072 13892
rect 35124 13880 35130 13932
rect 35250 13920 35256 13932
rect 35211 13892 35256 13920
rect 35250 13880 35256 13892
rect 35308 13880 35314 13932
rect 35345 13923 35403 13929
rect 35345 13889 35357 13923
rect 35391 13889 35403 13923
rect 35345 13883 35403 13889
rect 33318 13784 33324 13796
rect 33244 13756 33324 13784
rect 33318 13744 33324 13756
rect 33376 13744 33382 13796
rect 33410 13744 33416 13796
rect 33468 13784 33474 13796
rect 35158 13784 35164 13796
rect 33468 13756 35164 13784
rect 33468 13744 33474 13756
rect 35158 13744 35164 13756
rect 35216 13744 35222 13796
rect 35360 13784 35388 13883
rect 35434 13880 35440 13932
rect 35492 13929 35498 13932
rect 35492 13923 35523 13929
rect 35511 13889 35523 13923
rect 35492 13883 35523 13889
rect 35492 13880 35498 13883
rect 35894 13880 35900 13932
rect 35952 13920 35958 13932
rect 37277 13923 37335 13929
rect 37277 13920 37289 13923
rect 35952 13892 37289 13920
rect 35952 13880 35958 13892
rect 37277 13889 37289 13892
rect 37323 13889 37335 13923
rect 37550 13920 37556 13932
rect 37511 13892 37556 13920
rect 37277 13883 37335 13889
rect 37550 13880 37556 13892
rect 37608 13880 37614 13932
rect 37734 13929 37740 13932
rect 37697 13923 37740 13929
rect 37697 13889 37709 13923
rect 37697 13883 37740 13889
rect 37734 13880 37740 13883
rect 37792 13880 37798 13932
rect 38286 13920 38292 13932
rect 38247 13892 38292 13920
rect 38286 13880 38292 13892
rect 38344 13880 38350 13932
rect 38378 13880 38384 13932
rect 38436 13920 38442 13932
rect 39151 13920 39179 14028
rect 39298 14016 39304 14028
rect 39356 14016 39362 14068
rect 39390 14016 39396 14068
rect 39448 14056 39454 14068
rect 40589 14059 40647 14065
rect 40589 14056 40601 14059
rect 39448 14028 40601 14056
rect 39448 14016 39454 14028
rect 40589 14025 40601 14028
rect 40635 14025 40647 14059
rect 41414 14056 41420 14068
rect 40589 14019 40647 14025
rect 40972 14028 41420 14056
rect 40972 13988 41000 14028
rect 41414 14016 41420 14028
rect 41472 14016 41478 14068
rect 41506 14016 41512 14068
rect 41564 14056 41570 14068
rect 41564 14028 50936 14056
rect 41564 14016 41570 14028
rect 38436 13892 39179 13920
rect 39224 13960 41000 13988
rect 41049 13991 41107 13997
rect 38436 13880 38442 13892
rect 39224 13852 39252 13960
rect 41049 13957 41061 13991
rect 41095 13988 41107 13991
rect 42518 13988 42524 14000
rect 41095 13960 42524 13988
rect 41095 13957 41107 13960
rect 41049 13951 41107 13957
rect 42518 13948 42524 13960
rect 42576 13948 42582 14000
rect 42702 13948 42708 14000
rect 42760 13988 42766 14000
rect 45830 13988 45836 14000
rect 42760 13960 45836 13988
rect 42760 13948 42766 13960
rect 40957 13923 41015 13929
rect 40221 13907 40279 13913
rect 40221 13873 40233 13907
rect 40267 13904 40279 13907
rect 40267 13876 40356 13904
rect 40957 13889 40969 13923
rect 41003 13920 41015 13923
rect 41322 13920 41328 13932
rect 41003 13892 41328 13920
rect 41003 13889 41015 13892
rect 40957 13883 41015 13889
rect 41322 13880 41328 13892
rect 41380 13880 41386 13932
rect 41690 13920 41696 13932
rect 41651 13892 41696 13920
rect 41690 13880 41696 13892
rect 41748 13880 41754 13932
rect 42613 13923 42671 13929
rect 42613 13889 42625 13923
rect 42659 13920 42671 13923
rect 42978 13920 42984 13932
rect 42659 13892 42984 13920
rect 42659 13889 42671 13892
rect 42613 13883 42671 13889
rect 42978 13880 42984 13892
rect 43036 13880 43042 13932
rect 43824 13929 43852 13960
rect 45830 13948 45836 13960
rect 45888 13948 45894 14000
rect 46385 13991 46443 13997
rect 46385 13957 46397 13991
rect 46431 13988 46443 13991
rect 47762 13988 47768 14000
rect 46431 13960 47768 13988
rect 46431 13957 46443 13960
rect 46385 13951 46443 13957
rect 47762 13948 47768 13960
rect 47820 13948 47826 14000
rect 48590 13988 48596 14000
rect 47964 13960 48596 13988
rect 43809 13923 43867 13929
rect 43809 13889 43821 13923
rect 43855 13889 43867 13923
rect 43809 13883 43867 13889
rect 44076 13923 44134 13929
rect 44076 13889 44088 13923
rect 44122 13920 44134 13923
rect 44358 13920 44364 13932
rect 44122 13892 44364 13920
rect 44122 13889 44134 13892
rect 44076 13883 44134 13889
rect 44358 13880 44364 13892
rect 44416 13880 44422 13932
rect 44542 13880 44548 13932
rect 44600 13920 44606 13932
rect 45741 13923 45799 13929
rect 44600 13892 45508 13920
rect 44600 13880 44606 13892
rect 40267 13873 40279 13876
rect 40221 13867 40279 13873
rect 39390 13852 39396 13864
rect 37660 13824 39252 13852
rect 39351 13824 39396 13852
rect 35802 13784 35808 13796
rect 35360 13756 35808 13784
rect 35802 13744 35808 13756
rect 35860 13784 35866 13796
rect 37550 13784 37556 13796
rect 35860 13756 37556 13784
rect 35860 13744 35866 13756
rect 37550 13744 37556 13756
rect 37608 13744 37614 13796
rect 26476 13688 28488 13716
rect 26476 13676 26482 13688
rect 28626 13676 28632 13728
rect 28684 13716 28690 13728
rect 30466 13716 30472 13728
rect 28684 13688 30472 13716
rect 28684 13676 28690 13688
rect 30466 13676 30472 13688
rect 30524 13676 30530 13728
rect 30742 13676 30748 13728
rect 30800 13716 30806 13728
rect 37660 13716 37688 13824
rect 39390 13812 39396 13824
rect 39448 13812 39454 13864
rect 39577 13855 39635 13861
rect 39577 13821 39589 13855
rect 39623 13821 39635 13855
rect 39577 13815 39635 13821
rect 38565 13787 38623 13793
rect 38565 13753 38577 13787
rect 38611 13784 38623 13787
rect 39408 13784 39436 13812
rect 38611 13756 39436 13784
rect 38611 13753 38623 13756
rect 38565 13747 38623 13753
rect 30800 13688 37688 13716
rect 37829 13719 37887 13725
rect 30800 13676 30806 13688
rect 37829 13685 37841 13719
rect 37875 13716 37887 13719
rect 37918 13716 37924 13728
rect 37875 13688 37924 13716
rect 37875 13685 37887 13688
rect 37829 13679 37887 13685
rect 37918 13676 37924 13688
rect 37976 13676 37982 13728
rect 38102 13716 38108 13728
rect 38063 13688 38108 13716
rect 38102 13676 38108 13688
rect 38160 13676 38166 13728
rect 38746 13676 38752 13728
rect 38804 13716 38810 13728
rect 38933 13719 38991 13725
rect 38933 13716 38945 13719
rect 38804 13688 38945 13716
rect 38804 13676 38810 13688
rect 38933 13685 38945 13688
rect 38979 13685 38991 13719
rect 39592 13716 39620 13815
rect 39758 13812 39764 13864
rect 39816 13852 39822 13864
rect 39942 13852 39948 13864
rect 39816 13824 39948 13852
rect 39816 13812 39822 13824
rect 39942 13812 39948 13824
rect 40000 13812 40006 13864
rect 40328 13852 40356 13876
rect 40328 13824 40448 13852
rect 40037 13787 40095 13793
rect 40037 13753 40049 13787
rect 40083 13784 40095 13787
rect 40310 13784 40316 13796
rect 40083 13756 40316 13784
rect 40083 13753 40095 13756
rect 40037 13747 40095 13753
rect 40310 13744 40316 13756
rect 40368 13744 40374 13796
rect 40420 13784 40448 13824
rect 41046 13812 41052 13864
rect 41104 13852 41110 13864
rect 41141 13855 41199 13861
rect 41141 13852 41153 13855
rect 41104 13824 41153 13852
rect 41104 13812 41110 13824
rect 41141 13821 41153 13824
rect 41187 13821 41199 13855
rect 41340 13852 41368 13880
rect 42058 13852 42064 13864
rect 41340 13824 42064 13852
rect 41141 13815 41199 13821
rect 42058 13812 42064 13824
rect 42116 13852 42122 13864
rect 42886 13852 42892 13864
rect 42116 13824 42288 13852
rect 42847 13824 42892 13852
rect 42116 13812 42122 13824
rect 40770 13784 40776 13796
rect 40420 13756 40776 13784
rect 40770 13744 40776 13756
rect 40828 13744 40834 13796
rect 41877 13787 41935 13793
rect 41877 13753 41889 13787
rect 41923 13784 41935 13787
rect 42150 13784 42156 13796
rect 41923 13756 42156 13784
rect 41923 13753 41935 13756
rect 41877 13747 41935 13753
rect 42150 13744 42156 13756
rect 42208 13744 42214 13796
rect 42260 13784 42288 13824
rect 42886 13812 42892 13824
rect 42944 13812 42950 13864
rect 45186 13812 45192 13864
rect 45244 13812 45250 13864
rect 43162 13784 43168 13796
rect 42260 13756 43168 13784
rect 43162 13744 43168 13756
rect 43220 13744 43226 13796
rect 41046 13716 41052 13728
rect 39592 13688 41052 13716
rect 38933 13679 38991 13685
rect 41046 13676 41052 13688
rect 41104 13676 41110 13728
rect 41138 13676 41144 13728
rect 41196 13716 41202 13728
rect 45094 13716 45100 13728
rect 41196 13688 45100 13716
rect 41196 13676 41202 13688
rect 45094 13676 45100 13688
rect 45152 13676 45158 13728
rect 45204 13725 45232 13812
rect 45189 13719 45247 13725
rect 45189 13685 45201 13719
rect 45235 13685 45247 13719
rect 45480 13716 45508 13892
rect 45741 13889 45753 13923
rect 45787 13920 45799 13923
rect 46014 13920 46020 13932
rect 45787 13892 46020 13920
rect 45787 13889 45799 13892
rect 45741 13883 45799 13889
rect 46014 13880 46020 13892
rect 46072 13880 46078 13932
rect 46474 13880 46480 13932
rect 46532 13920 46538 13932
rect 46569 13923 46627 13929
rect 46569 13920 46581 13923
rect 46532 13892 46581 13920
rect 46532 13880 46538 13892
rect 46569 13889 46581 13892
rect 46615 13889 46627 13923
rect 46569 13883 46627 13889
rect 46937 13923 46995 13929
rect 46937 13889 46949 13923
rect 46983 13920 46995 13923
rect 47964 13920 47992 13960
rect 48590 13948 48596 13960
rect 48648 13948 48654 14000
rect 48774 13948 48780 14000
rect 48832 13988 48838 14000
rect 49234 13988 49240 14000
rect 48832 13960 49240 13988
rect 48832 13948 48838 13960
rect 49234 13948 49240 13960
rect 49292 13948 49298 14000
rect 50154 13948 50160 14000
rect 50212 13948 50218 14000
rect 50246 13948 50252 14000
rect 50304 13988 50310 14000
rect 50798 13988 50804 14000
rect 50304 13960 50804 13988
rect 50304 13948 50310 13960
rect 50798 13948 50804 13960
rect 50856 13948 50862 14000
rect 50908 13988 50936 14028
rect 50982 14016 50988 14068
rect 51040 14056 51046 14068
rect 51169 14059 51227 14065
rect 51169 14056 51181 14059
rect 51040 14028 51181 14056
rect 51040 14016 51046 14028
rect 51169 14025 51181 14028
rect 51215 14025 51227 14059
rect 51169 14019 51227 14025
rect 51994 14016 52000 14068
rect 52052 14056 52058 14068
rect 57983 14059 58041 14065
rect 52052 14028 57560 14056
rect 52052 14016 52058 14028
rect 52730 13988 52736 14000
rect 50908 13960 52736 13988
rect 52730 13948 52736 13960
rect 52788 13948 52794 14000
rect 54570 13988 54576 14000
rect 52932 13960 54576 13988
rect 46983 13892 47992 13920
rect 46983 13889 46995 13892
rect 46937 13883 46995 13889
rect 48038 13880 48044 13932
rect 48096 13920 48102 13932
rect 48205 13923 48263 13929
rect 48205 13920 48217 13923
rect 48096 13892 48217 13920
rect 48096 13880 48102 13892
rect 48205 13889 48217 13892
rect 48251 13889 48263 13923
rect 48205 13883 48263 13889
rect 48958 13880 48964 13932
rect 49016 13920 49022 13932
rect 50045 13923 50103 13929
rect 50045 13920 50057 13923
rect 49016 13892 50057 13920
rect 49016 13880 49022 13892
rect 50045 13889 50057 13892
rect 50091 13889 50103 13923
rect 50172 13920 50200 13948
rect 51442 13920 51448 13932
rect 50172 13892 51448 13920
rect 50045 13883 50103 13889
rect 51442 13880 51448 13892
rect 51500 13880 51506 13932
rect 51718 13880 51724 13932
rect 51776 13920 51782 13932
rect 52932 13929 52960 13960
rect 54570 13948 54576 13960
rect 54628 13988 54634 14000
rect 55582 13988 55588 14000
rect 54628 13960 55588 13988
rect 54628 13948 54634 13960
rect 55582 13948 55588 13960
rect 55640 13948 55646 14000
rect 56226 13948 56232 14000
rect 56284 13988 56290 14000
rect 57425 13991 57483 13997
rect 57425 13988 57437 13991
rect 56284 13960 57437 13988
rect 56284 13948 56290 13960
rect 57425 13957 57437 13960
rect 57471 13957 57483 13991
rect 57532 13988 57560 14028
rect 57983 14025 57995 14059
rect 58029 14056 58041 14059
rect 60550 14056 60556 14068
rect 58029 14028 60556 14056
rect 58029 14025 58041 14028
rect 57983 14019 58041 14025
rect 60550 14016 60556 14028
rect 60608 14016 60614 14068
rect 61562 14016 61568 14068
rect 61620 14056 61626 14068
rect 64233 14059 64291 14065
rect 61620 14028 63724 14056
rect 61620 14016 61626 14028
rect 61746 13988 61752 14000
rect 57532 13960 61752 13988
rect 57425 13951 57483 13957
rect 61746 13948 61752 13960
rect 61804 13948 61810 14000
rect 61938 13991 61996 13997
rect 61938 13957 61950 13991
rect 61984 13988 61996 13991
rect 62298 13988 62304 14000
rect 61984 13960 62304 13988
rect 61984 13957 61996 13960
rect 61938 13951 61996 13957
rect 62298 13948 62304 13960
rect 62356 13948 62362 14000
rect 63034 13988 63040 14000
rect 62995 13960 63040 13988
rect 63034 13948 63040 13960
rect 63092 13948 63098 14000
rect 63405 13991 63463 13997
rect 63405 13957 63417 13991
rect 63451 13988 63463 13991
rect 63586 13988 63592 14000
rect 63451 13960 63592 13988
rect 63451 13957 63463 13960
rect 63405 13951 63463 13957
rect 63586 13948 63592 13960
rect 63644 13948 63650 14000
rect 63696 13988 63724 14028
rect 64233 14025 64245 14059
rect 64279 14056 64291 14059
rect 64506 14056 64512 14068
rect 64279 14028 64512 14056
rect 64279 14025 64291 14028
rect 64233 14019 64291 14025
rect 64506 14016 64512 14028
rect 64564 14016 64570 14068
rect 64874 14016 64880 14068
rect 64932 14056 64938 14068
rect 65061 14059 65119 14065
rect 65061 14056 65073 14059
rect 64932 14028 65073 14056
rect 64932 14016 64938 14028
rect 65061 14025 65073 14028
rect 65107 14025 65119 14059
rect 65061 14019 65119 14025
rect 67545 14059 67603 14065
rect 67545 14025 67557 14059
rect 67591 14056 67603 14059
rect 67726 14056 67732 14068
rect 67591 14028 67732 14056
rect 67591 14025 67603 14028
rect 67545 14019 67603 14025
rect 67726 14016 67732 14028
rect 67784 14016 67790 14068
rect 68002 14016 68008 14068
rect 68060 14056 68066 14068
rect 69474 14056 69480 14068
rect 68060 14028 69480 14056
rect 68060 14016 68066 14028
rect 67450 13988 67456 14000
rect 63696 13960 67456 13988
rect 67450 13948 67456 13960
rect 67508 13948 67514 14000
rect 68388 13988 68416 14028
rect 69474 14016 69480 14028
rect 69532 14016 69538 14068
rect 70210 14016 70216 14068
rect 70268 14056 70274 14068
rect 70765 14059 70823 14065
rect 70765 14056 70777 14059
rect 70268 14028 70777 14056
rect 70268 14016 70274 14028
rect 70765 14025 70777 14028
rect 70811 14025 70823 14059
rect 70765 14019 70823 14025
rect 71774 14016 71780 14068
rect 71832 14056 71838 14068
rect 72421 14059 72479 14065
rect 72421 14056 72433 14059
rect 71832 14028 72433 14056
rect 71832 14016 71838 14028
rect 72421 14025 72433 14028
rect 72467 14025 72479 14059
rect 73890 14056 73896 14068
rect 73851 14028 73896 14056
rect 72421 14019 72479 14025
rect 73890 14016 73896 14028
rect 73948 14016 73954 14068
rect 80026 14028 84194 14056
rect 68388 13960 68508 13988
rect 67729 13932 67787 13933
rect 52917 13923 52975 13929
rect 51776 13892 51821 13920
rect 51776 13880 51782 13892
rect 52917 13889 52929 13923
rect 52963 13889 52975 13923
rect 52917 13883 52975 13889
rect 53184 13923 53242 13929
rect 53184 13889 53196 13923
rect 53230 13920 53242 13923
rect 55030 13920 55036 13932
rect 53230 13892 55036 13920
rect 53230 13889 53242 13892
rect 53184 13883 53242 13889
rect 55030 13880 55036 13892
rect 55088 13880 55094 13932
rect 55125 13923 55183 13929
rect 55125 13889 55137 13923
rect 55171 13920 55183 13923
rect 56778 13920 56784 13932
rect 55171 13892 56784 13920
rect 55171 13889 55183 13892
rect 55125 13883 55183 13889
rect 45557 13855 45615 13861
rect 45557 13821 45569 13855
rect 45603 13821 45615 13855
rect 45922 13852 45928 13864
rect 45883 13824 45928 13852
rect 45557 13815 45615 13821
rect 45572 13784 45600 13815
rect 45922 13812 45928 13824
rect 45980 13812 45986 13864
rect 46750 13812 46756 13864
rect 46808 13852 46814 13864
rect 47949 13855 48007 13861
rect 47949 13852 47961 13855
rect 46808 13824 47961 13852
rect 46808 13812 46814 13824
rect 47949 13821 47961 13824
rect 47995 13821 48007 13855
rect 49786 13852 49792 13864
rect 49747 13824 49792 13852
rect 47949 13815 48007 13821
rect 49786 13812 49792 13824
rect 49844 13812 49850 13864
rect 51534 13852 51540 13864
rect 51495 13824 51540 13852
rect 51534 13812 51540 13824
rect 51592 13812 51598 13864
rect 51905 13855 51963 13861
rect 51905 13821 51917 13855
rect 51951 13852 51963 13855
rect 51994 13852 52000 13864
rect 51951 13824 52000 13852
rect 51951 13821 51963 13824
rect 51905 13815 51963 13821
rect 51994 13812 52000 13824
rect 52052 13812 52058 13864
rect 54110 13812 54116 13864
rect 54168 13852 54174 13864
rect 55140 13852 55168 13883
rect 56778 13880 56784 13892
rect 56836 13880 56842 13932
rect 56870 13880 56876 13932
rect 56928 13920 56934 13932
rect 57057 13923 57115 13929
rect 57057 13920 57069 13923
rect 56928 13892 57069 13920
rect 56928 13880 56934 13892
rect 57057 13889 57069 13892
rect 57103 13889 57115 13923
rect 57238 13920 57244 13932
rect 57199 13892 57244 13920
rect 57057 13883 57115 13889
rect 57238 13880 57244 13892
rect 57296 13880 57302 13932
rect 57882 13920 57888 13932
rect 57843 13892 57888 13920
rect 57882 13880 57888 13892
rect 57940 13880 57946 13932
rect 58069 13923 58127 13929
rect 58069 13889 58081 13923
rect 58115 13889 58127 13923
rect 58069 13883 58127 13889
rect 58170 13926 58228 13929
rect 58342 13926 58348 13932
rect 58170 13923 58348 13926
rect 58170 13889 58182 13923
rect 58216 13898 58348 13923
rect 58216 13889 58228 13898
rect 58170 13883 58228 13889
rect 54168 13824 55168 13852
rect 54168 13812 54174 13824
rect 55214 13812 55220 13864
rect 55272 13852 55278 13864
rect 55309 13855 55367 13861
rect 55309 13852 55321 13855
rect 55272 13824 55321 13852
rect 55272 13812 55278 13824
rect 55309 13821 55321 13824
rect 55355 13821 55367 13855
rect 55674 13852 55680 13864
rect 55635 13824 55680 13852
rect 55309 13815 55367 13821
rect 55674 13812 55680 13824
rect 55732 13812 55738 13864
rect 55953 13855 56011 13861
rect 55953 13821 55965 13855
rect 55999 13852 56011 13855
rect 56962 13852 56968 13864
rect 55999 13824 56968 13852
rect 55999 13821 56011 13824
rect 55953 13815 56011 13821
rect 56962 13812 56968 13824
rect 57020 13812 57026 13864
rect 57330 13812 57336 13864
rect 57388 13852 57394 13864
rect 58084 13852 58112 13883
rect 58342 13880 58348 13898
rect 58400 13880 58406 13932
rect 59081 13923 59139 13929
rect 58452 13892 58940 13920
rect 58452 13852 58480 13892
rect 57388 13824 58480 13852
rect 57388 13812 57394 13824
rect 58526 13812 58532 13864
rect 58584 13852 58590 13864
rect 58805 13855 58863 13861
rect 58805 13852 58817 13855
rect 58584 13824 58817 13852
rect 58584 13812 58590 13824
rect 58805 13821 58817 13824
rect 58851 13821 58863 13855
rect 58912 13852 58940 13892
rect 59081 13889 59093 13923
rect 59127 13920 59139 13923
rect 59446 13920 59452 13932
rect 59127 13892 59452 13920
rect 59127 13889 59139 13892
rect 59081 13883 59139 13889
rect 59446 13880 59452 13892
rect 59504 13880 59510 13932
rect 61657 13923 61715 13929
rect 61657 13889 61669 13923
rect 61703 13889 61715 13923
rect 61838 13920 61844 13932
rect 61799 13892 61844 13920
rect 61657 13883 61715 13889
rect 59170 13852 59176 13864
rect 58912 13824 59176 13852
rect 58805 13815 58863 13821
rect 59170 13812 59176 13824
rect 59228 13812 59234 13864
rect 59262 13812 59268 13864
rect 59320 13852 59326 13864
rect 60461 13855 60519 13861
rect 60461 13852 60473 13855
rect 59320 13824 60473 13852
rect 59320 13812 59326 13824
rect 60461 13821 60473 13824
rect 60507 13852 60519 13855
rect 60642 13852 60648 13864
rect 60507 13824 60648 13852
rect 60507 13821 60519 13824
rect 60461 13815 60519 13821
rect 60642 13812 60648 13824
rect 60700 13812 60706 13864
rect 60737 13855 60795 13861
rect 60737 13821 60749 13855
rect 60783 13852 60795 13855
rect 61010 13852 61016 13864
rect 60783 13824 61016 13852
rect 60783 13821 60795 13824
rect 60737 13815 60795 13821
rect 61010 13812 61016 13824
rect 61068 13812 61074 13864
rect 61672 13852 61700 13883
rect 61838 13880 61844 13892
rect 61896 13880 61902 13932
rect 62022 13880 62028 13932
rect 62080 13929 62086 13932
rect 62080 13920 62088 13929
rect 62482 13920 62488 13932
rect 62080 13892 62488 13920
rect 62080 13883 62088 13892
rect 62080 13880 62086 13883
rect 62482 13880 62488 13892
rect 62540 13880 62546 13932
rect 63218 13920 63224 13932
rect 63179 13892 63224 13920
rect 63218 13880 63224 13892
rect 63276 13880 63282 13932
rect 63494 13920 63500 13932
rect 63455 13892 63500 13920
rect 63494 13880 63500 13892
rect 63552 13880 63558 13932
rect 64046 13920 64052 13932
rect 64007 13892 64052 13920
rect 64046 13880 64052 13892
rect 64104 13880 64110 13932
rect 64325 13923 64383 13929
rect 64325 13889 64337 13923
rect 64371 13889 64383 13923
rect 64325 13883 64383 13889
rect 62574 13852 62580 13864
rect 61672 13824 62580 13852
rect 62574 13812 62580 13824
rect 62632 13812 62638 13864
rect 63954 13812 63960 13864
rect 64012 13852 64018 13864
rect 64340 13852 64368 13883
rect 64598 13880 64604 13932
rect 64656 13918 64662 13932
rect 64785 13923 64843 13929
rect 64785 13918 64797 13923
rect 64656 13890 64797 13918
rect 64656 13880 64662 13890
rect 64785 13889 64797 13890
rect 64831 13889 64843 13923
rect 64785 13883 64843 13889
rect 64877 13923 64935 13929
rect 64877 13889 64889 13923
rect 64923 13920 64935 13923
rect 64966 13920 64972 13932
rect 64923 13892 64972 13920
rect 64923 13889 64935 13892
rect 64877 13883 64935 13889
rect 64966 13880 64972 13892
rect 65024 13880 65030 13932
rect 65150 13880 65156 13932
rect 65208 13920 65214 13932
rect 65208 13892 66254 13920
rect 65208 13880 65214 13892
rect 64012 13824 64368 13852
rect 66226 13852 66254 13892
rect 67726 13880 67732 13932
rect 67784 13920 67790 13932
rect 68370 13920 68376 13932
rect 67784 13892 67825 13920
rect 68189 13913 68247 13919
rect 67784 13880 67790 13892
rect 68189 13879 68201 13913
rect 68235 13879 68247 13913
rect 68331 13892 68376 13920
rect 68370 13880 68376 13892
rect 68428 13880 68434 13932
rect 68480 13929 68508 13960
rect 69106 13948 69112 14000
rect 69164 13988 69170 14000
rect 80026 13988 80054 14028
rect 69164 13960 80054 13988
rect 69164 13948 69170 13960
rect 68558 13929 68616 13935
rect 68465 13923 68523 13929
rect 68465 13889 68477 13923
rect 68511 13889 68523 13923
rect 68558 13895 68570 13929
rect 68604 13926 68616 13929
rect 68646 13926 68652 13932
rect 68604 13898 68652 13926
rect 68604 13895 68616 13898
rect 68558 13889 68616 13895
rect 68465 13883 68523 13889
rect 68646 13880 68652 13898
rect 68704 13880 68710 13932
rect 68922 13880 68928 13932
rect 68980 13920 68986 13932
rect 69641 13923 69699 13929
rect 69641 13920 69653 13923
rect 68980 13892 69653 13920
rect 68980 13880 68986 13892
rect 69641 13889 69653 13892
rect 69687 13889 69699 13923
rect 69641 13883 69699 13889
rect 70118 13880 70124 13932
rect 70176 13920 70182 13932
rect 71317 13923 71375 13929
rect 71317 13920 71329 13923
rect 70176 13892 71329 13920
rect 70176 13880 70182 13892
rect 71317 13889 71329 13892
rect 71363 13920 71375 13923
rect 71866 13920 71872 13932
rect 71363 13892 71872 13920
rect 71363 13889 71375 13892
rect 71317 13883 71375 13889
rect 71866 13880 71872 13892
rect 71924 13880 71930 13932
rect 71958 13880 71964 13932
rect 72016 13920 72022 13932
rect 72053 13923 72111 13929
rect 72053 13920 72065 13923
rect 72016 13892 72065 13920
rect 72016 13880 72022 13892
rect 72053 13889 72065 13892
rect 72099 13889 72111 13923
rect 72234 13920 72240 13932
rect 72195 13892 72240 13920
rect 72053 13883 72111 13889
rect 72234 13880 72240 13892
rect 72292 13880 72298 13932
rect 72326 13880 72332 13932
rect 72384 13920 72390 13932
rect 72513 13923 72571 13929
rect 72513 13920 72525 13923
rect 72384 13892 72525 13920
rect 72384 13880 72390 13892
rect 72513 13889 72525 13892
rect 72559 13889 72571 13923
rect 73706 13920 73712 13932
rect 73667 13892 73712 13920
rect 72513 13883 72571 13889
rect 73706 13880 73712 13892
rect 73764 13880 73770 13932
rect 84166 13920 84194 14028
rect 88245 13923 88303 13929
rect 88245 13920 88257 13923
rect 84166 13892 88257 13920
rect 88245 13889 88257 13892
rect 88291 13889 88303 13923
rect 88245 13883 88303 13889
rect 68189 13873 68247 13879
rect 68002 13852 68008 13864
rect 66226 13824 68008 13852
rect 64012 13812 64018 13824
rect 68002 13812 68008 13824
rect 68060 13812 68066 13864
rect 68204 13796 68232 13873
rect 69014 13812 69020 13864
rect 69072 13852 69078 13864
rect 69382 13852 69388 13864
rect 69072 13824 69388 13852
rect 69072 13812 69078 13824
rect 69382 13812 69388 13824
rect 69440 13812 69446 13864
rect 71222 13852 71228 13864
rect 71148 13824 71228 13852
rect 45572 13756 47992 13784
rect 47964 13728 47992 13756
rect 49050 13744 49056 13796
rect 49108 13784 49114 13796
rect 49329 13787 49387 13793
rect 49329 13784 49341 13787
rect 49108 13756 49341 13784
rect 49108 13744 49114 13756
rect 49329 13753 49341 13756
rect 49375 13784 49387 13787
rect 49510 13784 49516 13796
rect 49375 13756 49516 13784
rect 49375 13753 49387 13756
rect 49329 13747 49387 13753
rect 49510 13744 49516 13756
rect 49568 13744 49574 13796
rect 51350 13744 51356 13796
rect 51408 13784 51414 13796
rect 52914 13784 52920 13796
rect 51408 13756 52920 13784
rect 51408 13744 51414 13756
rect 52914 13744 52920 13756
rect 52972 13744 52978 13796
rect 53852 13756 66254 13784
rect 45830 13716 45836 13728
rect 45480 13688 45836 13716
rect 45189 13679 45247 13685
rect 45830 13676 45836 13688
rect 45888 13676 45894 13728
rect 47026 13716 47032 13728
rect 46987 13688 47032 13716
rect 47026 13676 47032 13688
rect 47084 13676 47090 13728
rect 47946 13676 47952 13728
rect 48004 13716 48010 13728
rect 50154 13716 50160 13728
rect 48004 13688 50160 13716
rect 48004 13676 48010 13688
rect 50154 13676 50160 13688
rect 50212 13676 50218 13728
rect 50430 13676 50436 13728
rect 50488 13716 50494 13728
rect 53852 13716 53880 13756
rect 50488 13688 53880 13716
rect 54297 13719 54355 13725
rect 50488 13676 50494 13688
rect 54297 13685 54309 13719
rect 54343 13716 54355 13719
rect 54386 13716 54392 13728
rect 54343 13688 54392 13716
rect 54343 13685 54355 13688
rect 54297 13679 54355 13685
rect 54386 13676 54392 13688
rect 54444 13716 54450 13728
rect 54662 13716 54668 13728
rect 54444 13688 54668 13716
rect 54444 13676 54450 13688
rect 54662 13676 54668 13688
rect 54720 13676 54726 13728
rect 54938 13676 54944 13728
rect 54996 13716 55002 13728
rect 62114 13716 62120 13728
rect 54996 13688 62120 13716
rect 54996 13676 55002 13688
rect 62114 13676 62120 13688
rect 62172 13676 62178 13728
rect 62209 13719 62267 13725
rect 62209 13685 62221 13719
rect 62255 13716 62267 13719
rect 62390 13716 62396 13728
rect 62255 13688 62396 13716
rect 62255 13685 62267 13688
rect 62209 13679 62267 13685
rect 62390 13676 62396 13688
rect 62448 13676 62454 13728
rect 63862 13716 63868 13728
rect 63823 13688 63868 13716
rect 63862 13676 63868 13688
rect 63920 13676 63926 13728
rect 66226 13716 66254 13756
rect 68186 13744 68192 13796
rect 68244 13744 68250 13796
rect 68833 13787 68891 13793
rect 68833 13753 68845 13787
rect 68879 13753 68891 13787
rect 68833 13747 68891 13753
rect 68848 13716 68876 13747
rect 70578 13744 70584 13796
rect 70636 13784 70642 13796
rect 71148 13784 71176 13824
rect 71222 13812 71228 13824
rect 71280 13852 71286 13864
rect 73525 13855 73583 13861
rect 73525 13852 73537 13855
rect 71280 13824 71373 13852
rect 71516 13824 73537 13852
rect 71280 13812 71286 13824
rect 70636 13756 71176 13784
rect 70636 13744 70642 13756
rect 71314 13744 71320 13796
rect 71372 13784 71378 13796
rect 71516 13784 71544 13824
rect 73525 13821 73537 13824
rect 73571 13821 73583 13855
rect 73525 13815 73583 13821
rect 71372 13756 71544 13784
rect 71372 13744 71378 13756
rect 66226 13688 68876 13716
rect 71038 13676 71044 13728
rect 71096 13716 71102 13728
rect 71685 13719 71743 13725
rect 71685 13716 71697 13719
rect 71096 13688 71697 13716
rect 71096 13676 71102 13688
rect 71685 13685 71697 13688
rect 71731 13685 71743 13719
rect 88058 13716 88064 13728
rect 88019 13688 88064 13716
rect 71685 13679 71743 13685
rect 88058 13676 88064 13688
rect 88116 13676 88122 13728
rect 1104 13626 88872 13648
rect 1104 13574 11924 13626
rect 11976 13574 11988 13626
rect 12040 13574 12052 13626
rect 12104 13574 12116 13626
rect 12168 13574 12180 13626
rect 12232 13574 33872 13626
rect 33924 13574 33936 13626
rect 33988 13574 34000 13626
rect 34052 13574 34064 13626
rect 34116 13574 34128 13626
rect 34180 13574 55820 13626
rect 55872 13574 55884 13626
rect 55936 13574 55948 13626
rect 56000 13574 56012 13626
rect 56064 13574 56076 13626
rect 56128 13574 77768 13626
rect 77820 13574 77832 13626
rect 77884 13574 77896 13626
rect 77948 13574 77960 13626
rect 78012 13574 78024 13626
rect 78076 13574 88872 13626
rect 1104 13552 88872 13574
rect 19058 13472 19064 13524
rect 19116 13512 19122 13524
rect 19978 13512 19984 13524
rect 19116 13484 19984 13512
rect 19116 13472 19122 13484
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 20806 13472 20812 13524
rect 20864 13512 20870 13524
rect 20901 13515 20959 13521
rect 20901 13512 20913 13515
rect 20864 13484 20913 13512
rect 20864 13472 20870 13484
rect 20901 13481 20913 13484
rect 20947 13481 20959 13515
rect 21818 13512 21824 13524
rect 20901 13475 20959 13481
rect 21284 13484 21824 13512
rect 19705 13447 19763 13453
rect 19705 13413 19717 13447
rect 19751 13413 19763 13447
rect 19886 13444 19892 13456
rect 19847 13416 19892 13444
rect 19705 13407 19763 13413
rect 19610 13376 19616 13388
rect 19571 13348 19616 13376
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 19720 13376 19748 13407
rect 19886 13404 19892 13416
rect 19944 13404 19950 13456
rect 20162 13404 20168 13456
rect 20220 13444 20226 13456
rect 21284 13444 21312 13484
rect 21818 13472 21824 13484
rect 21876 13512 21882 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 21876 13484 22109 13512
rect 21876 13472 21882 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 22554 13472 22560 13524
rect 22612 13512 22618 13524
rect 22925 13515 22983 13521
rect 22925 13512 22937 13515
rect 22612 13484 22937 13512
rect 22612 13472 22618 13484
rect 22925 13481 22937 13484
rect 22971 13481 22983 13515
rect 23290 13512 23296 13524
rect 23251 13484 23296 13512
rect 22925 13475 22983 13481
rect 23290 13472 23296 13484
rect 23348 13472 23354 13524
rect 23845 13515 23903 13521
rect 23845 13481 23857 13515
rect 23891 13512 23903 13515
rect 24762 13512 24768 13524
rect 23891 13484 24768 13512
rect 23891 13481 23903 13484
rect 23845 13475 23903 13481
rect 24762 13472 24768 13484
rect 24820 13472 24826 13524
rect 25685 13515 25743 13521
rect 25685 13481 25697 13515
rect 25731 13481 25743 13515
rect 25685 13475 25743 13481
rect 20220 13416 21312 13444
rect 21361 13447 21419 13453
rect 20220 13404 20226 13416
rect 21361 13413 21373 13447
rect 21407 13413 21419 13447
rect 25700 13444 25728 13475
rect 26050 13472 26056 13524
rect 26108 13512 26114 13524
rect 27522 13512 27528 13524
rect 26108 13484 27528 13512
rect 26108 13472 26114 13484
rect 27522 13472 27528 13484
rect 27580 13472 27586 13524
rect 28258 13472 28264 13524
rect 28316 13512 28322 13524
rect 28721 13515 28779 13521
rect 28721 13512 28733 13515
rect 28316 13484 28733 13512
rect 28316 13472 28322 13484
rect 28721 13481 28733 13484
rect 28767 13481 28779 13515
rect 28721 13475 28779 13481
rect 28994 13472 29000 13524
rect 29052 13512 29058 13524
rect 30282 13512 30288 13524
rect 29052 13484 30288 13512
rect 29052 13472 29058 13484
rect 30282 13472 30288 13484
rect 30340 13472 30346 13524
rect 30466 13472 30472 13524
rect 30524 13512 30530 13524
rect 31938 13512 31944 13524
rect 30524 13484 31944 13512
rect 30524 13472 30530 13484
rect 31938 13472 31944 13484
rect 31996 13512 32002 13524
rect 34606 13512 34612 13524
rect 31996 13484 34612 13512
rect 31996 13472 32002 13484
rect 34606 13472 34612 13484
rect 34664 13472 34670 13524
rect 37182 13472 37188 13524
rect 37240 13512 37246 13524
rect 37737 13515 37795 13521
rect 37737 13512 37749 13515
rect 37240 13484 37749 13512
rect 37240 13472 37246 13484
rect 37737 13481 37749 13484
rect 37783 13481 37795 13515
rect 37737 13475 37795 13481
rect 38838 13472 38844 13524
rect 38896 13512 38902 13524
rect 38933 13515 38991 13521
rect 38933 13512 38945 13515
rect 38896 13484 38945 13512
rect 38896 13472 38902 13484
rect 38933 13481 38945 13484
rect 38979 13481 38991 13515
rect 41782 13512 41788 13524
rect 38933 13475 38991 13481
rect 39132 13484 41788 13512
rect 21361 13407 21419 13413
rect 22388 13416 25728 13444
rect 20993 13379 21051 13385
rect 20993 13376 21005 13379
rect 19720 13348 21005 13376
rect 20993 13345 21005 13348
rect 21039 13345 21051 13379
rect 21376 13376 21404 13407
rect 22388 13376 22416 13416
rect 25866 13404 25872 13456
rect 25924 13444 25930 13456
rect 27890 13444 27896 13456
rect 25924 13416 27752 13444
rect 27851 13416 27896 13444
rect 25924 13404 25930 13416
rect 21376 13348 22416 13376
rect 22465 13379 22523 13385
rect 20993 13339 21051 13345
rect 22465 13345 22477 13379
rect 22511 13376 22523 13379
rect 23658 13376 23664 13388
rect 22511 13348 23664 13376
rect 22511 13345 22523 13348
rect 22465 13339 22523 13345
rect 23658 13336 23664 13348
rect 23716 13336 23722 13388
rect 24578 13376 24584 13388
rect 24491 13348 24584 13376
rect 24578 13336 24584 13348
rect 24636 13376 24642 13388
rect 25498 13376 25504 13388
rect 24636 13348 25504 13376
rect 24636 13336 24642 13348
rect 25498 13336 25504 13348
rect 25556 13336 25562 13388
rect 25682 13376 25688 13388
rect 25643 13348 25688 13376
rect 25682 13336 25688 13348
rect 25740 13336 25746 13388
rect 26418 13336 26424 13388
rect 26476 13376 26482 13388
rect 26476 13348 26832 13376
rect 26476 13336 26482 13348
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 6886 13280 15025 13308
rect 1397 13175 1455 13181
rect 1397 13141 1409 13175
rect 1443 13172 1455 13175
rect 6886 13172 6914 13280
rect 15013 13277 15025 13280
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13277 18015 13311
rect 18230 13308 18236 13320
rect 18191 13280 18236 13308
rect 17957 13271 18015 13277
rect 17972 13240 18000 13271
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 19058 13268 19064 13320
rect 19116 13308 19122 13320
rect 19521 13311 19579 13317
rect 19521 13308 19533 13311
rect 19116 13280 19533 13308
rect 19116 13268 19122 13280
rect 19521 13277 19533 13280
rect 19567 13277 19579 13311
rect 19702 13308 19708 13320
rect 19663 13280 19708 13308
rect 19521 13271 19579 13277
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 19978 13308 19984 13320
rect 19939 13280 19984 13308
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20070 13268 20076 13320
rect 20128 13308 20134 13320
rect 20714 13308 20720 13320
rect 20128 13280 20720 13308
rect 20128 13268 20134 13280
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 21082 13268 21088 13320
rect 21140 13308 21146 13320
rect 21177 13311 21235 13317
rect 21177 13308 21189 13311
rect 21140 13280 21189 13308
rect 21140 13268 21146 13280
rect 21177 13277 21189 13280
rect 21223 13277 21235 13311
rect 22002 13308 22008 13320
rect 21963 13280 22008 13308
rect 21177 13271 21235 13277
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 22370 13268 22376 13320
rect 22428 13308 22434 13320
rect 22554 13308 22560 13320
rect 22428 13280 22560 13308
rect 22428 13268 22434 13280
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 22833 13311 22891 13317
rect 22833 13277 22845 13311
rect 22879 13308 22891 13311
rect 23753 13311 23811 13317
rect 23753 13308 23765 13311
rect 22879 13280 23765 13308
rect 22879 13277 22891 13280
rect 22833 13271 22891 13277
rect 23753 13277 23765 13280
rect 23799 13308 23811 13311
rect 24118 13308 24124 13320
rect 23799 13280 24124 13308
rect 23799 13277 23811 13280
rect 23753 13271 23811 13277
rect 24118 13268 24124 13280
rect 24176 13268 24182 13320
rect 24210 13268 24216 13320
rect 24268 13308 24274 13320
rect 24489 13311 24547 13317
rect 24489 13308 24501 13311
rect 24268 13280 24501 13308
rect 24268 13268 24274 13280
rect 24489 13277 24501 13280
rect 24535 13277 24547 13311
rect 25038 13308 25044 13320
rect 24999 13280 25044 13308
rect 24489 13271 24547 13277
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 25406 13268 25412 13320
rect 25464 13308 25470 13320
rect 25869 13311 25927 13317
rect 25869 13308 25881 13311
rect 25464 13280 25881 13308
rect 25464 13268 25470 13280
rect 25869 13277 25881 13280
rect 25915 13277 25927 13311
rect 26510 13308 26516 13320
rect 26471 13280 26516 13308
rect 25869 13271 25927 13277
rect 26510 13268 26516 13280
rect 26568 13268 26574 13320
rect 26602 13268 26608 13320
rect 26660 13308 26666 13320
rect 26804 13317 26832 13348
rect 26896 13348 27568 13376
rect 26896 13317 26924 13348
rect 27540 13320 27568 13348
rect 26789 13311 26847 13317
rect 26660 13280 26705 13308
rect 26660 13268 26666 13280
rect 26789 13277 26801 13311
rect 26835 13277 26847 13311
rect 26789 13271 26847 13277
rect 26881 13311 26939 13317
rect 26881 13277 26893 13311
rect 26927 13277 26939 13311
rect 26881 13271 26939 13277
rect 26978 13311 27036 13317
rect 26978 13277 26990 13311
rect 27024 13277 27036 13311
rect 27522 13308 27528 13320
rect 27483 13280 27528 13308
rect 26978 13271 27036 13277
rect 20438 13240 20444 13252
rect 17972 13212 20444 13240
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 20901 13243 20959 13249
rect 20901 13209 20913 13243
rect 20947 13240 20959 13243
rect 23566 13240 23572 13252
rect 20947 13212 23572 13240
rect 20947 13209 20959 13212
rect 20901 13203 20959 13209
rect 23566 13200 23572 13212
rect 23624 13200 23630 13252
rect 23658 13200 23664 13252
rect 23716 13240 23722 13252
rect 23934 13240 23940 13252
rect 23716 13212 23940 13240
rect 23716 13200 23722 13212
rect 23934 13200 23940 13212
rect 23992 13200 23998 13252
rect 25593 13243 25651 13249
rect 25593 13240 25605 13243
rect 24044 13212 25605 13240
rect 1443 13144 6914 13172
rect 15105 13175 15163 13181
rect 1443 13141 1455 13144
rect 1397 13135 1455 13141
rect 15105 13141 15117 13175
rect 15151 13172 15163 13175
rect 20714 13172 20720 13184
rect 15151 13144 20720 13172
rect 15151 13141 15163 13144
rect 15105 13135 15163 13141
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 22462 13132 22468 13184
rect 22520 13172 22526 13184
rect 24044 13172 24072 13212
rect 25593 13209 25605 13212
rect 25639 13209 25651 13243
rect 26988 13240 27016 13271
rect 27522 13268 27528 13280
rect 27580 13268 27586 13320
rect 25593 13203 25651 13209
rect 25976 13212 27016 13240
rect 27724 13240 27752 13416
rect 27890 13404 27896 13416
rect 27948 13404 27954 13456
rect 28442 13404 28448 13456
rect 28500 13444 28506 13456
rect 28500 13416 32536 13444
rect 28500 13404 28506 13416
rect 29178 13376 29184 13388
rect 28644 13348 29184 13376
rect 28644 13317 28672 13348
rect 29178 13336 29184 13348
rect 29236 13336 29242 13388
rect 30926 13336 30932 13388
rect 30984 13376 30990 13388
rect 31294 13376 31300 13388
rect 30984 13348 31300 13376
rect 30984 13336 30990 13348
rect 31294 13336 31300 13348
rect 31352 13336 31358 13388
rect 31846 13376 31852 13388
rect 31807 13348 31852 13376
rect 31846 13336 31852 13348
rect 31904 13336 31910 13388
rect 32508 13376 32536 13416
rect 32582 13404 32588 13456
rect 32640 13444 32646 13456
rect 32950 13444 32956 13456
rect 32640 13416 32956 13444
rect 32640 13404 32646 13416
rect 32950 13404 32956 13416
rect 33008 13404 33014 13456
rect 33042 13404 33048 13456
rect 33100 13444 33106 13456
rect 33100 13416 34744 13444
rect 33100 13404 33106 13416
rect 32766 13376 32772 13388
rect 32508 13348 32772 13376
rect 32766 13336 32772 13348
rect 32824 13336 32830 13388
rect 34606 13376 34612 13388
rect 33040 13348 34612 13376
rect 28629 13311 28687 13317
rect 28629 13277 28641 13311
rect 28675 13277 28687 13311
rect 28629 13271 28687 13277
rect 29549 13311 29607 13317
rect 29549 13277 29561 13311
rect 29595 13308 29607 13311
rect 29595 13280 30052 13308
rect 29595 13277 29607 13280
rect 29549 13271 29607 13277
rect 29178 13240 29184 13252
rect 27724 13212 29184 13240
rect 22520 13144 24072 13172
rect 25133 13175 25191 13181
rect 22520 13132 22526 13144
rect 25133 13141 25145 13175
rect 25179 13172 25191 13175
rect 25976 13172 26004 13212
rect 29178 13200 29184 13212
rect 29236 13200 29242 13252
rect 29638 13240 29644 13252
rect 29599 13212 29644 13240
rect 29638 13200 29644 13212
rect 29696 13200 29702 13252
rect 30024 13240 30052 13280
rect 30098 13268 30104 13320
rect 30156 13308 30162 13320
rect 30834 13308 30840 13320
rect 30156 13280 30201 13308
rect 30795 13280 30840 13308
rect 30156 13268 30162 13280
rect 30834 13268 30840 13280
rect 30892 13268 30898 13320
rect 31573 13311 31631 13317
rect 31573 13277 31585 13311
rect 31619 13308 31631 13311
rect 31662 13308 31668 13320
rect 31619 13280 31668 13308
rect 31619 13277 31631 13280
rect 31573 13271 31631 13277
rect 31662 13268 31668 13280
rect 31720 13268 31726 13320
rect 32306 13268 32312 13320
rect 32364 13308 32370 13320
rect 32953 13311 33011 13317
rect 32953 13308 32965 13311
rect 32364 13280 32965 13308
rect 32364 13268 32370 13280
rect 32953 13277 32965 13280
rect 32999 13308 33011 13311
rect 33040 13308 33068 13348
rect 34606 13336 34612 13348
rect 34664 13336 34670 13388
rect 34716 13385 34744 13416
rect 35710 13404 35716 13456
rect 35768 13444 35774 13456
rect 38654 13444 38660 13456
rect 35768 13416 38660 13444
rect 35768 13404 35774 13416
rect 38654 13404 38660 13416
rect 38712 13404 38718 13456
rect 34701 13379 34759 13385
rect 34701 13345 34713 13379
rect 34747 13345 34759 13379
rect 34701 13339 34759 13345
rect 36814 13336 36820 13388
rect 36872 13376 36878 13388
rect 38746 13376 38752 13388
rect 36872 13348 38752 13376
rect 36872 13336 36878 13348
rect 38746 13336 38752 13348
rect 38804 13336 38810 13388
rect 32999 13280 33068 13308
rect 33505 13311 33563 13317
rect 32999 13277 33011 13280
rect 32953 13271 33011 13277
rect 33505 13277 33517 13311
rect 33551 13308 33563 13311
rect 33778 13308 33784 13320
rect 33551 13280 33784 13308
rect 33551 13277 33563 13280
rect 33505 13271 33563 13277
rect 33778 13268 33784 13280
rect 33836 13308 33842 13320
rect 33873 13311 33931 13317
rect 33873 13308 33885 13311
rect 33836 13280 33885 13308
rect 33836 13268 33842 13280
rect 33873 13277 33885 13280
rect 33919 13308 33931 13311
rect 34146 13308 34152 13320
rect 33919 13280 34152 13308
rect 33919 13277 33931 13280
rect 33873 13271 33931 13277
rect 34146 13268 34152 13280
rect 34204 13268 34210 13320
rect 34790 13268 34796 13320
rect 34848 13308 34854 13320
rect 39132 13317 39160 13484
rect 41782 13472 41788 13484
rect 41840 13472 41846 13524
rect 42426 13472 42432 13524
rect 42484 13512 42490 13524
rect 42978 13512 42984 13524
rect 42484 13484 42984 13512
rect 42484 13472 42490 13484
rect 42978 13472 42984 13484
rect 43036 13472 43042 13524
rect 43622 13512 43628 13524
rect 43583 13484 43628 13512
rect 43622 13472 43628 13484
rect 43680 13472 43686 13524
rect 44358 13512 44364 13524
rect 44319 13484 44364 13512
rect 44358 13472 44364 13484
rect 44416 13472 44422 13524
rect 44450 13472 44456 13524
rect 44508 13512 44514 13524
rect 44634 13512 44640 13524
rect 44508 13484 44640 13512
rect 44508 13472 44514 13484
rect 44634 13472 44640 13484
rect 44692 13472 44698 13524
rect 45094 13472 45100 13524
rect 45152 13512 45158 13524
rect 50430 13512 50436 13524
rect 45152 13484 50436 13512
rect 45152 13472 45158 13484
rect 50430 13472 50436 13484
rect 50488 13472 50494 13524
rect 50617 13515 50675 13521
rect 50617 13481 50629 13515
rect 50663 13512 50675 13515
rect 51258 13512 51264 13524
rect 50663 13484 51264 13512
rect 50663 13481 50675 13484
rect 50617 13475 50675 13481
rect 51258 13472 51264 13484
rect 51316 13472 51322 13524
rect 51534 13512 51540 13524
rect 51368 13484 51540 13512
rect 39942 13404 39948 13456
rect 40000 13444 40006 13456
rect 45278 13444 45284 13456
rect 40000 13416 40724 13444
rect 40000 13404 40006 13416
rect 39853 13379 39911 13385
rect 39853 13345 39865 13379
rect 39899 13376 39911 13379
rect 40402 13376 40408 13388
rect 39899 13348 40408 13376
rect 39899 13345 39911 13348
rect 39853 13339 39911 13345
rect 40402 13336 40408 13348
rect 40460 13336 40466 13388
rect 34957 13311 35015 13317
rect 34957 13308 34969 13311
rect 34848 13280 34969 13308
rect 34848 13268 34854 13280
rect 34957 13277 34969 13280
rect 35003 13277 35015 13311
rect 39117 13311 39175 13317
rect 34957 13271 35015 13277
rect 35084 13280 39068 13308
rect 30374 13240 30380 13252
rect 30024 13212 30380 13240
rect 30374 13200 30380 13212
rect 30432 13200 30438 13252
rect 30576 13212 31754 13240
rect 25179 13144 26004 13172
rect 25179 13141 25191 13144
rect 25133 13135 25191 13141
rect 26050 13132 26056 13184
rect 26108 13172 26114 13184
rect 26108 13144 26153 13172
rect 26108 13132 26114 13144
rect 26234 13132 26240 13184
rect 26292 13172 26298 13184
rect 27157 13175 27215 13181
rect 27157 13172 27169 13175
rect 26292 13144 27169 13172
rect 26292 13132 26298 13144
rect 27157 13141 27169 13144
rect 27203 13141 27215 13175
rect 27157 13135 27215 13141
rect 27798 13132 27804 13184
rect 27856 13172 27862 13184
rect 27985 13175 28043 13181
rect 27985 13172 27997 13175
rect 27856 13144 27997 13172
rect 27856 13132 27862 13144
rect 27985 13141 27997 13144
rect 28031 13141 28043 13175
rect 27985 13135 28043 13141
rect 29822 13132 29828 13184
rect 29880 13172 29886 13184
rect 30576 13172 30604 13212
rect 29880 13144 30604 13172
rect 29880 13132 29886 13144
rect 30650 13132 30656 13184
rect 30708 13172 30714 13184
rect 30929 13175 30987 13181
rect 30929 13172 30941 13175
rect 30708 13144 30941 13172
rect 30708 13132 30714 13144
rect 30929 13141 30941 13144
rect 30975 13141 30987 13175
rect 31726 13172 31754 13212
rect 32674 13200 32680 13252
rect 32732 13240 32738 13252
rect 32769 13243 32827 13249
rect 32769 13240 32781 13243
rect 32732 13212 32781 13240
rect 32732 13200 32738 13212
rect 32769 13209 32781 13212
rect 32815 13209 32827 13243
rect 33229 13243 33287 13249
rect 33229 13240 33241 13243
rect 32769 13203 32827 13209
rect 32876 13212 33241 13240
rect 32876 13172 32904 13212
rect 33229 13209 33241 13212
rect 33275 13209 33287 13243
rect 33229 13203 33287 13209
rect 33594 13200 33600 13252
rect 33652 13240 33658 13252
rect 35084 13240 35112 13280
rect 33652 13212 35112 13240
rect 36449 13243 36507 13249
rect 33652 13200 33658 13212
rect 36449 13209 36461 13243
rect 36495 13240 36507 13243
rect 38930 13240 38936 13252
rect 36495 13212 38936 13240
rect 36495 13209 36507 13212
rect 36449 13203 36507 13209
rect 38930 13200 38936 13212
rect 38988 13200 38994 13252
rect 39040 13240 39068 13280
rect 39117 13277 39129 13311
rect 39163 13277 39175 13311
rect 39298 13308 39304 13320
rect 39259 13280 39304 13308
rect 39117 13271 39175 13277
rect 39298 13268 39304 13280
rect 39356 13268 39362 13320
rect 39390 13268 39396 13320
rect 39448 13308 39454 13320
rect 40126 13308 40132 13320
rect 39448 13280 39493 13308
rect 40087 13280 40132 13308
rect 39448 13268 39454 13280
rect 40126 13268 40132 13280
rect 40184 13268 40190 13320
rect 40696 13308 40724 13416
rect 43272 13416 45284 13444
rect 40770 13336 40776 13388
rect 40828 13376 40834 13388
rect 40828 13348 41644 13376
rect 40828 13336 40834 13348
rect 41417 13311 41475 13317
rect 41417 13308 41429 13311
rect 40696 13280 41429 13308
rect 41417 13277 41429 13280
rect 41463 13308 41475 13311
rect 41506 13308 41512 13320
rect 41463 13280 41512 13308
rect 41463 13277 41475 13280
rect 41417 13271 41475 13277
rect 41506 13268 41512 13280
rect 41564 13268 41570 13320
rect 41616 13317 41644 13348
rect 41601 13311 41659 13317
rect 41601 13277 41613 13311
rect 41647 13277 41659 13311
rect 41601 13271 41659 13277
rect 41690 13268 41696 13320
rect 41748 13308 41754 13320
rect 41748 13280 42196 13308
rect 41748 13268 41754 13280
rect 41322 13240 41328 13252
rect 39040 13212 41328 13240
rect 41322 13200 41328 13212
rect 41380 13200 41386 13252
rect 42168 13240 42196 13280
rect 42242 13268 42248 13320
rect 42300 13308 42306 13320
rect 42300 13280 42748 13308
rect 42300 13268 42306 13280
rect 42720 13252 42748 13280
rect 42794 13268 42800 13320
rect 42852 13308 42858 13320
rect 43272 13308 43300 13416
rect 45278 13404 45284 13416
rect 45336 13404 45342 13456
rect 47213 13447 47271 13453
rect 47213 13413 47225 13447
rect 47259 13444 47271 13447
rect 47762 13444 47768 13456
rect 47259 13416 47768 13444
rect 47259 13413 47271 13416
rect 47213 13407 47271 13413
rect 47762 13404 47768 13416
rect 47820 13404 47826 13456
rect 47854 13404 47860 13456
rect 47912 13444 47918 13456
rect 48682 13444 48688 13456
rect 47912 13416 48688 13444
rect 47912 13404 47918 13416
rect 48682 13404 48688 13416
rect 48740 13404 48746 13456
rect 49145 13447 49203 13453
rect 49145 13413 49157 13447
rect 49191 13444 49203 13447
rect 49191 13416 49280 13444
rect 49191 13413 49203 13416
rect 49145 13407 49203 13413
rect 44266 13336 44272 13388
rect 44324 13376 44330 13388
rect 45462 13376 45468 13388
rect 44324 13348 45468 13376
rect 44324 13336 44330 13348
rect 45462 13336 45468 13348
rect 45520 13336 45526 13388
rect 45738 13336 45744 13388
rect 45796 13376 45802 13388
rect 45833 13379 45891 13385
rect 45833 13376 45845 13379
rect 45796 13348 45845 13376
rect 45796 13336 45802 13348
rect 45833 13345 45845 13348
rect 45879 13345 45891 13379
rect 45833 13339 45891 13345
rect 47670 13336 47676 13388
rect 47728 13376 47734 13388
rect 48866 13376 48872 13388
rect 47728 13348 48872 13376
rect 47728 13336 47734 13348
rect 48866 13336 48872 13348
rect 48924 13336 48930 13388
rect 49050 13376 49056 13388
rect 49011 13348 49056 13376
rect 49050 13336 49056 13348
rect 49108 13336 49114 13388
rect 49252 13376 49280 13416
rect 49786 13404 49792 13456
rect 49844 13444 49850 13456
rect 50338 13444 50344 13456
rect 49844 13416 50344 13444
rect 49844 13404 49850 13416
rect 50338 13404 50344 13416
rect 50396 13404 50402 13456
rect 50522 13404 50528 13456
rect 50580 13444 50586 13456
rect 51368 13444 51396 13484
rect 51534 13472 51540 13484
rect 51592 13472 51598 13524
rect 51718 13472 51724 13524
rect 51776 13512 51782 13524
rect 51997 13515 52055 13521
rect 51997 13512 52009 13515
rect 51776 13484 52009 13512
rect 51776 13472 51782 13484
rect 51997 13481 52009 13484
rect 52043 13481 52055 13515
rect 54938 13512 54944 13524
rect 51997 13475 52055 13481
rect 52380 13484 54944 13512
rect 52380 13444 52408 13484
rect 54938 13472 54944 13484
rect 54996 13472 55002 13524
rect 55030 13472 55036 13524
rect 55088 13512 55094 13524
rect 55309 13515 55367 13521
rect 55309 13512 55321 13515
rect 55088 13484 55321 13512
rect 55088 13472 55094 13484
rect 55309 13481 55321 13484
rect 55355 13481 55367 13515
rect 55309 13475 55367 13481
rect 55953 13515 56011 13521
rect 55953 13481 55965 13515
rect 55999 13512 56011 13515
rect 58342 13512 58348 13524
rect 55999 13484 58348 13512
rect 55999 13481 56011 13484
rect 55953 13475 56011 13481
rect 58342 13472 58348 13484
rect 58400 13472 58406 13524
rect 60001 13515 60059 13521
rect 60001 13481 60013 13515
rect 60047 13512 60059 13515
rect 61654 13512 61660 13524
rect 60047 13484 61660 13512
rect 60047 13481 60059 13484
rect 60001 13475 60059 13481
rect 61654 13472 61660 13484
rect 61712 13472 61718 13524
rect 61841 13515 61899 13521
rect 61841 13481 61853 13515
rect 61887 13512 61899 13515
rect 63586 13512 63592 13524
rect 61887 13484 63448 13512
rect 63547 13484 63592 13512
rect 61887 13481 61899 13484
rect 61841 13475 61899 13481
rect 50580 13416 51396 13444
rect 52012 13416 52408 13444
rect 52457 13447 52515 13453
rect 50580 13404 50586 13416
rect 50154 13376 50160 13388
rect 49252 13348 50160 13376
rect 50154 13336 50160 13348
rect 50212 13336 50218 13388
rect 51258 13376 51264 13388
rect 50264 13348 51264 13376
rect 42852 13280 43300 13308
rect 44545 13311 44603 13317
rect 42852 13268 42858 13280
rect 44545 13277 44557 13311
rect 44591 13308 44603 13311
rect 45922 13308 45928 13320
rect 44591 13280 45928 13308
rect 44591 13277 44603 13280
rect 44545 13271 44603 13277
rect 45922 13268 45928 13280
rect 45980 13268 45986 13320
rect 47026 13308 47032 13320
rect 46032 13280 47032 13308
rect 42490 13243 42548 13249
rect 42490 13240 42502 13243
rect 42168 13212 42502 13240
rect 42490 13209 42502 13212
rect 42536 13209 42548 13243
rect 42490 13203 42548 13209
rect 42702 13200 42708 13252
rect 42760 13200 42766 13252
rect 43070 13200 43076 13252
rect 43128 13240 43134 13252
rect 45281 13243 45339 13249
rect 45281 13240 45293 13243
rect 43128 13212 45293 13240
rect 43128 13200 43134 13212
rect 45281 13209 45293 13212
rect 45327 13240 45339 13243
rect 45646 13240 45652 13252
rect 45327 13212 45652 13240
rect 45327 13209 45339 13212
rect 45281 13203 45339 13209
rect 45646 13200 45652 13212
rect 45704 13240 45710 13252
rect 46032 13240 46060 13280
rect 47026 13268 47032 13280
rect 47084 13308 47090 13320
rect 47581 13311 47639 13317
rect 47581 13308 47593 13311
rect 47084 13280 47593 13308
rect 47084 13268 47090 13280
rect 47581 13277 47593 13280
rect 47627 13277 47639 13311
rect 47581 13271 47639 13277
rect 47857 13311 47915 13317
rect 47857 13277 47869 13311
rect 47903 13308 47915 13311
rect 47946 13308 47952 13320
rect 47903 13280 47952 13308
rect 47903 13277 47915 13280
rect 47857 13271 47915 13277
rect 47946 13268 47952 13280
rect 48004 13308 48010 13320
rect 48130 13308 48136 13320
rect 48004 13280 48136 13308
rect 48004 13268 48010 13280
rect 48130 13268 48136 13280
rect 48188 13268 48194 13320
rect 48682 13268 48688 13320
rect 48740 13308 48746 13320
rect 48961 13311 49019 13317
rect 48961 13308 48973 13311
rect 48740 13280 48973 13308
rect 48740 13268 48746 13280
rect 48961 13277 48973 13280
rect 49007 13277 49019 13311
rect 48961 13271 49019 13277
rect 49234 13268 49240 13320
rect 49292 13308 49298 13320
rect 49418 13308 49424 13320
rect 49292 13280 49337 13308
rect 49379 13280 49424 13308
rect 49292 13268 49298 13280
rect 49418 13268 49424 13280
rect 49476 13268 49482 13320
rect 49510 13268 49516 13320
rect 49568 13308 49574 13320
rect 50264 13317 50292 13348
rect 51258 13336 51264 13348
rect 51316 13336 51322 13388
rect 52012 13376 52040 13416
rect 52457 13413 52469 13447
rect 52503 13444 52515 13447
rect 54386 13444 54392 13456
rect 52503 13416 54392 13444
rect 52503 13413 52515 13416
rect 52457 13407 52515 13413
rect 54386 13404 54392 13416
rect 54444 13404 54450 13456
rect 56689 13447 56747 13453
rect 56689 13444 56701 13447
rect 55416 13416 56701 13444
rect 51368 13348 52040 13376
rect 50249 13311 50307 13317
rect 50249 13308 50261 13311
rect 49568 13280 50261 13308
rect 49568 13268 49574 13280
rect 50249 13277 50261 13280
rect 50295 13277 50307 13311
rect 50430 13308 50436 13320
rect 50391 13280 50436 13308
rect 50249 13271 50307 13277
rect 50430 13268 50436 13280
rect 50488 13268 50494 13320
rect 45704 13212 46060 13240
rect 46100 13243 46158 13249
rect 45704 13200 45710 13212
rect 46100 13209 46112 13243
rect 46146 13240 46158 13243
rect 46382 13240 46388 13252
rect 46146 13212 46388 13240
rect 46146 13209 46158 13212
rect 46100 13203 46158 13209
rect 46382 13200 46388 13212
rect 46440 13200 46446 13252
rect 48314 13240 48320 13252
rect 46492 13212 48320 13240
rect 31726 13144 32904 13172
rect 30929 13135 30987 13141
rect 32950 13132 32956 13184
rect 33008 13172 33014 13184
rect 33137 13175 33195 13181
rect 33137 13172 33149 13175
rect 33008 13144 33149 13172
rect 33008 13132 33014 13144
rect 33137 13141 33149 13144
rect 33183 13141 33195 13175
rect 33137 13135 33195 13141
rect 34057 13175 34115 13181
rect 34057 13141 34069 13175
rect 34103 13172 34115 13175
rect 34422 13172 34428 13184
rect 34103 13144 34428 13172
rect 34103 13141 34115 13144
rect 34057 13135 34115 13141
rect 34422 13132 34428 13144
rect 34480 13132 34486 13184
rect 34606 13132 34612 13184
rect 34664 13172 34670 13184
rect 35894 13172 35900 13184
rect 34664 13144 35900 13172
rect 34664 13132 34670 13144
rect 35894 13132 35900 13144
rect 35952 13132 35958 13184
rect 36081 13175 36139 13181
rect 36081 13141 36093 13175
rect 36127 13172 36139 13175
rect 36722 13172 36728 13184
rect 36127 13144 36728 13172
rect 36127 13141 36139 13144
rect 36081 13135 36139 13141
rect 36722 13132 36728 13144
rect 36780 13132 36786 13184
rect 36906 13132 36912 13184
rect 36964 13172 36970 13184
rect 41138 13172 41144 13184
rect 36964 13144 41144 13172
rect 36964 13132 36970 13144
rect 41138 13132 41144 13144
rect 41196 13132 41202 13184
rect 41785 13175 41843 13181
rect 41785 13141 41797 13175
rect 41831 13172 41843 13175
rect 42334 13172 42340 13184
rect 41831 13144 42340 13172
rect 41831 13141 41843 13144
rect 41785 13135 41843 13141
rect 42334 13132 42340 13144
rect 42392 13132 42398 13184
rect 43438 13132 43444 13184
rect 43496 13172 43502 13184
rect 46492 13172 46520 13212
rect 48314 13200 48320 13212
rect 48372 13200 48378 13252
rect 48777 13243 48835 13249
rect 48777 13209 48789 13243
rect 48823 13240 48835 13243
rect 51368 13240 51396 13348
rect 52086 13336 52092 13388
rect 52144 13376 52150 13388
rect 52917 13379 52975 13385
rect 52917 13376 52929 13379
rect 52144 13348 52929 13376
rect 52144 13336 52150 13348
rect 52917 13345 52929 13348
rect 52963 13345 52975 13379
rect 52917 13339 52975 13345
rect 53101 13379 53159 13385
rect 53101 13345 53113 13379
rect 53147 13376 53159 13379
rect 53466 13376 53472 13388
rect 53147 13348 53472 13376
rect 53147 13345 53159 13348
rect 53101 13339 53159 13345
rect 53466 13336 53472 13348
rect 53524 13336 53530 13388
rect 55416 13376 55444 13416
rect 56689 13413 56701 13416
rect 56735 13444 56747 13447
rect 59446 13444 59452 13456
rect 56735 13416 59452 13444
rect 56735 13413 56747 13416
rect 56689 13407 56747 13413
rect 59446 13404 59452 13416
rect 59504 13404 59510 13456
rect 60274 13404 60280 13456
rect 60332 13444 60338 13456
rect 60734 13444 60740 13456
rect 60332 13416 60740 13444
rect 60332 13404 60338 13416
rect 60734 13404 60740 13416
rect 60792 13404 60798 13456
rect 60826 13404 60832 13456
rect 60884 13404 60890 13456
rect 61013 13447 61071 13453
rect 61013 13413 61025 13447
rect 61059 13444 61071 13447
rect 61102 13444 61108 13456
rect 61059 13416 61108 13444
rect 61059 13413 61071 13416
rect 61013 13407 61071 13413
rect 61102 13404 61108 13416
rect 61160 13404 61166 13456
rect 60844 13376 60872 13404
rect 63420 13376 63448 13484
rect 63586 13472 63592 13484
rect 63644 13472 63650 13524
rect 64506 13472 64512 13524
rect 64564 13512 64570 13524
rect 69382 13512 69388 13524
rect 64564 13484 69388 13512
rect 64564 13472 64570 13484
rect 69382 13472 69388 13484
rect 69440 13472 69446 13524
rect 72326 13512 72332 13524
rect 69492 13484 72332 13512
rect 64414 13404 64420 13456
rect 64472 13444 64478 13456
rect 64472 13416 65840 13444
rect 64472 13404 64478 13416
rect 53576 13348 55444 13376
rect 55968 13348 59492 13376
rect 60844 13348 62344 13376
rect 63420 13348 64828 13376
rect 53576 13324 53604 13348
rect 51445 13311 51503 13317
rect 51445 13277 51457 13311
rect 51491 13277 51503 13311
rect 51810 13308 51816 13320
rect 51771 13280 51816 13308
rect 51445 13271 51503 13277
rect 48823 13212 51396 13240
rect 48823 13209 48835 13212
rect 48777 13203 48835 13209
rect 43496 13144 46520 13172
rect 43496 13132 43502 13144
rect 47762 13132 47768 13184
rect 47820 13172 47826 13184
rect 48682 13172 48688 13184
rect 47820 13144 48688 13172
rect 47820 13132 47826 13144
rect 48682 13132 48688 13144
rect 48740 13132 48746 13184
rect 51460 13172 51488 13271
rect 51810 13268 51816 13280
rect 51868 13268 51874 13320
rect 52178 13268 52184 13320
rect 52236 13308 52242 13320
rect 52236 13280 52776 13308
rect 52236 13268 52242 13280
rect 51626 13240 51632 13252
rect 51587 13212 51632 13240
rect 51626 13200 51632 13212
rect 51684 13200 51690 13252
rect 51721 13243 51779 13249
rect 51721 13209 51733 13243
rect 51767 13240 51779 13243
rect 52454 13240 52460 13252
rect 51767 13212 52460 13240
rect 51767 13209 51779 13212
rect 51721 13203 51779 13209
rect 52454 13200 52460 13212
rect 52512 13200 52518 13252
rect 52748 13240 52776 13280
rect 52822 13268 52828 13320
rect 52880 13308 52886 13320
rect 53573 13308 53604 13324
rect 53668 13317 53880 13318
rect 52880 13280 52925 13308
rect 53484 13296 53604 13308
rect 53653 13311 53880 13317
rect 53484 13280 53601 13296
rect 52880 13268 52886 13280
rect 53484 13240 53512 13280
rect 53653 13277 53665 13311
rect 53699 13308 53880 13311
rect 54110 13308 54116 13320
rect 53699 13290 54116 13308
rect 53699 13277 53711 13290
rect 53852 13280 54116 13290
rect 53653 13271 53711 13277
rect 54110 13268 54116 13280
rect 54168 13268 54174 13320
rect 54386 13268 54392 13320
rect 54444 13308 54450 13320
rect 55493 13311 55551 13317
rect 55493 13308 55505 13311
rect 54444 13280 55505 13308
rect 54444 13268 54450 13280
rect 55493 13277 55505 13280
rect 55539 13277 55551 13311
rect 55493 13271 55551 13277
rect 55861 13311 55919 13317
rect 55861 13277 55873 13311
rect 55907 13277 55919 13311
rect 55861 13271 55919 13277
rect 52748 13212 53512 13240
rect 53837 13243 53895 13249
rect 53837 13209 53849 13243
rect 53883 13209 53895 13243
rect 53837 13203 53895 13209
rect 52546 13172 52552 13184
rect 51460 13144 52552 13172
rect 52546 13132 52552 13144
rect 52604 13132 52610 13184
rect 53852 13172 53880 13203
rect 53926 13200 53932 13252
rect 53984 13240 53990 13252
rect 54297 13243 54355 13249
rect 54297 13240 54309 13243
rect 53984 13212 54309 13240
rect 53984 13200 53990 13212
rect 54297 13209 54309 13212
rect 54343 13240 54355 13243
rect 55122 13240 55128 13252
rect 54343 13212 55128 13240
rect 54343 13209 54355 13212
rect 54297 13203 54355 13209
rect 55122 13200 55128 13212
rect 55180 13200 55186 13252
rect 55306 13200 55312 13252
rect 55364 13240 55370 13252
rect 55876 13240 55904 13271
rect 55364 13212 55904 13240
rect 55364 13200 55370 13212
rect 54110 13172 54116 13184
rect 53852 13144 54116 13172
rect 54110 13132 54116 13144
rect 54168 13132 54174 13184
rect 54386 13132 54392 13184
rect 54444 13172 54450 13184
rect 54444 13144 54489 13172
rect 54444 13132 54450 13144
rect 55398 13132 55404 13184
rect 55456 13172 55462 13184
rect 55968 13172 55996 13348
rect 56962 13268 56968 13320
rect 57020 13308 57026 13320
rect 57057 13311 57115 13317
rect 57057 13308 57069 13311
rect 57020 13280 57069 13308
rect 57020 13268 57026 13280
rect 57057 13277 57069 13280
rect 57103 13277 57115 13311
rect 57057 13271 57115 13277
rect 57333 13311 57391 13317
rect 57333 13277 57345 13311
rect 57379 13308 57391 13311
rect 57882 13308 57888 13320
rect 57379 13280 57888 13308
rect 57379 13277 57391 13280
rect 57333 13271 57391 13277
rect 56042 13200 56048 13252
rect 56100 13240 56106 13252
rect 56505 13243 56563 13249
rect 56505 13240 56517 13243
rect 56100 13212 56517 13240
rect 56100 13200 56106 13212
rect 56505 13209 56517 13212
rect 56551 13209 56563 13243
rect 57072 13240 57100 13271
rect 57882 13268 57888 13280
rect 57940 13268 57946 13320
rect 58158 13268 58164 13320
rect 58216 13308 58222 13320
rect 58253 13311 58311 13317
rect 58253 13308 58265 13311
rect 58216 13280 58265 13308
rect 58216 13268 58222 13280
rect 58253 13277 58265 13280
rect 58299 13277 58311 13311
rect 58253 13271 58311 13277
rect 58342 13268 58348 13320
rect 58400 13308 58406 13320
rect 59354 13308 59360 13320
rect 58400 13280 59360 13308
rect 58400 13268 58406 13280
rect 59354 13268 59360 13280
rect 59412 13268 59418 13320
rect 59464 13317 59492 13348
rect 59449 13311 59507 13317
rect 59449 13277 59461 13311
rect 59495 13277 59507 13311
rect 59814 13308 59820 13320
rect 59775 13280 59820 13308
rect 59449 13271 59507 13277
rect 59814 13268 59820 13280
rect 59872 13268 59878 13320
rect 60461 13311 60519 13317
rect 60461 13277 60473 13311
rect 60507 13277 60519 13311
rect 60461 13271 60519 13277
rect 59262 13240 59268 13252
rect 57072 13212 59268 13240
rect 56505 13203 56563 13209
rect 59262 13200 59268 13212
rect 59320 13200 59326 13252
rect 59630 13240 59636 13252
rect 59591 13212 59636 13240
rect 59630 13200 59636 13212
rect 59688 13200 59694 13252
rect 59725 13243 59783 13249
rect 59725 13209 59737 13243
rect 59771 13209 59783 13243
rect 59725 13203 59783 13209
rect 55456 13144 55996 13172
rect 55456 13132 55462 13144
rect 56134 13132 56140 13184
rect 56192 13172 56198 13184
rect 57514 13172 57520 13184
rect 56192 13144 57520 13172
rect 56192 13132 56198 13144
rect 57514 13132 57520 13144
rect 57572 13172 57578 13184
rect 58483 13175 58541 13181
rect 58483 13172 58495 13175
rect 57572 13144 58495 13172
rect 57572 13132 57578 13144
rect 58483 13141 58495 13144
rect 58529 13172 58541 13175
rect 58894 13172 58900 13184
rect 58529 13144 58900 13172
rect 58529 13141 58541 13144
rect 58483 13135 58541 13141
rect 58894 13132 58900 13144
rect 58952 13172 58958 13184
rect 59740 13172 59768 13203
rect 58952 13144 59768 13172
rect 60476 13172 60504 13271
rect 60550 13268 60556 13320
rect 60608 13308 60614 13320
rect 60734 13311 60792 13317
rect 60734 13308 60746 13311
rect 60608 13280 60746 13308
rect 60608 13268 60614 13280
rect 60734 13277 60746 13280
rect 60780 13277 60792 13311
rect 60734 13271 60792 13277
rect 60826 13268 60832 13320
rect 60884 13317 60890 13320
rect 60884 13308 60892 13317
rect 60884 13280 60929 13308
rect 60884 13271 60892 13280
rect 60884 13268 60890 13271
rect 61010 13268 61016 13320
rect 61068 13308 61074 13320
rect 61473 13311 61531 13317
rect 61473 13308 61485 13311
rect 61068 13280 61485 13308
rect 61068 13268 61074 13280
rect 61473 13277 61485 13280
rect 61519 13277 61531 13311
rect 61654 13308 61660 13320
rect 61615 13280 61660 13308
rect 61473 13271 61531 13277
rect 61654 13268 61660 13280
rect 61712 13268 61718 13320
rect 62206 13308 62212 13320
rect 62167 13280 62212 13308
rect 62206 13268 62212 13280
rect 62264 13268 62270 13320
rect 62316 13308 62344 13348
rect 64800 13317 64828 13348
rect 65812 13317 65840 13416
rect 66254 13404 66260 13456
rect 66312 13444 66318 13456
rect 67637 13447 67695 13453
rect 67637 13444 67649 13447
rect 66312 13416 67649 13444
rect 66312 13404 66318 13416
rect 67637 13413 67649 13416
rect 67683 13413 67695 13447
rect 67637 13407 67695 13413
rect 68281 13447 68339 13453
rect 68281 13413 68293 13447
rect 68327 13413 68339 13447
rect 68281 13407 68339 13413
rect 68296 13376 68324 13407
rect 68922 13404 68928 13456
rect 68980 13444 68986 13456
rect 69492 13444 69520 13484
rect 68980 13416 69520 13444
rect 68980 13404 68986 13416
rect 68296 13348 68968 13376
rect 63957 13311 64015 13317
rect 63957 13308 63969 13311
rect 62316 13280 63969 13308
rect 63957 13277 63969 13280
rect 64003 13277 64015 13311
rect 63957 13271 64015 13277
rect 64785 13311 64843 13317
rect 64785 13277 64797 13311
rect 64831 13277 64843 13311
rect 64785 13271 64843 13277
rect 65797 13311 65855 13317
rect 65797 13277 65809 13311
rect 65843 13277 65855 13311
rect 65797 13271 65855 13277
rect 67913 13311 67971 13317
rect 67913 13277 67925 13311
rect 67959 13308 67971 13311
rect 68462 13308 68468 13320
rect 67959 13280 68468 13308
rect 67959 13277 67971 13280
rect 67913 13271 67971 13277
rect 68462 13268 68468 13280
rect 68520 13268 68526 13320
rect 68557 13311 68615 13317
rect 68557 13277 68569 13311
rect 68603 13308 68615 13311
rect 68830 13308 68836 13320
rect 68603 13280 68836 13308
rect 68603 13277 68615 13280
rect 68557 13271 68615 13277
rect 68830 13268 68836 13280
rect 68888 13268 68894 13320
rect 68940 13317 68968 13348
rect 69124 13348 69888 13376
rect 69124 13317 69152 13348
rect 69860 13317 69888 13348
rect 68925 13311 68983 13317
rect 68925 13277 68937 13311
rect 68971 13277 68983 13311
rect 68925 13271 68983 13277
rect 69109 13311 69167 13317
rect 69109 13277 69121 13311
rect 69155 13277 69167 13311
rect 69109 13271 69167 13277
rect 69293 13311 69351 13317
rect 69293 13277 69305 13311
rect 69339 13277 69351 13311
rect 69293 13271 69351 13277
rect 69845 13311 69903 13317
rect 69845 13277 69857 13311
rect 69891 13277 69903 13311
rect 69845 13271 69903 13277
rect 70029 13311 70087 13317
rect 70029 13277 70041 13311
rect 70075 13277 70087 13311
rect 70210 13308 70216 13320
rect 70171 13280 70216 13308
rect 70029 13271 70087 13277
rect 60642 13240 60648 13252
rect 60603 13212 60648 13240
rect 60642 13200 60648 13212
rect 60700 13200 60706 13252
rect 62476 13243 62534 13249
rect 62476 13209 62488 13243
rect 62522 13240 62534 13243
rect 62522 13212 65656 13240
rect 62522 13209 62534 13212
rect 62476 13203 62534 13209
rect 62666 13172 62672 13184
rect 60476 13144 62672 13172
rect 58952 13132 58958 13144
rect 62666 13132 62672 13144
rect 62724 13132 62730 13184
rect 63310 13132 63316 13184
rect 63368 13172 63374 13184
rect 64141 13175 64199 13181
rect 64141 13172 64153 13175
rect 63368 13144 64153 13172
rect 63368 13132 63374 13144
rect 64141 13141 64153 13144
rect 64187 13172 64199 13175
rect 64322 13172 64328 13184
rect 64187 13144 64328 13172
rect 64187 13141 64199 13144
rect 64141 13135 64199 13141
rect 64322 13132 64328 13144
rect 64380 13132 64386 13184
rect 64598 13172 64604 13184
rect 64559 13144 64604 13172
rect 64598 13132 64604 13144
rect 64656 13132 64662 13184
rect 65628 13181 65656 13212
rect 67634 13200 67640 13252
rect 67692 13240 67698 13252
rect 68186 13240 68192 13252
rect 67692 13212 68192 13240
rect 67692 13200 67698 13212
rect 68186 13200 68192 13212
rect 68244 13240 68250 13252
rect 68281 13243 68339 13249
rect 68281 13240 68293 13243
rect 68244 13212 68293 13240
rect 68244 13200 68250 13212
rect 68281 13209 68293 13212
rect 68327 13209 68339 13243
rect 68281 13203 68339 13209
rect 68370 13200 68376 13252
rect 68428 13240 68434 13252
rect 69201 13243 69259 13249
rect 69201 13240 69213 13243
rect 68428 13212 69213 13240
rect 68428 13200 68434 13212
rect 69201 13209 69213 13212
rect 69247 13209 69259 13243
rect 69201 13203 69259 13209
rect 65613 13175 65671 13181
rect 65613 13141 65625 13175
rect 65659 13141 65671 13175
rect 65613 13135 65671 13141
rect 67821 13175 67879 13181
rect 67821 13141 67833 13175
rect 67867 13172 67879 13175
rect 68094 13172 68100 13184
rect 67867 13144 68100 13172
rect 67867 13141 67879 13144
rect 67821 13135 67879 13141
rect 68094 13132 68100 13144
rect 68152 13172 68158 13184
rect 68465 13175 68523 13181
rect 68465 13172 68477 13175
rect 68152 13144 68477 13172
rect 68152 13132 68158 13144
rect 68465 13141 68477 13144
rect 68511 13141 68523 13175
rect 68465 13135 68523 13141
rect 68554 13132 68560 13184
rect 68612 13172 68618 13184
rect 69308 13172 69336 13271
rect 69658 13200 69664 13252
rect 69716 13240 69722 13252
rect 70044 13240 70072 13271
rect 70210 13268 70216 13280
rect 70268 13268 70274 13320
rect 70320 13317 70348 13484
rect 72326 13472 72332 13484
rect 72384 13472 72390 13524
rect 71866 13404 71872 13456
rect 71924 13444 71930 13456
rect 72145 13447 72203 13453
rect 72145 13444 72157 13447
rect 71924 13416 72157 13444
rect 71924 13404 71930 13416
rect 72145 13413 72157 13416
rect 72191 13413 72203 13447
rect 72145 13407 72203 13413
rect 70305 13311 70363 13317
rect 70305 13277 70317 13311
rect 70351 13277 70363 13311
rect 70762 13308 70768 13320
rect 70723 13280 70768 13308
rect 70305 13271 70363 13277
rect 70762 13268 70768 13280
rect 70820 13268 70826 13320
rect 71038 13317 71044 13320
rect 71032 13308 71044 13317
rect 70999 13280 71044 13308
rect 71032 13271 71044 13280
rect 71038 13268 71044 13271
rect 71096 13268 71102 13320
rect 86770 13268 86776 13320
rect 86828 13308 86834 13320
rect 88245 13311 88303 13317
rect 88245 13308 88257 13311
rect 86828 13280 88257 13308
rect 86828 13268 86834 13280
rect 88245 13277 88257 13280
rect 88291 13277 88303 13311
rect 88245 13271 88303 13277
rect 72234 13240 72240 13252
rect 69716 13212 72240 13240
rect 69716 13200 69722 13212
rect 72234 13200 72240 13212
rect 72292 13200 72298 13252
rect 68612 13144 69336 13172
rect 68612 13132 68618 13144
rect 69382 13132 69388 13184
rect 69440 13172 69446 13184
rect 69477 13175 69535 13181
rect 69477 13172 69489 13175
rect 69440 13144 69489 13172
rect 69440 13132 69446 13144
rect 69477 13141 69489 13144
rect 69523 13172 69535 13175
rect 72510 13172 72516 13184
rect 69523 13144 72516 13172
rect 69523 13141 69535 13144
rect 69477 13135 69535 13141
rect 72510 13132 72516 13144
rect 72568 13132 72574 13184
rect 88058 13172 88064 13184
rect 88019 13144 88064 13172
rect 88058 13132 88064 13144
rect 88116 13132 88122 13184
rect 1104 13082 88872 13104
rect 1104 13030 22898 13082
rect 22950 13030 22962 13082
rect 23014 13030 23026 13082
rect 23078 13030 23090 13082
rect 23142 13030 23154 13082
rect 23206 13030 44846 13082
rect 44898 13030 44910 13082
rect 44962 13030 44974 13082
rect 45026 13030 45038 13082
rect 45090 13030 45102 13082
rect 45154 13030 66794 13082
rect 66846 13030 66858 13082
rect 66910 13030 66922 13082
rect 66974 13030 66986 13082
rect 67038 13030 67050 13082
rect 67102 13030 88872 13082
rect 1104 13008 88872 13030
rect 6886 12940 22692 12968
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 6886 12832 6914 12940
rect 22002 12900 22008 12912
rect 19628 12872 22008 12900
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 1719 12804 6914 12832
rect 12406 12804 18613 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 3326 12724 3332 12776
rect 3384 12764 3390 12776
rect 3970 12764 3976 12776
rect 3384 12736 3976 12764
rect 3384 12724 3390 12736
rect 3970 12724 3976 12736
rect 4028 12764 4034 12776
rect 12406 12764 12434 12804
rect 18601 12801 18613 12804
rect 18647 12832 18659 12835
rect 19518 12832 19524 12844
rect 18647 12804 19524 12832
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 19518 12792 19524 12804
rect 19576 12792 19582 12844
rect 19058 12764 19064 12776
rect 4028 12736 12434 12764
rect 19019 12736 19064 12764
rect 4028 12724 4034 12736
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 19628 12696 19656 12872
rect 22002 12860 22008 12872
rect 22060 12860 22066 12912
rect 19797 12835 19855 12841
rect 19797 12801 19809 12835
rect 19843 12832 19855 12835
rect 19886 12832 19892 12844
rect 19843 12804 19892 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 19886 12792 19892 12804
rect 19944 12832 19950 12844
rect 20162 12832 20168 12844
rect 19944 12804 20168 12832
rect 19944 12792 19950 12804
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20404 12804 20637 12832
rect 20404 12792 20410 12804
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 22664 12832 22692 12940
rect 22738 12928 22744 12980
rect 22796 12968 22802 12980
rect 23477 12971 23535 12977
rect 23477 12968 23489 12971
rect 22796 12940 23489 12968
rect 22796 12928 22802 12940
rect 23477 12937 23489 12940
rect 23523 12937 23535 12971
rect 24486 12968 24492 12980
rect 24447 12940 24492 12968
rect 23477 12931 23535 12937
rect 24486 12928 24492 12940
rect 24544 12928 24550 12980
rect 25222 12968 25228 12980
rect 24964 12940 25228 12968
rect 24964 12909 24992 12940
rect 25222 12928 25228 12940
rect 25280 12928 25286 12980
rect 25406 12968 25412 12980
rect 25367 12940 25412 12968
rect 25406 12928 25412 12940
rect 25464 12928 25470 12980
rect 25498 12928 25504 12980
rect 25556 12968 25562 12980
rect 26421 12971 26479 12977
rect 26421 12968 26433 12971
rect 25556 12940 26433 12968
rect 25556 12928 25562 12940
rect 26421 12937 26433 12940
rect 26467 12937 26479 12971
rect 26421 12931 26479 12937
rect 26510 12928 26516 12980
rect 26568 12968 26574 12980
rect 28534 12968 28540 12980
rect 26568 12940 28540 12968
rect 26568 12928 26574 12940
rect 28534 12928 28540 12940
rect 28592 12928 28598 12980
rect 29089 12971 29147 12977
rect 29089 12937 29101 12971
rect 29135 12937 29147 12971
rect 29089 12931 29147 12937
rect 23661 12903 23719 12909
rect 23661 12869 23673 12903
rect 23707 12900 23719 12903
rect 24949 12903 25007 12909
rect 23707 12872 24808 12900
rect 23707 12869 23719 12872
rect 23661 12863 23719 12869
rect 24394 12832 24400 12844
rect 20772 12804 22600 12832
rect 22664 12804 24164 12832
rect 24355 12804 24400 12832
rect 20772 12792 20778 12804
rect 19702 12724 19708 12776
rect 19760 12764 19766 12776
rect 19760 12736 20024 12764
rect 19760 12724 19766 12736
rect 19628 12668 19932 12696
rect 18877 12631 18935 12637
rect 18877 12597 18889 12631
rect 18923 12628 18935 12631
rect 19794 12628 19800 12640
rect 18923 12600 19800 12628
rect 18923 12597 18935 12600
rect 18877 12591 18935 12597
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 19904 12637 19932 12668
rect 19889 12631 19947 12637
rect 19889 12597 19901 12631
rect 19935 12597 19947 12631
rect 19996 12628 20024 12736
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 20496 12736 22094 12764
rect 20496 12724 20502 12736
rect 20898 12696 20904 12708
rect 20732 12668 20904 12696
rect 20732 12637 20760 12668
rect 20898 12656 20904 12668
rect 20956 12656 20962 12708
rect 20257 12631 20315 12637
rect 20257 12628 20269 12631
rect 19996 12600 20269 12628
rect 19889 12591 19947 12597
rect 20257 12597 20269 12600
rect 20303 12597 20315 12631
rect 20257 12591 20315 12597
rect 20717 12631 20775 12637
rect 20717 12597 20729 12631
rect 20763 12597 20775 12631
rect 20717 12591 20775 12597
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21085 12631 21143 12637
rect 21085 12628 21097 12631
rect 20864 12600 21097 12628
rect 20864 12588 20870 12600
rect 21085 12597 21097 12600
rect 21131 12597 21143 12631
rect 22066 12628 22094 12736
rect 22572 12696 22600 12804
rect 23474 12724 23480 12776
rect 23532 12764 23538 12776
rect 23569 12767 23627 12773
rect 23569 12764 23581 12767
rect 23532 12736 23581 12764
rect 23532 12724 23538 12736
rect 23569 12733 23581 12736
rect 23615 12733 23627 12767
rect 23569 12727 23627 12733
rect 23750 12724 23756 12776
rect 23808 12764 23814 12776
rect 24029 12767 24087 12773
rect 23808 12736 23853 12764
rect 23808 12724 23814 12736
rect 24029 12733 24041 12767
rect 24075 12733 24087 12767
rect 24136 12764 24164 12804
rect 24394 12792 24400 12804
rect 24452 12792 24458 12844
rect 24780 12832 24808 12872
rect 24949 12869 24961 12903
rect 24995 12869 25007 12903
rect 26142 12900 26148 12912
rect 24949 12863 25007 12869
rect 25148 12872 26148 12900
rect 24854 12832 24860 12844
rect 24780 12804 24860 12832
rect 24854 12792 24860 12804
rect 24912 12792 24918 12844
rect 25148 12841 25176 12872
rect 26142 12860 26148 12872
rect 26200 12860 26206 12912
rect 29104 12900 29132 12931
rect 29178 12928 29184 12980
rect 29236 12968 29242 12980
rect 33870 12968 33876 12980
rect 29236 12940 33876 12968
rect 29236 12928 29242 12940
rect 33870 12928 33876 12940
rect 33928 12928 33934 12980
rect 36446 12968 36452 12980
rect 33980 12940 36452 12968
rect 30193 12903 30251 12909
rect 30193 12900 30205 12903
rect 26252 12872 29132 12900
rect 29196 12872 30205 12900
rect 26252 12841 26280 12872
rect 25133 12835 25191 12841
rect 25133 12801 25145 12835
rect 25179 12801 25191 12835
rect 25133 12795 25191 12801
rect 25225 12835 25283 12841
rect 25225 12801 25237 12835
rect 25271 12832 25283 12835
rect 25777 12835 25835 12841
rect 25777 12832 25789 12835
rect 25271 12804 25789 12832
rect 25271 12801 25283 12804
rect 25225 12795 25283 12801
rect 25777 12801 25789 12804
rect 25823 12801 25835 12835
rect 25777 12795 25835 12801
rect 26237 12835 26295 12841
rect 26237 12801 26249 12835
rect 26283 12801 26295 12835
rect 26510 12832 26516 12844
rect 26471 12804 26516 12832
rect 26237 12795 26295 12801
rect 26510 12792 26516 12804
rect 26568 12792 26574 12844
rect 29196 12832 29224 12872
rect 30193 12869 30205 12872
rect 30239 12869 30251 12903
rect 30193 12863 30251 12869
rect 31297 12903 31355 12909
rect 31297 12869 31309 12903
rect 31343 12900 31355 12903
rect 32490 12900 32496 12912
rect 31343 12872 32496 12900
rect 31343 12869 31355 12872
rect 31297 12863 31355 12869
rect 32490 12860 32496 12872
rect 32548 12900 32554 12912
rect 32548 12872 33088 12900
rect 32548 12860 32554 12872
rect 26620 12804 29224 12832
rect 30101 12835 30159 12841
rect 26620 12764 26648 12804
rect 30101 12801 30113 12835
rect 30147 12832 30159 12835
rect 30374 12832 30380 12844
rect 30147 12804 30380 12832
rect 30147 12801 30159 12804
rect 30101 12795 30159 12801
rect 30374 12792 30380 12804
rect 30432 12832 30438 12844
rect 30926 12832 30932 12844
rect 30432 12804 30932 12832
rect 30432 12792 30438 12804
rect 30926 12792 30932 12804
rect 30984 12792 30990 12844
rect 31665 12835 31723 12841
rect 31665 12801 31677 12835
rect 31711 12832 31723 12835
rect 31938 12832 31944 12844
rect 31711 12804 31944 12832
rect 31711 12801 31723 12804
rect 31665 12795 31723 12801
rect 31938 12792 31944 12804
rect 31996 12792 32002 12844
rect 32030 12792 32036 12844
rect 32088 12832 32094 12844
rect 32398 12832 32404 12844
rect 32088 12804 32404 12832
rect 32088 12792 32094 12804
rect 32398 12792 32404 12804
rect 32456 12792 32462 12844
rect 32582 12832 32588 12844
rect 32543 12804 32588 12832
rect 32582 12792 32588 12804
rect 32640 12792 32646 12844
rect 32677 12835 32735 12841
rect 32677 12801 32689 12835
rect 32723 12832 32735 12835
rect 32766 12832 32772 12844
rect 32723 12804 32772 12832
rect 32723 12801 32735 12804
rect 32677 12795 32735 12801
rect 32766 12792 32772 12804
rect 32824 12792 32830 12844
rect 33060 12841 33088 12872
rect 33045 12835 33103 12841
rect 33045 12801 33057 12835
rect 33091 12832 33103 12835
rect 33134 12832 33140 12844
rect 33091 12804 33140 12832
rect 33091 12801 33103 12804
rect 33045 12795 33103 12801
rect 33134 12792 33140 12804
rect 33192 12792 33198 12844
rect 33873 12835 33931 12841
rect 33873 12801 33885 12835
rect 33919 12832 33931 12835
rect 33980 12832 34008 12940
rect 36446 12928 36452 12940
rect 36504 12928 36510 12980
rect 36817 12971 36875 12977
rect 36817 12937 36829 12971
rect 36863 12968 36875 12971
rect 38286 12968 38292 12980
rect 36863 12940 38292 12968
rect 36863 12937 36875 12940
rect 36817 12931 36875 12937
rect 38286 12928 38292 12940
rect 38344 12928 38350 12980
rect 38470 12928 38476 12980
rect 38528 12968 38534 12980
rect 38565 12971 38623 12977
rect 38565 12968 38577 12971
rect 38528 12940 38577 12968
rect 38528 12928 38534 12940
rect 38565 12937 38577 12940
rect 38611 12937 38623 12971
rect 38565 12931 38623 12937
rect 41506 12928 41512 12980
rect 41564 12968 41570 12980
rect 42659 12971 42717 12977
rect 42659 12968 42671 12971
rect 41564 12940 42671 12968
rect 41564 12928 41570 12940
rect 42659 12937 42671 12940
rect 42705 12937 42717 12971
rect 45646 12968 45652 12980
rect 42659 12931 42717 12937
rect 43824 12940 45652 12968
rect 34057 12903 34115 12909
rect 34057 12869 34069 12903
rect 34103 12900 34115 12903
rect 34238 12900 34244 12912
rect 34103 12872 34244 12900
rect 34103 12869 34115 12872
rect 34057 12863 34115 12869
rect 34238 12860 34244 12872
rect 34296 12860 34302 12912
rect 34606 12900 34612 12912
rect 34348 12872 34612 12900
rect 33919 12804 34008 12832
rect 34149 12835 34207 12841
rect 33919 12801 33931 12804
rect 33873 12795 33931 12801
rect 34149 12801 34161 12835
rect 34195 12832 34207 12835
rect 34348 12832 34376 12872
rect 34606 12860 34612 12872
rect 34664 12860 34670 12912
rect 34793 12903 34851 12909
rect 34793 12869 34805 12903
rect 34839 12900 34851 12903
rect 35802 12900 35808 12912
rect 34839 12872 35808 12900
rect 34839 12869 34851 12872
rect 34793 12863 34851 12869
rect 35802 12860 35808 12872
rect 35860 12860 35866 12912
rect 36998 12860 37004 12912
rect 37056 12900 37062 12912
rect 38105 12903 38163 12909
rect 38105 12900 38117 12903
rect 37056 12872 38117 12900
rect 37056 12860 37062 12872
rect 38105 12869 38117 12872
rect 38151 12900 38163 12903
rect 38378 12900 38384 12912
rect 38151 12872 38384 12900
rect 38151 12869 38163 12872
rect 38105 12863 38163 12869
rect 38378 12860 38384 12872
rect 38436 12860 38442 12912
rect 38930 12860 38936 12912
rect 38988 12900 38994 12912
rect 39025 12903 39083 12909
rect 39025 12900 39037 12903
rect 38988 12872 39037 12900
rect 38988 12860 38994 12872
rect 39025 12869 39037 12872
rect 39071 12900 39083 12903
rect 39114 12900 39120 12912
rect 39071 12872 39120 12900
rect 39071 12869 39083 12872
rect 39025 12863 39083 12869
rect 39114 12860 39120 12872
rect 39172 12860 39178 12912
rect 40034 12860 40040 12912
rect 40092 12900 40098 12912
rect 40589 12903 40647 12909
rect 40589 12900 40601 12903
rect 40092 12872 40601 12900
rect 40092 12860 40098 12872
rect 40589 12869 40601 12872
rect 40635 12900 40647 12903
rect 40954 12900 40960 12912
rect 40635 12872 40960 12900
rect 40635 12869 40647 12872
rect 40589 12863 40647 12869
rect 40954 12860 40960 12872
rect 41012 12900 41018 12912
rect 42242 12900 42248 12912
rect 41012 12872 42248 12900
rect 41012 12860 41018 12872
rect 42242 12860 42248 12872
rect 42300 12860 42306 12912
rect 42886 12900 42892 12912
rect 42352 12872 42892 12900
rect 34514 12832 34520 12844
rect 34195 12804 34376 12832
rect 34475 12804 34520 12832
rect 34195 12801 34207 12804
rect 34149 12795 34207 12801
rect 34514 12792 34520 12804
rect 34572 12792 34578 12844
rect 34701 12835 34759 12841
rect 34701 12801 34713 12835
rect 34747 12801 34759 12835
rect 34882 12832 34888 12844
rect 34843 12804 34888 12832
rect 34701 12795 34759 12801
rect 24136 12736 26648 12764
rect 24029 12727 24087 12733
rect 23934 12696 23940 12708
rect 22572 12668 23940 12696
rect 23934 12656 23940 12668
rect 23992 12656 23998 12708
rect 24044 12696 24072 12727
rect 26694 12724 26700 12776
rect 26752 12764 26758 12776
rect 27433 12767 27491 12773
rect 27433 12764 27445 12767
rect 26752 12736 27445 12764
rect 26752 12724 26758 12736
rect 27433 12733 27445 12736
rect 27479 12764 27491 12767
rect 27801 12767 27859 12773
rect 27801 12764 27813 12767
rect 27479 12736 27813 12764
rect 27479 12733 27491 12736
rect 27433 12727 27491 12733
rect 27801 12733 27813 12736
rect 27847 12764 27859 12767
rect 27847 12736 28396 12764
rect 27847 12733 27859 12736
rect 27801 12727 27859 12733
rect 24210 12696 24216 12708
rect 24044 12668 24216 12696
rect 24210 12656 24216 12668
rect 24268 12656 24274 12708
rect 26145 12699 26203 12705
rect 26145 12665 26157 12699
rect 26191 12696 26203 12699
rect 26191 12668 27568 12696
rect 26191 12665 26203 12668
rect 26145 12659 26203 12665
rect 23382 12628 23388 12640
rect 22066 12600 23388 12628
rect 21085 12591 21143 12597
rect 23382 12588 23388 12600
rect 23440 12588 23446 12640
rect 25222 12588 25228 12640
rect 25280 12628 25286 12640
rect 26053 12631 26111 12637
rect 25280 12600 25325 12628
rect 25280 12588 25286 12600
rect 26053 12597 26065 12631
rect 26099 12628 26111 12631
rect 27246 12628 27252 12640
rect 26099 12600 27252 12628
rect 26099 12597 26111 12600
rect 26053 12591 26111 12597
rect 27246 12588 27252 12600
rect 27304 12588 27310 12640
rect 27540 12628 27568 12668
rect 27614 12656 27620 12708
rect 27672 12696 27678 12708
rect 28077 12699 28135 12705
rect 28077 12696 28089 12699
rect 27672 12668 28089 12696
rect 27672 12656 27678 12668
rect 28077 12665 28089 12668
rect 28123 12696 28135 12699
rect 28166 12696 28172 12708
rect 28123 12668 28172 12696
rect 28123 12665 28135 12668
rect 28077 12659 28135 12665
rect 28166 12656 28172 12668
rect 28224 12656 28230 12708
rect 28261 12631 28319 12637
rect 28261 12628 28273 12631
rect 27540 12600 28273 12628
rect 28261 12597 28273 12600
rect 28307 12597 28319 12631
rect 28368 12628 28396 12736
rect 28442 12724 28448 12776
rect 28500 12764 28506 12776
rect 28629 12767 28687 12773
rect 28629 12764 28641 12767
rect 28500 12736 28641 12764
rect 28500 12724 28506 12736
rect 28629 12733 28641 12736
rect 28675 12733 28687 12767
rect 28629 12727 28687 12733
rect 30285 12767 30343 12773
rect 30285 12733 30297 12767
rect 30331 12764 30343 12767
rect 32858 12764 32864 12776
rect 30331 12736 32864 12764
rect 30331 12733 30343 12736
rect 30285 12727 30343 12733
rect 32858 12724 32864 12736
rect 32916 12724 32922 12776
rect 33594 12764 33600 12776
rect 33060 12736 33600 12764
rect 28902 12696 28908 12708
rect 28863 12668 28908 12696
rect 28902 12656 28908 12668
rect 28960 12656 28966 12708
rect 33060 12696 33088 12736
rect 33594 12724 33600 12736
rect 33652 12724 33658 12776
rect 33689 12767 33747 12773
rect 33689 12733 33701 12767
rect 33735 12764 33747 12767
rect 34716 12764 34744 12795
rect 34882 12792 34888 12804
rect 34940 12792 34946 12844
rect 35434 12792 35440 12844
rect 35492 12832 35498 12844
rect 35529 12835 35587 12841
rect 35529 12832 35541 12835
rect 35492 12804 35541 12832
rect 35492 12792 35498 12804
rect 35529 12801 35541 12804
rect 35575 12801 35587 12835
rect 35529 12795 35587 12801
rect 35710 12792 35716 12844
rect 35768 12832 35774 12844
rect 35897 12835 35955 12841
rect 35768 12804 35813 12832
rect 35768 12792 35774 12804
rect 35897 12801 35909 12835
rect 35943 12801 35955 12835
rect 36538 12832 36544 12844
rect 36499 12804 36544 12832
rect 35897 12795 35955 12801
rect 33735 12736 34744 12764
rect 35912 12764 35940 12795
rect 36538 12792 36544 12804
rect 36596 12792 36602 12844
rect 36633 12835 36691 12841
rect 36633 12801 36645 12835
rect 36679 12801 36691 12835
rect 36633 12795 36691 12801
rect 36648 12764 36676 12795
rect 37642 12792 37648 12844
rect 37700 12832 37706 12844
rect 37737 12835 37795 12841
rect 37737 12832 37749 12835
rect 37700 12804 37749 12832
rect 37700 12792 37706 12804
rect 37737 12801 37749 12804
rect 37783 12801 37795 12835
rect 37737 12795 37795 12801
rect 38473 12835 38531 12841
rect 38473 12801 38485 12835
rect 38519 12832 38531 12835
rect 40402 12832 40408 12844
rect 38519 12804 40408 12832
rect 38519 12801 38531 12804
rect 38473 12795 38531 12801
rect 40402 12792 40408 12804
rect 40460 12792 40466 12844
rect 41506 12832 41512 12844
rect 41467 12804 41512 12832
rect 41506 12792 41512 12804
rect 41564 12792 41570 12844
rect 41693 12835 41751 12841
rect 41693 12801 41705 12835
rect 41739 12801 41751 12835
rect 41693 12795 41751 12801
rect 41785 12835 41843 12841
rect 41785 12801 41797 12835
rect 41831 12832 41843 12835
rect 42352 12832 42380 12872
rect 42886 12860 42892 12872
rect 42944 12860 42950 12912
rect 41831 12804 42380 12832
rect 41831 12801 41843 12804
rect 41785 12795 41843 12801
rect 37918 12764 37924 12776
rect 35912 12736 36124 12764
rect 36648 12736 37924 12764
rect 33735 12733 33747 12736
rect 33689 12727 33747 12733
rect 34422 12696 34428 12708
rect 29012 12668 33088 12696
rect 33152 12668 34428 12696
rect 29012 12628 29040 12668
rect 28368 12600 29040 12628
rect 28261 12591 28319 12597
rect 29086 12588 29092 12640
rect 29144 12628 29150 12640
rect 29733 12631 29791 12637
rect 29733 12628 29745 12631
rect 29144 12600 29745 12628
rect 29144 12588 29150 12600
rect 29733 12597 29745 12600
rect 29779 12597 29791 12631
rect 29733 12591 29791 12597
rect 30006 12588 30012 12640
rect 30064 12628 30070 12640
rect 32030 12628 32036 12640
rect 30064 12600 32036 12628
rect 30064 12588 30070 12600
rect 32030 12588 32036 12600
rect 32088 12588 32094 12640
rect 32214 12628 32220 12640
rect 32175 12600 32220 12628
rect 32214 12588 32220 12600
rect 32272 12588 32278 12640
rect 32950 12588 32956 12640
rect 33008 12628 33014 12640
rect 33152 12628 33180 12668
rect 34422 12656 34428 12668
rect 34480 12656 34486 12708
rect 35912 12696 35940 12736
rect 34624 12668 35940 12696
rect 36096 12696 36124 12736
rect 37918 12724 37924 12736
rect 37976 12724 37982 12776
rect 38010 12724 38016 12776
rect 38068 12764 38074 12776
rect 41524 12764 41552 12792
rect 38068 12736 41552 12764
rect 41708 12764 41736 12795
rect 42426 12792 42432 12844
rect 42484 12832 42490 12844
rect 42484 12804 42529 12832
rect 42484 12792 42490 12804
rect 42610 12792 42616 12844
rect 42668 12832 42674 12844
rect 43824 12832 43852 12940
rect 45646 12928 45652 12940
rect 45704 12928 45710 12980
rect 46382 12968 46388 12980
rect 46343 12940 46388 12968
rect 46382 12928 46388 12940
rect 46440 12928 46446 12980
rect 48314 12968 48320 12980
rect 48275 12940 48320 12968
rect 48314 12928 48320 12940
rect 48372 12928 48378 12980
rect 50430 12968 50436 12980
rect 49620 12940 50436 12968
rect 46661 12903 46719 12909
rect 46661 12869 46673 12903
rect 46707 12900 46719 12903
rect 47670 12900 47676 12912
rect 46707 12872 47676 12900
rect 46707 12869 46719 12872
rect 46661 12863 46719 12869
rect 47670 12860 47676 12872
rect 47728 12860 47734 12912
rect 47762 12860 47768 12912
rect 47820 12900 47826 12912
rect 47949 12903 48007 12909
rect 47949 12900 47961 12903
rect 47820 12872 47961 12900
rect 47820 12860 47826 12872
rect 47949 12869 47961 12872
rect 47995 12869 48007 12903
rect 48165 12903 48223 12909
rect 48165 12900 48177 12903
rect 47949 12863 48007 12869
rect 48056 12872 48177 12900
rect 43990 12832 43996 12844
rect 42668 12804 43852 12832
rect 43951 12804 43996 12832
rect 42668 12792 42674 12804
rect 43990 12792 43996 12804
rect 44048 12792 44054 12844
rect 44545 12835 44603 12841
rect 44545 12801 44557 12835
rect 44591 12801 44603 12835
rect 44726 12832 44732 12844
rect 44687 12804 44732 12832
rect 44545 12795 44603 12801
rect 41708 12736 42012 12764
rect 38068 12724 38074 12736
rect 41782 12696 41788 12708
rect 36096 12668 41788 12696
rect 33008 12600 33180 12628
rect 33229 12631 33287 12637
rect 33008 12588 33014 12600
rect 33229 12597 33241 12631
rect 33275 12628 33287 12631
rect 33502 12628 33508 12640
rect 33275 12600 33508 12628
rect 33275 12597 33287 12600
rect 33229 12591 33287 12597
rect 33502 12588 33508 12600
rect 33560 12588 33566 12640
rect 33870 12588 33876 12640
rect 33928 12628 33934 12640
rect 34624 12628 34652 12668
rect 41782 12656 41788 12668
rect 41840 12656 41846 12708
rect 35066 12628 35072 12640
rect 33928 12600 34652 12628
rect 35027 12600 35072 12628
rect 33928 12588 33934 12600
rect 35066 12588 35072 12600
rect 35124 12588 35130 12640
rect 36081 12631 36139 12637
rect 36081 12597 36093 12631
rect 36127 12628 36139 12631
rect 36538 12628 36544 12640
rect 36127 12600 36544 12628
rect 36127 12597 36139 12600
rect 36081 12591 36139 12597
rect 36538 12588 36544 12600
rect 36596 12588 36602 12640
rect 36630 12588 36636 12640
rect 36688 12628 36694 12640
rect 39942 12628 39948 12640
rect 36688 12600 39948 12628
rect 36688 12588 36694 12600
rect 39942 12588 39948 12600
rect 40000 12588 40006 12640
rect 40218 12588 40224 12640
rect 40276 12628 40282 12640
rect 41325 12631 41383 12637
rect 41325 12628 41337 12631
rect 40276 12600 41337 12628
rect 40276 12588 40282 12600
rect 41325 12597 41337 12600
rect 41371 12597 41383 12631
rect 41984 12628 42012 12736
rect 42978 12724 42984 12776
rect 43036 12764 43042 12776
rect 43806 12764 43812 12776
rect 43036 12736 43812 12764
rect 43036 12724 43042 12736
rect 43806 12724 43812 12736
rect 43864 12724 43870 12776
rect 43898 12724 43904 12776
rect 43956 12764 43962 12776
rect 43956 12736 44001 12764
rect 43956 12724 43962 12736
rect 44082 12724 44088 12776
rect 44140 12764 44146 12776
rect 44560 12764 44588 12795
rect 44726 12792 44732 12804
rect 44784 12792 44790 12844
rect 44818 12792 44824 12844
rect 44876 12832 44882 12844
rect 44876 12804 44921 12832
rect 44876 12792 44882 12804
rect 45646 12792 45652 12844
rect 45704 12832 45710 12844
rect 46106 12832 46112 12844
rect 45704 12804 46112 12832
rect 45704 12792 45710 12804
rect 46106 12792 46112 12804
rect 46164 12792 46170 12844
rect 46566 12832 46572 12844
rect 46527 12804 46572 12832
rect 46566 12792 46572 12804
rect 46624 12792 46630 12844
rect 46750 12832 46756 12844
rect 46711 12804 46756 12832
rect 46750 12792 46756 12804
rect 46808 12792 46814 12844
rect 46842 12792 46848 12844
rect 46900 12841 46906 12844
rect 46900 12835 46929 12841
rect 46917 12801 46929 12835
rect 47026 12832 47032 12844
rect 46987 12804 47032 12832
rect 46900 12795 46929 12801
rect 46900 12792 46906 12795
rect 47026 12792 47032 12804
rect 47084 12792 47090 12844
rect 47210 12792 47216 12844
rect 47268 12832 47274 12844
rect 48056 12832 48084 12872
rect 48165 12869 48177 12872
rect 48211 12900 48223 12903
rect 49620 12900 49648 12940
rect 50430 12928 50436 12940
rect 50488 12928 50494 12980
rect 51442 12928 51448 12980
rect 51500 12968 51506 12980
rect 52733 12971 52791 12977
rect 52733 12968 52745 12971
rect 51500 12940 52745 12968
rect 51500 12928 51506 12940
rect 52733 12937 52745 12940
rect 52779 12937 52791 12971
rect 52733 12931 52791 12937
rect 52822 12928 52828 12980
rect 52880 12968 52886 12980
rect 55950 12968 55956 12980
rect 52880 12940 55956 12968
rect 52880 12928 52886 12940
rect 55950 12928 55956 12940
rect 56008 12928 56014 12980
rect 57054 12968 57060 12980
rect 56060 12940 57060 12968
rect 48211 12872 49648 12900
rect 49697 12903 49755 12909
rect 48211 12869 48223 12872
rect 48165 12863 48223 12869
rect 49697 12869 49709 12903
rect 49743 12900 49755 12903
rect 50798 12900 50804 12912
rect 49743 12872 50804 12900
rect 49743 12869 49755 12872
rect 49697 12863 49755 12869
rect 50798 12860 50804 12872
rect 50856 12860 50862 12912
rect 51718 12903 51776 12909
rect 51718 12869 51730 12903
rect 51764 12900 51776 12903
rect 52086 12900 52092 12912
rect 51764 12872 52092 12900
rect 51764 12869 51776 12872
rect 51718 12863 51776 12869
rect 52086 12860 52092 12872
rect 52144 12860 52150 12912
rect 52178 12860 52184 12912
rect 52236 12900 52242 12912
rect 54573 12903 54631 12909
rect 54573 12900 54585 12903
rect 52236 12872 54585 12900
rect 52236 12860 52242 12872
rect 54573 12869 54585 12872
rect 54619 12900 54631 12903
rect 56060 12900 56088 12940
rect 57054 12928 57060 12940
rect 57112 12928 57118 12980
rect 57514 12968 57520 12980
rect 57164 12940 57520 12968
rect 54619 12872 56088 12900
rect 56965 12903 57023 12909
rect 54619 12869 54631 12872
rect 54573 12863 54631 12869
rect 56965 12869 56977 12903
rect 57011 12900 57023 12903
rect 57164 12900 57192 12940
rect 57514 12928 57520 12940
rect 57572 12928 57578 12980
rect 57606 12928 57612 12980
rect 57664 12968 57670 12980
rect 59078 12968 59084 12980
rect 57664 12940 59084 12968
rect 57664 12928 57670 12940
rect 59078 12928 59084 12940
rect 59136 12928 59142 12980
rect 59170 12928 59176 12980
rect 59228 12968 59234 12980
rect 59265 12971 59323 12977
rect 59265 12968 59277 12971
rect 59228 12940 59277 12968
rect 59228 12928 59234 12940
rect 59265 12937 59277 12940
rect 59311 12937 59323 12971
rect 59265 12931 59323 12937
rect 59446 12928 59452 12980
rect 59504 12968 59510 12980
rect 61010 12968 61016 12980
rect 59504 12940 61016 12968
rect 59504 12928 59510 12940
rect 61010 12928 61016 12940
rect 61068 12928 61074 12980
rect 62206 12968 62212 12980
rect 61580 12940 62212 12968
rect 59814 12900 59820 12912
rect 57011 12872 57192 12900
rect 57532 12872 59820 12900
rect 57011 12869 57023 12872
rect 56965 12863 57023 12869
rect 57532 12844 57560 12872
rect 59814 12860 59820 12872
rect 59872 12860 59878 12912
rect 60550 12860 60556 12912
rect 60608 12900 60614 12912
rect 61580 12909 61608 12940
rect 62206 12928 62212 12940
rect 62264 12928 62270 12980
rect 63494 12968 63500 12980
rect 62408 12940 63500 12968
rect 61565 12903 61623 12909
rect 61565 12900 61577 12903
rect 60608 12872 61577 12900
rect 60608 12860 60614 12872
rect 61565 12869 61577 12872
rect 61611 12869 61623 12903
rect 61565 12863 61623 12869
rect 61838 12860 61844 12912
rect 61896 12900 61902 12912
rect 62301 12903 62359 12909
rect 62301 12900 62313 12903
rect 61896 12872 62313 12900
rect 61896 12860 61902 12872
rect 62301 12869 62313 12872
rect 62347 12869 62359 12903
rect 62301 12863 62359 12869
rect 47268 12804 48084 12832
rect 48777 12835 48835 12841
rect 47268 12792 47274 12804
rect 48777 12801 48789 12835
rect 48823 12832 48835 12835
rect 49142 12832 49148 12844
rect 48823 12804 49148 12832
rect 48823 12801 48835 12804
rect 48777 12795 48835 12801
rect 49142 12792 49148 12804
rect 49200 12832 49206 12844
rect 49602 12832 49608 12844
rect 49200 12804 49608 12832
rect 49200 12792 49206 12804
rect 49602 12792 49608 12804
rect 49660 12792 49666 12844
rect 50982 12792 50988 12844
rect 51040 12832 51046 12844
rect 51445 12835 51503 12841
rect 51445 12832 51457 12835
rect 51040 12822 51074 12832
rect 51184 12822 51457 12832
rect 51040 12804 51457 12822
rect 51040 12794 51212 12804
rect 51445 12801 51457 12804
rect 51491 12801 51503 12835
rect 51445 12795 51503 12801
rect 51629 12835 51687 12841
rect 51629 12801 51641 12835
rect 51675 12801 51687 12835
rect 51810 12832 51816 12844
rect 51769 12804 51816 12832
rect 51629 12795 51687 12801
rect 51040 12792 51046 12794
rect 45278 12764 45284 12776
rect 44140 12736 44185 12764
rect 44560 12736 45284 12764
rect 44140 12724 44146 12736
rect 45278 12724 45284 12736
rect 45336 12724 45342 12776
rect 45462 12724 45468 12776
rect 45520 12764 45526 12776
rect 45558 12767 45616 12773
rect 45558 12764 45570 12767
rect 45520 12736 45570 12764
rect 45520 12724 45526 12736
rect 45558 12733 45570 12736
rect 45604 12733 45616 12767
rect 45738 12764 45744 12776
rect 45699 12736 45744 12764
rect 45558 12727 45616 12733
rect 45738 12724 45744 12736
rect 45796 12724 45802 12776
rect 45833 12767 45891 12773
rect 45833 12733 45845 12767
rect 45879 12764 45891 12767
rect 46014 12764 46020 12776
rect 45879 12736 46020 12764
rect 45879 12733 45891 12736
rect 45833 12727 45891 12733
rect 46014 12724 46020 12736
rect 46072 12724 46078 12776
rect 48038 12724 48044 12776
rect 48096 12764 48102 12776
rect 49881 12767 49939 12773
rect 49881 12764 49893 12767
rect 48096 12736 49893 12764
rect 48096 12724 48102 12736
rect 49881 12733 49893 12736
rect 49927 12764 49939 12767
rect 49973 12767 50031 12773
rect 49973 12764 49985 12767
rect 49927 12736 49985 12764
rect 49927 12733 49939 12736
rect 49881 12727 49939 12733
rect 49973 12733 49985 12736
rect 50019 12733 50031 12767
rect 49973 12727 50031 12733
rect 50154 12724 50160 12776
rect 50212 12764 50218 12776
rect 50249 12767 50307 12773
rect 50249 12764 50261 12767
rect 50212 12736 50261 12764
rect 50212 12724 50218 12736
rect 50249 12733 50261 12736
rect 50295 12733 50307 12767
rect 50249 12727 50307 12733
rect 50430 12724 50436 12776
rect 50488 12764 50494 12776
rect 50798 12764 50804 12776
rect 50488 12736 50804 12764
rect 50488 12724 50494 12736
rect 50798 12724 50804 12736
rect 50856 12724 50862 12776
rect 51644 12764 51672 12795
rect 51810 12792 51816 12804
rect 51868 12841 51874 12844
rect 51868 12835 51917 12841
rect 51868 12801 51871 12835
rect 51905 12832 51917 12835
rect 52270 12832 52276 12844
rect 51905 12804 52276 12832
rect 51905 12801 51917 12804
rect 51868 12795 51917 12801
rect 51868 12792 51874 12795
rect 52270 12792 52276 12804
rect 52328 12792 52334 12844
rect 52822 12792 52828 12844
rect 52880 12832 52886 12844
rect 52917 12835 52975 12841
rect 52917 12832 52929 12835
rect 52880 12804 52929 12832
rect 52880 12792 52886 12804
rect 52917 12801 52929 12804
rect 52963 12801 52975 12835
rect 53098 12832 53104 12844
rect 53059 12804 53104 12832
rect 52917 12795 52975 12801
rect 53098 12792 53104 12804
rect 53156 12792 53162 12844
rect 53190 12792 53196 12844
rect 53248 12832 53254 12844
rect 53561 12835 53619 12841
rect 53248 12804 53293 12832
rect 53248 12792 53254 12804
rect 53561 12801 53573 12835
rect 53607 12832 53619 12835
rect 53650 12832 53656 12844
rect 53607 12804 53656 12832
rect 53607 12801 53619 12804
rect 53561 12795 53619 12801
rect 53650 12792 53656 12804
rect 53708 12792 53714 12844
rect 53745 12835 53803 12841
rect 53745 12801 53757 12835
rect 53791 12801 53803 12835
rect 53745 12795 53803 12801
rect 52730 12764 52736 12776
rect 51644 12736 52736 12764
rect 52730 12724 52736 12736
rect 52788 12724 52794 12776
rect 53282 12724 53288 12776
rect 53340 12764 53346 12776
rect 53760 12764 53788 12795
rect 53834 12792 53840 12844
rect 53892 12832 53898 12844
rect 53892 12804 53937 12832
rect 53892 12792 53898 12804
rect 54478 12792 54484 12844
rect 54536 12832 54542 12844
rect 55306 12832 55312 12844
rect 54536 12804 55312 12832
rect 54536 12792 54542 12804
rect 55306 12792 55312 12804
rect 55364 12792 55370 12844
rect 55674 12792 55680 12844
rect 55732 12832 55738 12844
rect 56410 12832 56416 12844
rect 55732 12804 56416 12832
rect 55732 12792 55738 12804
rect 56410 12792 56416 12804
rect 56468 12792 56474 12844
rect 56686 12832 56692 12844
rect 56647 12804 56692 12832
rect 56686 12792 56692 12804
rect 56744 12792 56750 12844
rect 56778 12792 56784 12844
rect 56836 12841 56842 12844
rect 56836 12835 56885 12841
rect 56836 12801 56839 12835
rect 56873 12801 56885 12835
rect 56836 12795 56885 12801
rect 57057 12835 57115 12841
rect 57057 12801 57069 12835
rect 57103 12801 57115 12835
rect 57057 12795 57115 12801
rect 57164 12804 57468 12832
rect 56836 12792 56842 12795
rect 53340 12736 53788 12764
rect 53340 12724 53346 12736
rect 54570 12724 54576 12776
rect 54628 12764 54634 12776
rect 56134 12764 56140 12776
rect 54628 12736 56140 12764
rect 54628 12724 54634 12736
rect 56134 12724 56140 12736
rect 56192 12724 56198 12776
rect 56962 12724 56968 12776
rect 57020 12764 57026 12776
rect 57072 12764 57100 12795
rect 57020 12736 57100 12764
rect 57020 12724 57026 12736
rect 43625 12699 43683 12705
rect 43625 12665 43637 12699
rect 43671 12696 43683 12699
rect 50890 12696 50896 12708
rect 43671 12668 48452 12696
rect 43671 12665 43683 12668
rect 43625 12659 43683 12665
rect 42242 12628 42248 12640
rect 41984 12600 42248 12628
rect 41325 12591 41383 12597
rect 42242 12588 42248 12600
rect 42300 12588 42306 12640
rect 43714 12588 43720 12640
rect 43772 12628 43778 12640
rect 43898 12628 43904 12640
rect 43772 12600 43904 12628
rect 43772 12588 43778 12600
rect 43898 12588 43904 12600
rect 43956 12588 43962 12640
rect 44545 12631 44603 12637
rect 44545 12597 44557 12631
rect 44591 12628 44603 12631
rect 44634 12628 44640 12640
rect 44591 12600 44640 12628
rect 44591 12597 44603 12600
rect 44545 12591 44603 12597
rect 44634 12588 44640 12600
rect 44692 12588 44698 12640
rect 45373 12631 45431 12637
rect 45373 12597 45385 12631
rect 45419 12628 45431 12631
rect 45554 12628 45560 12640
rect 45419 12600 45560 12628
rect 45419 12597 45431 12600
rect 45373 12591 45431 12597
rect 45554 12588 45560 12600
rect 45612 12588 45618 12640
rect 45922 12588 45928 12640
rect 45980 12628 45986 12640
rect 48038 12628 48044 12640
rect 45980 12600 48044 12628
rect 45980 12588 45986 12600
rect 48038 12588 48044 12600
rect 48096 12588 48102 12640
rect 48130 12588 48136 12640
rect 48188 12628 48194 12640
rect 48424 12628 48452 12668
rect 48700 12668 50896 12696
rect 48700 12628 48728 12668
rect 50890 12656 50896 12668
rect 50948 12656 50954 12708
rect 51169 12699 51227 12705
rect 51169 12665 51181 12699
rect 51215 12696 51227 12699
rect 51810 12696 51816 12708
rect 51215 12668 51816 12696
rect 51215 12665 51227 12668
rect 51169 12659 51227 12665
rect 51810 12656 51816 12668
rect 51868 12656 51874 12708
rect 52362 12656 52368 12708
rect 52420 12696 52426 12708
rect 57164 12696 57192 12804
rect 57330 12764 57336 12776
rect 57256 12736 57336 12764
rect 57256 12705 57284 12736
rect 57330 12724 57336 12736
rect 57388 12724 57394 12776
rect 57440 12764 57468 12804
rect 57514 12792 57520 12844
rect 57572 12792 57578 12844
rect 57606 12792 57612 12844
rect 57664 12832 57670 12844
rect 57885 12835 57943 12841
rect 57885 12832 57897 12835
rect 57664 12804 57897 12832
rect 57664 12792 57670 12804
rect 57885 12801 57897 12804
rect 57931 12801 57943 12835
rect 57885 12795 57943 12801
rect 57974 12792 57980 12844
rect 58032 12832 58038 12844
rect 58710 12832 58716 12844
rect 58032 12804 58716 12832
rect 58032 12792 58038 12804
rect 58710 12792 58716 12804
rect 58768 12832 58774 12844
rect 59081 12835 59139 12841
rect 59081 12832 59093 12835
rect 58768 12804 59093 12832
rect 58768 12792 58774 12804
rect 59081 12801 59093 12804
rect 59127 12801 59139 12835
rect 59081 12795 59139 12801
rect 59357 12835 59415 12841
rect 59357 12801 59369 12835
rect 59403 12801 59415 12835
rect 59357 12795 59415 12801
rect 57440 12736 57974 12764
rect 52420 12668 57192 12696
rect 57241 12699 57299 12705
rect 52420 12656 52426 12668
rect 57241 12665 57253 12699
rect 57287 12665 57299 12699
rect 57946 12696 57974 12736
rect 58066 12724 58072 12776
rect 58124 12764 58130 12776
rect 58161 12767 58219 12773
rect 58161 12764 58173 12767
rect 58124 12736 58173 12764
rect 58124 12724 58130 12736
rect 58161 12733 58173 12736
rect 58207 12733 58219 12767
rect 59372 12764 59400 12795
rect 60642 12792 60648 12844
rect 60700 12832 60706 12844
rect 62408 12841 62436 12940
rect 63494 12928 63500 12940
rect 63552 12928 63558 12980
rect 63954 12928 63960 12980
rect 64012 12968 64018 12980
rect 64877 12971 64935 12977
rect 64012 12940 64828 12968
rect 64012 12928 64018 12940
rect 63304 12903 63362 12909
rect 63304 12869 63316 12903
rect 63350 12900 63362 12903
rect 64598 12900 64604 12912
rect 63350 12872 64604 12900
rect 63350 12869 63362 12872
rect 63304 12863 63362 12869
rect 64598 12860 64604 12872
rect 64656 12860 64662 12912
rect 64800 12900 64828 12940
rect 64877 12937 64889 12971
rect 64923 12968 64935 12971
rect 65058 12968 65064 12980
rect 64923 12940 65064 12968
rect 64923 12937 64935 12940
rect 64877 12931 64935 12937
rect 65058 12928 65064 12940
rect 65116 12928 65122 12980
rect 66346 12928 66352 12980
rect 66404 12968 66410 12980
rect 68370 12968 68376 12980
rect 66404 12940 68376 12968
rect 66404 12928 66410 12940
rect 68370 12928 68376 12940
rect 68428 12928 68434 12980
rect 70026 12968 70032 12980
rect 69032 12940 70032 12968
rect 66441 12903 66499 12909
rect 64800 12872 65472 12900
rect 61933 12835 61991 12841
rect 61933 12832 61945 12835
rect 60700 12804 61945 12832
rect 60700 12792 60706 12804
rect 61933 12801 61945 12804
rect 61979 12801 61991 12835
rect 61933 12795 61991 12801
rect 62117 12835 62175 12841
rect 62117 12801 62129 12835
rect 62163 12801 62175 12835
rect 62117 12795 62175 12801
rect 62393 12835 62451 12841
rect 62393 12801 62405 12835
rect 62439 12801 62451 12835
rect 62393 12795 62451 12801
rect 58161 12727 58219 12733
rect 58268 12736 59400 12764
rect 58268 12696 58296 12736
rect 59446 12724 59452 12776
rect 59504 12764 59510 12776
rect 62132 12764 62160 12795
rect 62666 12792 62672 12844
rect 62724 12832 62730 12844
rect 65150 12832 65156 12844
rect 62724 12804 65156 12832
rect 62724 12792 62730 12804
rect 65150 12792 65156 12804
rect 65208 12792 65214 12844
rect 65334 12832 65340 12844
rect 65247 12804 65340 12832
rect 63034 12764 63040 12776
rect 59504 12736 62160 12764
rect 62995 12736 63040 12764
rect 59504 12724 59510 12736
rect 63034 12724 63040 12736
rect 63092 12724 63098 12776
rect 64046 12724 64052 12776
rect 64104 12764 64110 12776
rect 65061 12767 65119 12773
rect 65061 12764 65073 12767
rect 64104 12736 65073 12764
rect 64104 12724 64110 12736
rect 65061 12733 65073 12736
rect 65107 12733 65119 12767
rect 65260 12764 65288 12804
rect 65334 12792 65340 12804
rect 65392 12792 65398 12844
rect 65061 12727 65119 12733
rect 65168 12736 65288 12764
rect 65444 12764 65472 12872
rect 66441 12869 66453 12903
rect 66487 12900 66499 12903
rect 67177 12903 67235 12909
rect 67177 12900 67189 12903
rect 66487 12872 67189 12900
rect 66487 12869 66499 12872
rect 66441 12863 66499 12869
rect 67177 12869 67189 12872
rect 67223 12869 67235 12903
rect 67177 12863 67235 12869
rect 67545 12903 67603 12909
rect 67545 12869 67557 12903
rect 67591 12900 67603 12903
rect 67910 12900 67916 12912
rect 67591 12872 67916 12900
rect 67591 12869 67603 12872
rect 67545 12863 67603 12869
rect 67910 12860 67916 12872
rect 67968 12860 67974 12912
rect 68922 12900 68928 12912
rect 68664 12872 68928 12900
rect 66254 12832 66260 12844
rect 66215 12804 66260 12832
rect 66254 12792 66260 12804
rect 66312 12792 66318 12844
rect 66346 12792 66352 12844
rect 66404 12832 66410 12844
rect 66533 12835 66591 12841
rect 66533 12832 66545 12835
rect 66404 12804 66545 12832
rect 66404 12792 66410 12804
rect 66533 12801 66545 12804
rect 66579 12801 66591 12835
rect 66533 12795 66591 12801
rect 66625 12835 66683 12841
rect 66625 12801 66637 12835
rect 66671 12801 66683 12835
rect 66625 12795 66683 12801
rect 66640 12764 66668 12795
rect 66714 12792 66720 12844
rect 66772 12832 66778 12844
rect 67361 12835 67419 12841
rect 67361 12832 67373 12835
rect 66772 12804 67373 12832
rect 66772 12792 66778 12804
rect 67361 12801 67373 12804
rect 67407 12801 67419 12835
rect 67361 12795 67419 12801
rect 65444 12736 66668 12764
rect 67376 12764 67404 12795
rect 67450 12792 67456 12844
rect 67508 12832 67514 12844
rect 67637 12835 67695 12841
rect 67637 12832 67649 12835
rect 67508 12804 67649 12832
rect 67508 12792 67514 12804
rect 67637 12801 67649 12804
rect 67683 12832 67695 12835
rect 68664 12832 68692 12872
rect 68922 12860 68928 12872
rect 68980 12860 68986 12912
rect 67683 12804 68692 12832
rect 68741 12835 68799 12841
rect 67683 12801 67695 12804
rect 67637 12795 67695 12801
rect 68741 12801 68753 12835
rect 68787 12832 68799 12835
rect 69032 12832 69060 12940
rect 70026 12928 70032 12940
rect 70084 12928 70090 12980
rect 86770 12968 86776 12980
rect 86731 12940 86776 12968
rect 86770 12928 86776 12940
rect 86828 12928 86834 12980
rect 69216 12872 70256 12900
rect 68787 12804 69060 12832
rect 68787 12801 68799 12804
rect 68741 12795 68799 12801
rect 69106 12792 69112 12844
rect 69164 12832 69170 12844
rect 69216 12841 69244 12872
rect 69201 12835 69259 12841
rect 69201 12832 69213 12835
rect 69164 12804 69213 12832
rect 69164 12792 69170 12804
rect 69201 12801 69213 12804
rect 69247 12801 69259 12835
rect 69201 12795 69259 12801
rect 69293 12835 69351 12841
rect 69293 12801 69305 12835
rect 69339 12832 69351 12835
rect 69382 12832 69388 12844
rect 69339 12804 69388 12832
rect 69339 12801 69351 12804
rect 69293 12795 69351 12801
rect 69382 12792 69388 12804
rect 69440 12792 69446 12844
rect 69474 12792 69480 12844
rect 69532 12832 69538 12844
rect 69532 12804 69577 12832
rect 69532 12792 69538 12804
rect 69750 12792 69756 12844
rect 69808 12832 69814 12844
rect 70112 12836 70170 12841
rect 70044 12835 70170 12836
rect 70044 12832 70124 12835
rect 69808 12808 70124 12832
rect 69808 12804 70072 12808
rect 69808 12792 69814 12804
rect 70112 12801 70124 12808
rect 70158 12801 70170 12835
rect 70228 12832 70256 12872
rect 70302 12860 70308 12912
rect 70360 12900 70366 12912
rect 88150 12900 88156 12912
rect 70360 12872 88156 12900
rect 70360 12860 70366 12872
rect 88150 12860 88156 12872
rect 88208 12860 88214 12912
rect 71593 12835 71651 12841
rect 71593 12832 71605 12835
rect 70228 12804 71605 12832
rect 70112 12795 70170 12801
rect 71593 12801 71605 12804
rect 71639 12801 71651 12835
rect 71593 12795 71651 12801
rect 71682 12792 71688 12844
rect 71740 12832 71746 12844
rect 71777 12835 71835 12841
rect 71777 12832 71789 12835
rect 71740 12804 71789 12832
rect 71740 12792 71746 12804
rect 71777 12801 71789 12804
rect 71823 12832 71835 12835
rect 71866 12832 71872 12844
rect 71823 12804 71872 12832
rect 71823 12801 71835 12804
rect 71777 12795 71835 12801
rect 71866 12792 71872 12804
rect 71924 12792 71930 12844
rect 72326 12832 72332 12844
rect 72287 12804 72332 12832
rect 72326 12792 72332 12804
rect 72384 12792 72390 12844
rect 86954 12832 86960 12844
rect 86915 12804 86960 12832
rect 86954 12792 86960 12804
rect 87012 12792 87018 12844
rect 87046 12792 87052 12844
rect 87104 12832 87110 12844
rect 88245 12835 88303 12841
rect 88245 12832 88257 12835
rect 87104 12804 88257 12832
rect 87104 12792 87110 12804
rect 88245 12801 88257 12804
rect 88291 12801 88303 12835
rect 88245 12795 88303 12801
rect 69658 12764 69664 12776
rect 67376 12736 69664 12764
rect 57946 12668 58296 12696
rect 59081 12699 59139 12705
rect 57241 12659 57299 12665
rect 59081 12665 59093 12699
rect 59127 12696 59139 12699
rect 60458 12696 60464 12708
rect 59127 12668 60464 12696
rect 59127 12665 59139 12668
rect 59081 12659 59139 12665
rect 60458 12656 60464 12668
rect 60516 12656 60522 12708
rect 60642 12656 60648 12708
rect 60700 12696 60706 12708
rect 60700 12668 61139 12696
rect 60700 12656 60706 12668
rect 48866 12628 48872 12640
rect 48188 12600 48233 12628
rect 48424 12600 48728 12628
rect 48827 12600 48872 12628
rect 48188 12588 48194 12600
rect 48866 12588 48872 12600
rect 48924 12588 48930 12640
rect 50614 12588 50620 12640
rect 50672 12628 50678 12640
rect 51997 12631 52055 12637
rect 51997 12628 52009 12631
rect 50672 12600 52009 12628
rect 50672 12588 50678 12600
rect 51997 12597 52009 12600
rect 52043 12597 52055 12631
rect 51997 12591 52055 12597
rect 52546 12588 52552 12640
rect 52604 12628 52610 12640
rect 53561 12631 53619 12637
rect 53561 12628 53573 12631
rect 52604 12600 53573 12628
rect 52604 12588 52610 12600
rect 53561 12597 53573 12600
rect 53607 12597 53619 12631
rect 53561 12591 53619 12597
rect 54386 12588 54392 12640
rect 54444 12628 54450 12640
rect 55306 12628 55312 12640
rect 54444 12600 55312 12628
rect 54444 12588 54450 12600
rect 55306 12588 55312 12600
rect 55364 12588 55370 12640
rect 55582 12588 55588 12640
rect 55640 12628 55646 12640
rect 55861 12631 55919 12637
rect 55861 12628 55873 12631
rect 55640 12600 55873 12628
rect 55640 12588 55646 12600
rect 55861 12597 55873 12600
rect 55907 12597 55919 12631
rect 55861 12591 55919 12597
rect 55950 12588 55956 12640
rect 56008 12628 56014 12640
rect 59998 12628 60004 12640
rect 56008 12600 60004 12628
rect 56008 12588 56014 12600
rect 59998 12588 60004 12600
rect 60056 12588 60062 12640
rect 60090 12588 60096 12640
rect 60148 12628 60154 12640
rect 61010 12628 61016 12640
rect 60148 12600 61016 12628
rect 60148 12588 60154 12600
rect 61010 12588 61016 12600
rect 61068 12588 61074 12640
rect 61111 12628 61139 12668
rect 64506 12656 64512 12708
rect 64564 12696 64570 12708
rect 65168 12696 65196 12736
rect 69658 12724 69664 12736
rect 69716 12724 69722 12776
rect 69842 12764 69848 12776
rect 69803 12736 69848 12764
rect 69842 12724 69848 12736
rect 69900 12724 69906 12776
rect 64564 12668 65196 12696
rect 65245 12699 65303 12705
rect 64564 12656 64570 12668
rect 65245 12665 65257 12699
rect 65291 12696 65303 12699
rect 68557 12699 68615 12705
rect 65291 12668 68508 12696
rect 65291 12665 65303 12668
rect 65245 12659 65303 12665
rect 64417 12631 64475 12637
rect 64417 12628 64429 12631
rect 61111 12600 64429 12628
rect 64417 12597 64429 12600
rect 64463 12597 64475 12631
rect 64417 12591 64475 12597
rect 66254 12588 66260 12640
rect 66312 12628 66318 12640
rect 66809 12631 66867 12637
rect 66809 12628 66821 12631
rect 66312 12600 66821 12628
rect 66312 12588 66318 12600
rect 66809 12597 66821 12600
rect 66855 12597 66867 12631
rect 68480 12628 68508 12668
rect 68557 12665 68569 12699
rect 68603 12696 68615 12699
rect 69750 12696 69756 12708
rect 68603 12668 69756 12696
rect 68603 12665 68615 12668
rect 68557 12659 68615 12665
rect 69750 12656 69756 12668
rect 69808 12656 69814 12708
rect 71961 12699 72019 12705
rect 71961 12696 71973 12699
rect 70780 12668 71973 12696
rect 69290 12628 69296 12640
rect 68480 12600 69296 12628
rect 66809 12591 66867 12597
rect 69290 12588 69296 12600
rect 69348 12588 69354 12640
rect 70026 12588 70032 12640
rect 70084 12628 70090 12640
rect 70780 12628 70808 12668
rect 71961 12665 71973 12668
rect 72007 12665 72019 12699
rect 71961 12659 72019 12665
rect 70084 12600 70808 12628
rect 71225 12631 71283 12637
rect 70084 12588 70090 12600
rect 71225 12597 71237 12631
rect 71271 12628 71283 12631
rect 71774 12628 71780 12640
rect 71271 12600 71780 12628
rect 71271 12597 71283 12600
rect 71225 12591 71283 12597
rect 71774 12588 71780 12600
rect 71832 12588 71838 12640
rect 72418 12628 72424 12640
rect 72379 12600 72424 12628
rect 72418 12588 72424 12600
rect 72476 12588 72482 12640
rect 88058 12628 88064 12640
rect 88019 12600 88064 12628
rect 88058 12588 88064 12600
rect 88116 12588 88122 12640
rect 1104 12538 88872 12560
rect 1104 12486 11924 12538
rect 11976 12486 11988 12538
rect 12040 12486 12052 12538
rect 12104 12486 12116 12538
rect 12168 12486 12180 12538
rect 12232 12486 33872 12538
rect 33924 12486 33936 12538
rect 33988 12486 34000 12538
rect 34052 12486 34064 12538
rect 34116 12486 34128 12538
rect 34180 12486 55820 12538
rect 55872 12486 55884 12538
rect 55936 12486 55948 12538
rect 56000 12486 56012 12538
rect 56064 12486 56076 12538
rect 56128 12486 77768 12538
rect 77820 12486 77832 12538
rect 77884 12486 77896 12538
rect 77948 12486 77960 12538
rect 78012 12486 78024 12538
rect 78076 12486 88872 12538
rect 1104 12464 88872 12486
rect 20070 12424 20076 12436
rect 20031 12396 20076 12424
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 20220 12396 21312 12424
rect 20220 12384 20226 12396
rect 18966 12316 18972 12368
rect 19024 12356 19030 12368
rect 20993 12359 21051 12365
rect 19024 12328 20944 12356
rect 19024 12316 19030 12328
rect 20806 12288 20812 12300
rect 20767 12260 20812 12288
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 20916 12288 20944 12328
rect 20993 12325 21005 12359
rect 21039 12356 21051 12359
rect 21082 12356 21088 12368
rect 21039 12328 21088 12356
rect 21039 12325 21051 12328
rect 20993 12319 21051 12325
rect 21082 12316 21088 12328
rect 21140 12316 21146 12368
rect 21284 12356 21312 12396
rect 21358 12384 21364 12436
rect 21416 12424 21422 12436
rect 25130 12424 25136 12436
rect 21416 12396 25136 12424
rect 21416 12384 21422 12396
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 25222 12384 25228 12436
rect 25280 12424 25286 12436
rect 25777 12427 25835 12433
rect 25777 12424 25789 12427
rect 25280 12396 25789 12424
rect 25280 12384 25286 12396
rect 25777 12393 25789 12396
rect 25823 12393 25835 12427
rect 26237 12427 26295 12433
rect 25777 12387 25835 12393
rect 25884 12396 26065 12424
rect 25884 12356 25912 12396
rect 21284 12328 25912 12356
rect 26037 12356 26065 12396
rect 26237 12393 26249 12427
rect 26283 12424 26295 12427
rect 27798 12424 27804 12436
rect 26283 12396 27804 12424
rect 26283 12393 26295 12396
rect 26237 12387 26295 12393
rect 27798 12384 27804 12396
rect 27856 12384 27862 12436
rect 28534 12384 28540 12436
rect 28592 12424 28598 12436
rect 28629 12427 28687 12433
rect 28629 12424 28641 12427
rect 28592 12396 28641 12424
rect 28592 12384 28598 12396
rect 28629 12393 28641 12396
rect 28675 12393 28687 12427
rect 28629 12387 28687 12393
rect 28810 12384 28816 12436
rect 28868 12424 28874 12436
rect 30926 12424 30932 12436
rect 28868 12396 29408 12424
rect 30887 12396 30932 12424
rect 28868 12384 28874 12396
rect 26789 12359 26847 12365
rect 26789 12356 26801 12359
rect 26037 12328 26801 12356
rect 26789 12325 26801 12328
rect 26835 12356 26847 12359
rect 28258 12356 28264 12368
rect 26835 12328 26985 12356
rect 26835 12325 26847 12328
rect 26789 12319 26847 12325
rect 24946 12288 24952 12300
rect 20916 12260 24952 12288
rect 24946 12248 24952 12260
rect 25004 12248 25010 12300
rect 26050 12288 26056 12300
rect 26011 12260 26056 12288
rect 26050 12248 26056 12260
rect 26108 12248 26114 12300
rect 26957 12288 26985 12328
rect 28092 12328 28264 12356
rect 27617 12291 27675 12297
rect 27617 12288 27629 12291
rect 26957 12260 27629 12288
rect 27617 12257 27629 12260
rect 27663 12257 27675 12291
rect 27617 12251 27675 12257
rect 27801 12291 27859 12297
rect 27801 12257 27813 12291
rect 27847 12288 27859 12291
rect 28092 12288 28120 12328
rect 28258 12316 28264 12328
rect 28316 12316 28322 12368
rect 28353 12359 28411 12365
rect 28353 12325 28365 12359
rect 28399 12356 28411 12359
rect 28905 12359 28963 12365
rect 28399 12328 28580 12356
rect 28399 12325 28411 12328
rect 28353 12319 28411 12325
rect 27847 12260 28120 12288
rect 28445 12291 28503 12297
rect 27847 12257 27859 12260
rect 27801 12251 27859 12257
rect 28445 12257 28457 12291
rect 28491 12257 28503 12291
rect 28445 12251 28503 12257
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12220 19947 12223
rect 20714 12220 20720 12232
rect 19935 12192 20720 12220
rect 19935 12189 19947 12192
rect 19889 12183 19947 12189
rect 20714 12180 20720 12192
rect 20772 12180 20778 12232
rect 20990 12220 20996 12232
rect 20951 12192 20996 12220
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 21082 12180 21088 12232
rect 21140 12220 21146 12232
rect 21269 12223 21327 12229
rect 21140 12192 21185 12220
rect 21140 12180 21146 12192
rect 21269 12189 21281 12223
rect 21315 12220 21327 12223
rect 21542 12220 21548 12232
rect 21315 12192 21548 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 23474 12180 23480 12232
rect 23532 12220 23538 12232
rect 25222 12229 25228 12232
rect 25179 12223 25228 12229
rect 25179 12220 25191 12223
rect 23532 12192 25191 12220
rect 23532 12180 23538 12192
rect 25179 12189 25191 12192
rect 25225 12189 25228 12223
rect 25179 12183 25228 12189
rect 25222 12180 25228 12183
rect 25280 12180 25286 12232
rect 25419 12223 25477 12229
rect 25419 12189 25431 12223
rect 25465 12220 25477 12223
rect 26142 12220 26148 12232
rect 25465 12192 25544 12220
rect 26103 12192 26148 12220
rect 25465 12189 25477 12192
rect 25419 12183 25477 12189
rect 20901 12155 20959 12161
rect 20901 12152 20913 12155
rect 20364 12124 20913 12152
rect 1670 12044 1676 12096
rect 1728 12084 1734 12096
rect 20162 12084 20168 12096
rect 1728 12056 20168 12084
rect 1728 12044 1734 12056
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 20364 12093 20392 12124
rect 20901 12121 20913 12124
rect 20947 12121 20959 12155
rect 20901 12115 20959 12121
rect 24394 12112 24400 12164
rect 24452 12152 24458 12164
rect 25516 12152 25544 12192
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 26326 12220 26332 12232
rect 26287 12192 26332 12220
rect 26326 12180 26332 12192
rect 26384 12180 26390 12232
rect 26513 12223 26571 12229
rect 26513 12189 26525 12223
rect 26559 12220 26571 12223
rect 26786 12220 26792 12232
rect 26559 12192 26792 12220
rect 26559 12189 26571 12192
rect 26513 12183 26571 12189
rect 26786 12180 26792 12192
rect 26844 12180 26850 12232
rect 28184 12214 28304 12220
rect 28460 12214 28488 12251
rect 28552 12229 28580 12328
rect 28905 12325 28917 12359
rect 28951 12356 28963 12359
rect 28951 12328 29316 12356
rect 28951 12325 28963 12328
rect 28905 12319 28963 12325
rect 28184 12192 28488 12214
rect 27525 12155 27583 12161
rect 27525 12152 27537 12155
rect 24452 12124 27537 12152
rect 24452 12112 24458 12124
rect 27525 12121 27537 12124
rect 27571 12152 27583 12155
rect 27614 12152 27620 12164
rect 27571 12124 27620 12152
rect 27571 12121 27583 12124
rect 27525 12115 27583 12121
rect 27614 12112 27620 12124
rect 27672 12112 27678 12164
rect 27985 12155 28043 12161
rect 27985 12121 27997 12155
rect 28031 12152 28043 12155
rect 28074 12152 28080 12164
rect 28031 12124 28080 12152
rect 28031 12121 28043 12124
rect 27985 12115 28043 12121
rect 28074 12112 28080 12124
rect 28132 12112 28138 12164
rect 20349 12087 20407 12093
rect 20349 12053 20361 12087
rect 20395 12053 20407 12087
rect 20349 12047 20407 12053
rect 20530 12044 20536 12096
rect 20588 12084 20594 12096
rect 21542 12084 21548 12096
rect 20588 12056 21548 12084
rect 20588 12044 20594 12056
rect 21542 12044 21548 12056
rect 21600 12044 21606 12096
rect 24946 12084 24952 12096
rect 24907 12056 24952 12084
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 25038 12044 25044 12096
rect 25096 12084 25102 12096
rect 25317 12087 25375 12093
rect 25317 12084 25329 12087
rect 25096 12056 25329 12084
rect 25096 12044 25102 12056
rect 25317 12053 25329 12056
rect 25363 12053 25375 12087
rect 27154 12084 27160 12096
rect 27115 12056 27160 12084
rect 25317 12047 25375 12053
rect 27154 12044 27160 12056
rect 27212 12044 27218 12096
rect 27246 12044 27252 12096
rect 27304 12084 27310 12096
rect 28184 12084 28212 12192
rect 28276 12186 28488 12192
rect 28537 12223 28595 12229
rect 28537 12189 28549 12223
rect 28583 12220 28595 12223
rect 28626 12220 28632 12232
rect 28583 12192 28632 12220
rect 28583 12189 28595 12192
rect 28537 12183 28595 12189
rect 28626 12180 28632 12192
rect 28684 12180 28690 12232
rect 29086 12220 29092 12232
rect 29047 12192 29092 12220
rect 29086 12180 29092 12192
rect 29144 12180 29150 12232
rect 29288 12152 29316 12328
rect 29380 12220 29408 12396
rect 30926 12384 30932 12396
rect 30984 12384 30990 12436
rect 31570 12424 31576 12436
rect 31531 12396 31576 12424
rect 31570 12384 31576 12396
rect 31628 12384 31634 12436
rect 33042 12384 33048 12436
rect 33100 12424 33106 12436
rect 33873 12427 33931 12433
rect 33873 12424 33885 12427
rect 33100 12396 33885 12424
rect 33100 12384 33106 12396
rect 33873 12393 33885 12396
rect 33919 12393 33931 12427
rect 33873 12387 33931 12393
rect 34514 12384 34520 12436
rect 34572 12424 34578 12436
rect 35802 12424 35808 12436
rect 34572 12396 35808 12424
rect 34572 12384 34578 12396
rect 35802 12384 35808 12396
rect 35860 12384 35866 12436
rect 35986 12424 35992 12436
rect 35947 12396 35992 12424
rect 35986 12384 35992 12396
rect 36044 12384 36050 12436
rect 36170 12384 36176 12436
rect 36228 12424 36234 12436
rect 36228 12396 39344 12424
rect 36228 12384 36234 12396
rect 32122 12316 32128 12368
rect 32180 12356 32186 12368
rect 32180 12328 32352 12356
rect 32180 12316 32186 12328
rect 29546 12288 29552 12300
rect 29507 12260 29552 12288
rect 29546 12248 29552 12260
rect 29604 12248 29610 12300
rect 32214 12288 32220 12300
rect 30576 12260 32220 12288
rect 30576 12220 30604 12260
rect 32214 12248 32220 12260
rect 32272 12248 32278 12300
rect 32324 12297 32352 12328
rect 32858 12316 32864 12368
rect 32916 12356 32922 12368
rect 34793 12359 34851 12365
rect 32916 12328 34284 12356
rect 32916 12316 32922 12328
rect 32309 12291 32367 12297
rect 32309 12257 32321 12291
rect 32355 12257 32367 12291
rect 32309 12251 32367 12257
rect 33502 12248 33508 12300
rect 33560 12288 33566 12300
rect 33560 12260 33605 12288
rect 33560 12248 33566 12260
rect 29380 12192 30604 12220
rect 31754 12180 31760 12232
rect 31812 12220 31818 12232
rect 32125 12223 32183 12229
rect 31812 12192 31857 12220
rect 31812 12180 31818 12192
rect 32125 12189 32137 12223
rect 32171 12220 32183 12223
rect 33042 12220 33048 12232
rect 32171 12192 33048 12220
rect 32171 12189 32183 12192
rect 32125 12183 32183 12189
rect 33042 12180 33048 12192
rect 33100 12180 33106 12232
rect 33137 12223 33195 12229
rect 33137 12189 33149 12223
rect 33183 12198 33195 12223
rect 33183 12189 33272 12198
rect 33137 12183 33272 12189
rect 33152 12170 33272 12183
rect 33318 12180 33324 12232
rect 33376 12220 33382 12232
rect 33376 12192 33421 12220
rect 33376 12180 33382 12192
rect 33778 12180 33784 12232
rect 33836 12220 33842 12232
rect 34057 12223 34115 12229
rect 34057 12220 34069 12223
rect 33836 12192 34069 12220
rect 33836 12180 33842 12192
rect 34057 12189 34069 12192
rect 34103 12189 34115 12223
rect 34057 12183 34115 12189
rect 29794 12155 29852 12161
rect 29794 12152 29806 12155
rect 29288 12124 29806 12152
rect 29794 12121 29806 12124
rect 29840 12121 29852 12155
rect 32858 12152 32864 12164
rect 29794 12115 29852 12121
rect 32140 12124 32864 12152
rect 27304 12056 28212 12084
rect 27304 12044 27310 12056
rect 28902 12044 28908 12096
rect 28960 12084 28966 12096
rect 32140 12084 32168 12124
rect 32858 12112 32864 12124
rect 32916 12112 32922 12164
rect 33244 12152 33272 12170
rect 34256 12152 34284 12328
rect 34793 12325 34805 12359
rect 34839 12356 34851 12359
rect 34839 12328 35204 12356
rect 34839 12325 34851 12328
rect 34793 12319 34851 12325
rect 34330 12248 34336 12300
rect 34388 12288 34394 12300
rect 35176 12288 35204 12328
rect 35250 12316 35256 12368
rect 35308 12356 35314 12368
rect 36357 12359 36415 12365
rect 36357 12356 36369 12359
rect 35308 12328 36369 12356
rect 35308 12316 35314 12328
rect 36357 12325 36369 12328
rect 36403 12325 36415 12359
rect 36357 12319 36415 12325
rect 36538 12316 36544 12368
rect 36596 12356 36602 12368
rect 38010 12356 38016 12368
rect 36596 12328 38016 12356
rect 36596 12316 36602 12328
rect 38010 12316 38016 12328
rect 38068 12316 38074 12368
rect 39316 12356 39344 12396
rect 39390 12384 39396 12436
rect 39448 12424 39454 12436
rect 39448 12396 39493 12424
rect 40972 12396 42196 12424
rect 39448 12384 39454 12396
rect 40972 12356 41000 12396
rect 39316 12328 41000 12356
rect 42168 12356 42196 12396
rect 42242 12384 42248 12436
rect 42300 12424 42306 12436
rect 42337 12427 42395 12433
rect 42337 12424 42349 12427
rect 42300 12396 42349 12424
rect 42300 12384 42306 12396
rect 42337 12393 42349 12396
rect 42383 12393 42395 12427
rect 42337 12387 42395 12393
rect 43901 12427 43959 12433
rect 43901 12393 43913 12427
rect 43947 12424 43959 12427
rect 44082 12424 44088 12436
rect 43947 12396 44088 12424
rect 43947 12393 43959 12396
rect 43901 12387 43959 12393
rect 44082 12384 44088 12396
rect 44140 12384 44146 12436
rect 44174 12384 44180 12436
rect 44232 12424 44238 12436
rect 45738 12424 45744 12436
rect 44232 12396 45744 12424
rect 44232 12384 44238 12396
rect 45738 12384 45744 12396
rect 45796 12424 45802 12436
rect 45796 12396 46704 12424
rect 45796 12384 45802 12396
rect 45373 12359 45431 12365
rect 42168 12328 44128 12356
rect 35526 12288 35532 12300
rect 34388 12260 35112 12288
rect 35176 12260 35532 12288
rect 34388 12248 34394 12260
rect 34606 12180 34612 12232
rect 34664 12220 34670 12232
rect 34977 12223 35035 12229
rect 34977 12220 34989 12223
rect 34664 12192 34989 12220
rect 34664 12180 34670 12192
rect 34977 12189 34989 12192
rect 35023 12189 35035 12223
rect 35084 12220 35112 12260
rect 35526 12248 35532 12260
rect 35584 12248 35590 12300
rect 35618 12248 35624 12300
rect 35676 12288 35682 12300
rect 35676 12260 35848 12288
rect 35676 12248 35682 12260
rect 35820 12229 35848 12260
rect 36078 12248 36084 12300
rect 36136 12288 36142 12300
rect 37461 12291 37519 12297
rect 36136 12260 36860 12288
rect 36136 12248 36142 12260
rect 36832 12232 36860 12260
rect 37461 12257 37473 12291
rect 37507 12288 37519 12291
rect 37550 12288 37556 12300
rect 37507 12260 37556 12288
rect 37507 12257 37519 12260
rect 37461 12251 37519 12257
rect 37550 12248 37556 12260
rect 37608 12248 37614 12300
rect 40954 12288 40960 12300
rect 39859 12260 40356 12288
rect 40915 12260 40960 12288
rect 35713 12223 35771 12229
rect 35713 12220 35725 12223
rect 35084 12192 35725 12220
rect 34977 12183 35035 12189
rect 35713 12189 35725 12192
rect 35759 12189 35771 12223
rect 35713 12183 35771 12189
rect 35805 12223 35863 12229
rect 35805 12189 35817 12223
rect 35851 12189 35863 12223
rect 36538 12220 36544 12232
rect 36499 12192 36544 12220
rect 35805 12183 35863 12189
rect 35250 12152 35256 12164
rect 33244 12124 33609 12152
rect 34256 12124 35256 12152
rect 28960 12056 32168 12084
rect 28960 12044 28966 12056
rect 32214 12044 32220 12096
rect 32272 12084 32278 12096
rect 32950 12084 32956 12096
rect 32272 12056 32956 12084
rect 32272 12044 32278 12056
rect 32950 12044 32956 12056
rect 33008 12044 33014 12096
rect 33581 12084 33609 12124
rect 35250 12112 35256 12124
rect 35308 12112 35314 12164
rect 35728 12152 35756 12183
rect 36538 12180 36544 12192
rect 36596 12180 36602 12232
rect 36722 12220 36728 12232
rect 36683 12192 36728 12220
rect 36722 12180 36728 12192
rect 36780 12180 36786 12232
rect 36814 12180 36820 12232
rect 36872 12220 36878 12232
rect 36872 12192 36917 12220
rect 36872 12180 36878 12192
rect 37090 12180 37096 12232
rect 37148 12220 37154 12232
rect 37185 12223 37243 12229
rect 37185 12220 37197 12223
rect 37148 12192 37197 12220
rect 37148 12180 37154 12192
rect 37185 12189 37197 12192
rect 37231 12189 37243 12223
rect 38010 12220 38016 12232
rect 37971 12192 38016 12220
rect 37185 12183 37243 12189
rect 38010 12180 38016 12192
rect 38068 12180 38074 12232
rect 38102 12180 38108 12232
rect 38160 12220 38166 12232
rect 38269 12223 38327 12229
rect 38269 12220 38281 12223
rect 38160 12192 38281 12220
rect 38160 12180 38166 12192
rect 38269 12189 38281 12192
rect 38315 12189 38327 12223
rect 38269 12183 38327 12189
rect 38562 12180 38568 12232
rect 38620 12220 38626 12232
rect 39859 12220 39887 12260
rect 40034 12220 40040 12232
rect 38620 12192 39887 12220
rect 39995 12192 40040 12220
rect 38620 12180 38626 12192
rect 40034 12180 40040 12192
rect 40092 12180 40098 12232
rect 40218 12220 40224 12232
rect 40179 12192 40224 12220
rect 40218 12180 40224 12192
rect 40276 12180 40282 12232
rect 40328 12220 40356 12260
rect 40954 12248 40960 12260
rect 41012 12248 41018 12300
rect 42705 12291 42763 12297
rect 42705 12257 42717 12291
rect 42751 12288 42763 12291
rect 43346 12288 43352 12300
rect 42751 12260 43352 12288
rect 42751 12257 42763 12260
rect 42705 12251 42763 12257
rect 43346 12248 43352 12260
rect 43404 12248 43410 12300
rect 44100 12288 44128 12328
rect 45373 12325 45385 12359
rect 45419 12356 45431 12359
rect 46014 12356 46020 12368
rect 45419 12328 46020 12356
rect 45419 12325 45431 12328
rect 45373 12319 45431 12325
rect 46014 12316 46020 12328
rect 46072 12316 46078 12368
rect 46290 12356 46296 12368
rect 46251 12328 46296 12356
rect 46290 12316 46296 12328
rect 46348 12316 46354 12368
rect 44100 12260 44496 12288
rect 40405 12223 40463 12229
rect 40405 12220 40417 12223
rect 40328 12192 40417 12220
rect 40405 12189 40417 12192
rect 40451 12216 40463 12223
rect 40494 12216 40500 12232
rect 40451 12189 40500 12216
rect 40405 12188 40500 12189
rect 40405 12183 40463 12188
rect 40494 12180 40500 12188
rect 40552 12180 40558 12232
rect 42978 12220 42984 12232
rect 42939 12192 42984 12220
rect 42978 12180 42984 12192
rect 43036 12180 43042 12232
rect 44100 12229 44128 12260
rect 44085 12223 44143 12229
rect 44085 12189 44097 12223
rect 44131 12189 44143 12223
rect 44358 12220 44364 12232
rect 44319 12192 44364 12220
rect 44085 12183 44143 12189
rect 44358 12180 44364 12192
rect 44416 12180 44422 12232
rect 44468 12220 44496 12260
rect 45462 12248 45468 12300
rect 45520 12288 45526 12300
rect 46198 12288 46204 12300
rect 45520 12260 46204 12288
rect 45520 12248 45526 12260
rect 46198 12248 46204 12260
rect 46256 12288 46262 12300
rect 46676 12297 46704 12396
rect 48222 12384 48228 12436
rect 48280 12424 48286 12436
rect 49421 12427 49479 12433
rect 48280 12396 48544 12424
rect 48280 12384 48286 12396
rect 48038 12316 48044 12368
rect 48096 12356 48102 12368
rect 48516 12356 48544 12396
rect 49421 12393 49433 12427
rect 49467 12424 49479 12427
rect 50982 12424 50988 12436
rect 49467 12396 50988 12424
rect 49467 12393 49479 12396
rect 49421 12387 49479 12393
rect 50982 12384 50988 12396
rect 51040 12384 51046 12436
rect 53009 12427 53067 12433
rect 51092 12396 52592 12424
rect 51092 12356 51120 12396
rect 48096 12328 48452 12356
rect 48516 12328 51120 12356
rect 52564 12356 52592 12396
rect 53009 12393 53021 12427
rect 53055 12424 53067 12427
rect 53098 12424 53104 12436
rect 53055 12396 53104 12424
rect 53055 12393 53067 12396
rect 53009 12387 53067 12393
rect 53098 12384 53104 12396
rect 53156 12384 53162 12436
rect 53282 12384 53288 12436
rect 53340 12424 53346 12436
rect 53926 12424 53932 12436
rect 53340 12396 53932 12424
rect 53340 12384 53346 12396
rect 53926 12384 53932 12396
rect 53984 12384 53990 12436
rect 54021 12427 54079 12433
rect 54021 12393 54033 12427
rect 54067 12424 54079 12427
rect 55398 12424 55404 12436
rect 54067 12396 55404 12424
rect 54067 12393 54079 12396
rect 54021 12387 54079 12393
rect 55398 12384 55404 12396
rect 55456 12384 55462 12436
rect 57054 12424 57060 12436
rect 55508 12396 57060 12424
rect 53374 12356 53380 12368
rect 52564 12328 53380 12356
rect 48096 12316 48102 12328
rect 46477 12291 46535 12297
rect 46477 12288 46489 12291
rect 46256 12260 46489 12288
rect 46256 12248 46262 12260
rect 46477 12257 46489 12260
rect 46523 12257 46535 12291
rect 46477 12251 46535 12257
rect 46661 12291 46719 12297
rect 46661 12257 46673 12291
rect 46707 12257 46719 12291
rect 46661 12251 46719 12257
rect 46842 12248 46848 12300
rect 46900 12288 46906 12300
rect 47302 12288 47308 12300
rect 46900 12260 47308 12288
rect 46900 12248 46906 12260
rect 47302 12248 47308 12260
rect 47360 12248 47366 12300
rect 45554 12220 45560 12232
rect 44468 12192 45560 12220
rect 45554 12180 45560 12192
rect 45612 12180 45618 12232
rect 45833 12223 45891 12229
rect 45833 12214 45845 12223
rect 45756 12189 45845 12214
rect 45879 12189 45891 12223
rect 46566 12220 46572 12232
rect 46527 12192 46572 12220
rect 45756 12186 45891 12189
rect 39666 12152 39672 12164
rect 35728 12124 39672 12152
rect 39666 12112 39672 12124
rect 39724 12112 39730 12164
rect 40126 12112 40132 12164
rect 40184 12152 40190 12164
rect 41230 12161 41236 12164
rect 40313 12155 40371 12161
rect 40313 12152 40325 12155
rect 40184 12124 40325 12152
rect 40184 12112 40190 12124
rect 40313 12121 40325 12124
rect 40359 12121 40371 12155
rect 40313 12115 40371 12121
rect 40420 12124 40724 12152
rect 34974 12084 34980 12096
rect 33581 12056 34980 12084
rect 34974 12044 34980 12056
rect 35032 12044 35038 12096
rect 35158 12084 35164 12096
rect 35119 12056 35164 12084
rect 35158 12044 35164 12056
rect 35216 12044 35222 12096
rect 35894 12044 35900 12096
rect 35952 12084 35958 12096
rect 36170 12084 36176 12096
rect 35952 12056 36176 12084
rect 35952 12044 35958 12056
rect 36170 12044 36176 12056
rect 36228 12044 36234 12096
rect 36262 12044 36268 12096
rect 36320 12084 36326 12096
rect 40420 12084 40448 12124
rect 40586 12084 40592 12096
rect 36320 12056 40448 12084
rect 40547 12056 40592 12084
rect 36320 12044 36326 12056
rect 40586 12044 40592 12056
rect 40644 12044 40650 12096
rect 40696 12084 40724 12124
rect 41224 12115 41236 12161
rect 41288 12152 41294 12164
rect 41288 12124 41324 12152
rect 41230 12112 41236 12115
rect 41288 12112 41294 12124
rect 43162 12112 43168 12164
rect 43220 12152 43226 12164
rect 45756 12152 45784 12186
rect 45833 12183 45891 12186
rect 46566 12180 46572 12192
rect 46624 12180 46630 12232
rect 46753 12223 46811 12229
rect 46753 12189 46765 12223
rect 46799 12220 46811 12223
rect 47578 12220 47584 12232
rect 46799 12192 47584 12220
rect 46799 12189 46811 12192
rect 46753 12183 46811 12189
rect 47578 12180 47584 12192
rect 47636 12180 47642 12232
rect 48041 12223 48099 12229
rect 48041 12189 48053 12223
rect 48087 12220 48099 12223
rect 48314 12220 48320 12232
rect 48087 12192 48320 12220
rect 48087 12189 48099 12192
rect 48041 12183 48099 12189
rect 48314 12180 48320 12192
rect 48372 12180 48378 12232
rect 48424 12229 48452 12328
rect 53374 12316 53380 12328
rect 53432 12316 53438 12368
rect 53834 12316 53840 12368
rect 53892 12356 53898 12368
rect 54757 12359 54815 12365
rect 54757 12356 54769 12359
rect 53892 12328 54769 12356
rect 53892 12316 53898 12328
rect 54757 12325 54769 12328
rect 54803 12325 54815 12359
rect 55508 12356 55536 12396
rect 57054 12384 57060 12396
rect 57112 12384 57118 12436
rect 57146 12384 57152 12436
rect 57204 12424 57210 12436
rect 57514 12424 57520 12436
rect 57204 12396 57520 12424
rect 57204 12384 57210 12396
rect 57514 12384 57520 12396
rect 57572 12384 57578 12436
rect 58345 12427 58403 12433
rect 58345 12393 58357 12427
rect 58391 12424 58403 12427
rect 59630 12424 59636 12436
rect 58391 12396 59636 12424
rect 58391 12393 58403 12396
rect 58345 12387 58403 12393
rect 59630 12384 59636 12396
rect 59688 12384 59694 12436
rect 59906 12384 59912 12436
rect 59964 12424 59970 12436
rect 61838 12424 61844 12436
rect 59964 12396 61700 12424
rect 61799 12396 61844 12424
rect 59964 12384 59970 12396
rect 54757 12319 54815 12325
rect 55232 12328 55536 12356
rect 55232 12300 55260 12328
rect 56594 12316 56600 12368
rect 56652 12356 56658 12368
rect 57790 12356 57796 12368
rect 56652 12328 57796 12356
rect 56652 12316 56658 12328
rect 57790 12316 57796 12328
rect 57848 12316 57854 12368
rect 57882 12316 57888 12368
rect 57940 12356 57946 12368
rect 61672 12356 61700 12396
rect 61838 12384 61844 12396
rect 61896 12384 61902 12436
rect 61948 12396 63448 12424
rect 61948 12356 61976 12396
rect 63420 12356 63448 12396
rect 63494 12384 63500 12436
rect 63552 12424 63558 12436
rect 64049 12427 64107 12433
rect 64049 12424 64061 12427
rect 63552 12396 64061 12424
rect 63552 12384 63558 12396
rect 64049 12393 64061 12396
rect 64095 12424 64107 12427
rect 64782 12424 64788 12436
rect 64095 12396 64788 12424
rect 64095 12393 64107 12396
rect 64049 12387 64107 12393
rect 64782 12384 64788 12396
rect 64840 12384 64846 12436
rect 64877 12427 64935 12433
rect 64877 12393 64889 12427
rect 64923 12424 64935 12427
rect 65150 12424 65156 12436
rect 64923 12396 65156 12424
rect 64923 12393 64935 12396
rect 64877 12387 64935 12393
rect 65150 12384 65156 12396
rect 65208 12384 65214 12436
rect 65705 12427 65763 12433
rect 65705 12393 65717 12427
rect 65751 12424 65763 12427
rect 65978 12424 65984 12436
rect 65751 12396 65984 12424
rect 65751 12393 65763 12396
rect 65705 12387 65763 12393
rect 65978 12384 65984 12396
rect 66036 12384 66042 12436
rect 67542 12424 67548 12436
rect 66088 12396 67548 12424
rect 66088 12365 66116 12396
rect 67542 12384 67548 12396
rect 67600 12384 67606 12436
rect 67910 12424 67916 12436
rect 67871 12396 67916 12424
rect 67910 12384 67916 12396
rect 67968 12384 67974 12436
rect 68554 12384 68560 12436
rect 68612 12424 68618 12436
rect 69106 12424 69112 12436
rect 68612 12396 69112 12424
rect 68612 12384 68618 12396
rect 69106 12384 69112 12396
rect 69164 12384 69170 12436
rect 69290 12384 69296 12436
rect 69348 12424 69354 12436
rect 69474 12424 69480 12436
rect 69348 12396 69480 12424
rect 69348 12384 69354 12396
rect 69474 12384 69480 12396
rect 69532 12384 69538 12436
rect 70029 12427 70087 12433
rect 70029 12424 70041 12427
rect 69584 12396 70041 12424
rect 66073 12359 66131 12365
rect 57940 12328 59492 12356
rect 61672 12328 61976 12356
rect 62040 12328 62519 12356
rect 63420 12328 65932 12356
rect 57940 12316 57946 12328
rect 48501 12291 48559 12297
rect 48501 12257 48513 12291
rect 48547 12288 48559 12291
rect 48958 12288 48964 12300
rect 48547 12260 48964 12288
rect 48547 12257 48559 12260
rect 48501 12251 48559 12257
rect 48958 12248 48964 12260
rect 49016 12248 49022 12300
rect 50430 12288 50436 12300
rect 49436 12260 50436 12288
rect 48409 12223 48467 12229
rect 48409 12189 48421 12223
rect 48455 12189 48467 12223
rect 48590 12220 48596 12232
rect 48551 12192 48596 12220
rect 48409 12183 48467 12189
rect 48590 12180 48596 12192
rect 48648 12180 48654 12232
rect 49436 12164 49464 12260
rect 50430 12248 50436 12260
rect 50488 12248 50494 12300
rect 55122 12288 55128 12300
rect 53398 12260 55128 12288
rect 49694 12220 49700 12232
rect 49655 12192 49700 12220
rect 49694 12180 49700 12192
rect 49752 12180 49758 12232
rect 49970 12180 49976 12232
rect 50028 12220 50034 12232
rect 50157 12223 50215 12229
rect 50157 12220 50169 12223
rect 50028 12192 50169 12220
rect 50028 12180 50034 12192
rect 50157 12189 50169 12192
rect 50203 12220 50215 12223
rect 50246 12220 50252 12232
rect 50203 12192 50252 12220
rect 50203 12189 50215 12192
rect 50157 12183 50215 12189
rect 50246 12180 50252 12192
rect 50304 12180 50310 12232
rect 50338 12180 50344 12232
rect 50396 12220 50402 12232
rect 51629 12223 51687 12229
rect 51629 12220 51641 12223
rect 50396 12192 51641 12220
rect 50396 12180 50402 12192
rect 51629 12189 51641 12192
rect 51675 12189 51687 12223
rect 53398 12220 53426 12260
rect 55122 12248 55128 12260
rect 55180 12248 55186 12300
rect 55214 12248 55220 12300
rect 55272 12248 55278 12300
rect 55324 12260 55628 12288
rect 51629 12183 51687 12189
rect 51828 12192 53426 12220
rect 53469 12223 53527 12229
rect 43220 12124 45784 12152
rect 43220 12112 43226 12124
rect 46290 12112 46296 12164
rect 46348 12152 46354 12164
rect 47762 12152 47768 12164
rect 46348 12124 47768 12152
rect 46348 12112 46354 12124
rect 47762 12112 47768 12124
rect 47820 12112 47826 12164
rect 48222 12112 48228 12164
rect 48280 12152 48286 12164
rect 49418 12152 49424 12164
rect 48280 12112 48314 12152
rect 49379 12124 49424 12152
rect 49418 12112 49424 12124
rect 49476 12112 49482 12164
rect 49605 12155 49663 12161
rect 49605 12121 49617 12155
rect 49651 12152 49663 12155
rect 51828 12152 51856 12192
rect 53469 12189 53481 12223
rect 53515 12222 53527 12223
rect 53558 12222 53564 12232
rect 53515 12194 53564 12222
rect 53515 12189 53527 12194
rect 53469 12183 53527 12189
rect 53558 12180 53564 12194
rect 53616 12180 53622 12232
rect 54294 12220 54300 12232
rect 53668 12192 54156 12220
rect 54255 12192 54300 12220
rect 49651 12124 51856 12152
rect 51896 12155 51954 12161
rect 49651 12121 49663 12124
rect 49605 12115 49663 12121
rect 51896 12121 51908 12155
rect 51942 12152 51954 12155
rect 52086 12152 52092 12164
rect 51942 12124 52092 12152
rect 51942 12121 51954 12124
rect 51896 12115 51954 12121
rect 52086 12112 52092 12124
rect 52144 12112 52150 12164
rect 53668 12152 53696 12192
rect 52196 12124 53696 12152
rect 41598 12084 41604 12096
rect 40696 12056 41604 12084
rect 41598 12044 41604 12056
rect 41656 12044 41662 12096
rect 43806 12044 43812 12096
rect 43864 12084 43870 12096
rect 44269 12087 44327 12093
rect 44269 12084 44281 12087
rect 43864 12056 44281 12084
rect 43864 12044 43870 12056
rect 44269 12053 44281 12056
rect 44315 12084 44327 12087
rect 45741 12087 45799 12093
rect 45741 12084 45753 12087
rect 44315 12056 45753 12084
rect 44315 12053 44327 12056
rect 44269 12047 44327 12053
rect 45741 12053 45753 12056
rect 45787 12084 45799 12087
rect 47670 12084 47676 12096
rect 45787 12056 47676 12084
rect 45787 12053 45799 12056
rect 45741 12047 45799 12053
rect 47670 12044 47676 12056
rect 47728 12044 47734 12096
rect 47854 12044 47860 12096
rect 47912 12084 47918 12096
rect 48286 12084 48314 12112
rect 52196 12084 52224 12124
rect 53742 12112 53748 12164
rect 53800 12152 53806 12164
rect 54021 12155 54079 12161
rect 54021 12152 54033 12155
rect 53800 12124 54033 12152
rect 53800 12112 53806 12124
rect 54021 12121 54033 12124
rect 54067 12121 54079 12155
rect 54128 12152 54156 12192
rect 54294 12180 54300 12192
rect 54352 12180 54358 12232
rect 54662 12220 54668 12232
rect 54623 12192 54668 12220
rect 54662 12180 54668 12192
rect 54720 12180 54726 12232
rect 55324 12152 55352 12260
rect 55398 12180 55404 12232
rect 55456 12222 55462 12232
rect 55493 12223 55551 12229
rect 55493 12222 55505 12223
rect 55456 12194 55505 12222
rect 55456 12180 55462 12194
rect 55493 12189 55505 12194
rect 55539 12189 55551 12223
rect 55600 12220 55628 12260
rect 56778 12248 56784 12300
rect 56836 12288 56842 12300
rect 57241 12291 57299 12297
rect 57241 12288 57253 12291
rect 56836 12260 57253 12288
rect 56836 12248 56842 12260
rect 57241 12257 57253 12260
rect 57287 12257 57299 12291
rect 57241 12251 57299 12257
rect 57532 12260 58572 12288
rect 55600 12192 55904 12220
rect 55493 12183 55551 12189
rect 54128 12124 55352 12152
rect 54021 12115 54079 12121
rect 55582 12112 55588 12164
rect 55640 12152 55646 12164
rect 55738 12155 55796 12161
rect 55738 12152 55750 12155
rect 55640 12124 55750 12152
rect 55640 12112 55646 12124
rect 55738 12121 55750 12124
rect 55784 12121 55796 12155
rect 55876 12152 55904 12192
rect 57054 12180 57060 12232
rect 57112 12220 57118 12232
rect 57425 12223 57483 12229
rect 57425 12220 57437 12223
rect 57112 12192 57437 12220
rect 57112 12180 57118 12192
rect 57425 12189 57437 12192
rect 57471 12220 57483 12223
rect 57532 12220 57560 12260
rect 57471 12192 57560 12220
rect 57471 12189 57483 12192
rect 57425 12183 57483 12189
rect 57606 12180 57612 12232
rect 57664 12220 57670 12232
rect 57701 12223 57759 12229
rect 57701 12220 57713 12223
rect 57664 12192 57713 12220
rect 57664 12180 57670 12192
rect 57701 12189 57713 12192
rect 57747 12220 57759 12223
rect 57790 12220 57796 12232
rect 57747 12192 57796 12220
rect 57747 12189 57759 12192
rect 57701 12183 57759 12189
rect 57790 12180 57796 12192
rect 57848 12180 57854 12232
rect 57974 12180 57980 12232
rect 58032 12220 58038 12232
rect 58544 12229 58572 12260
rect 59170 12248 59176 12300
rect 59228 12288 59234 12300
rect 59228 12260 59273 12288
rect 59228 12248 59234 12260
rect 59464 12229 59492 12328
rect 60458 12288 60464 12300
rect 60419 12260 60464 12288
rect 60458 12248 60464 12260
rect 60516 12248 60522 12300
rect 58529 12223 58587 12229
rect 58032 12192 58480 12220
rect 58032 12180 58038 12192
rect 58342 12152 58348 12164
rect 55876 12124 58348 12152
rect 55738 12115 55796 12121
rect 58342 12112 58348 12124
rect 58400 12112 58406 12164
rect 58452 12152 58480 12192
rect 58529 12189 58541 12223
rect 58575 12189 58587 12223
rect 58529 12183 58587 12189
rect 58805 12223 58863 12229
rect 58805 12189 58817 12223
rect 58851 12220 58863 12223
rect 59449 12223 59507 12229
rect 58851 12192 59216 12220
rect 58851 12189 58863 12192
rect 58805 12183 58863 12189
rect 58820 12152 58848 12183
rect 59188 12164 59216 12192
rect 59449 12189 59461 12223
rect 59495 12189 59507 12223
rect 59449 12183 59507 12189
rect 58452 12124 58848 12152
rect 59170 12112 59176 12164
rect 59228 12112 59234 12164
rect 59464 12152 59492 12183
rect 59998 12180 60004 12232
rect 60056 12220 60062 12232
rect 62040 12220 62068 12328
rect 62491 12288 62519 12328
rect 65904 12297 65932 12328
rect 66073 12325 66085 12359
rect 66119 12325 66131 12359
rect 66073 12319 66131 12325
rect 68646 12316 68652 12368
rect 68704 12356 68710 12368
rect 69382 12356 69388 12368
rect 68704 12328 69388 12356
rect 68704 12316 68710 12328
rect 69382 12316 69388 12328
rect 69440 12316 69446 12368
rect 64233 12291 64291 12297
rect 64233 12288 64245 12291
rect 62491 12260 64245 12288
rect 64233 12257 64245 12260
rect 64279 12257 64291 12291
rect 64233 12251 64291 12257
rect 64417 12291 64475 12297
rect 64417 12257 64429 12291
rect 64463 12288 64475 12291
rect 65889 12291 65947 12297
rect 64463 12260 65288 12288
rect 64463 12257 64475 12260
rect 64417 12251 64475 12257
rect 62396 12233 62454 12239
rect 62298 12220 62304 12232
rect 60056 12192 62068 12220
rect 62259 12192 62304 12220
rect 60056 12180 60062 12192
rect 62298 12180 62304 12192
rect 62356 12180 62362 12232
rect 62396 12199 62408 12233
rect 62442 12220 62454 12233
rect 62442 12199 62519 12220
rect 62396 12193 62519 12199
rect 62411 12192 62519 12193
rect 60734 12161 60740 12164
rect 59464 12124 60688 12152
rect 60660 12096 60688 12124
rect 60728 12115 60740 12161
rect 60792 12152 60798 12164
rect 60792 12124 60828 12152
rect 60734 12112 60740 12115
rect 60792 12112 60798 12124
rect 62390 12112 62396 12164
rect 62448 12152 62454 12164
rect 62491 12152 62519 12192
rect 62666 12180 62672 12232
rect 62724 12220 62730 12232
rect 63037 12223 63095 12229
rect 63037 12220 63049 12223
rect 62724 12192 63049 12220
rect 62724 12180 62730 12192
rect 63037 12189 63049 12192
rect 63083 12189 63095 12223
rect 63218 12220 63224 12232
rect 63179 12192 63224 12220
rect 63037 12183 63095 12189
rect 63218 12180 63224 12192
rect 63276 12180 63282 12232
rect 64046 12180 64052 12232
rect 64104 12220 64110 12232
rect 64506 12220 64512 12232
rect 64104 12192 64512 12220
rect 64104 12180 64110 12192
rect 64506 12180 64512 12192
rect 64564 12180 64570 12232
rect 64690 12180 64696 12232
rect 64748 12220 64754 12232
rect 65153 12223 65211 12229
rect 65153 12220 65165 12223
rect 64748 12192 65165 12220
rect 64748 12180 64754 12192
rect 65153 12189 65165 12192
rect 65199 12189 65211 12223
rect 65153 12183 65211 12189
rect 62448 12124 62519 12152
rect 62577 12155 62635 12161
rect 62448 12112 62454 12124
rect 62577 12121 62589 12155
rect 62623 12152 62635 12155
rect 64414 12152 64420 12164
rect 62623 12124 64420 12152
rect 62623 12121 62635 12124
rect 62577 12115 62635 12121
rect 64414 12112 64420 12124
rect 64472 12112 64478 12164
rect 64874 12152 64880 12164
rect 64835 12124 64880 12152
rect 64874 12112 64880 12124
rect 64932 12112 64938 12164
rect 65260 12152 65288 12260
rect 65889 12257 65901 12291
rect 65935 12257 65947 12291
rect 69584 12288 69612 12396
rect 70029 12393 70041 12396
rect 70075 12393 70087 12427
rect 70029 12387 70087 12393
rect 70210 12384 70216 12436
rect 70268 12424 70274 12436
rect 82170 12424 82176 12436
rect 70268 12396 82176 12424
rect 70268 12384 70274 12396
rect 82170 12384 82176 12396
rect 82228 12384 82234 12436
rect 72145 12359 72203 12365
rect 72145 12325 72157 12359
rect 72191 12356 72203 12359
rect 72326 12356 72332 12368
rect 72191 12328 72332 12356
rect 72191 12325 72203 12328
rect 72145 12319 72203 12325
rect 72326 12316 72332 12328
rect 72384 12316 72390 12368
rect 72513 12359 72571 12365
rect 72513 12325 72525 12359
rect 72559 12356 72571 12359
rect 87138 12356 87144 12368
rect 72559 12328 72832 12356
rect 72559 12325 72571 12328
rect 72513 12319 72571 12325
rect 70762 12288 70768 12300
rect 65889 12251 65947 12257
rect 67560 12260 68692 12288
rect 65334 12180 65340 12232
rect 65392 12220 65398 12232
rect 66165 12223 66223 12229
rect 66165 12220 66177 12223
rect 65392 12192 66177 12220
rect 65392 12180 65398 12192
rect 66165 12189 66177 12192
rect 66211 12189 66223 12223
rect 66530 12220 66536 12232
rect 66491 12192 66536 12220
rect 66165 12183 66223 12189
rect 66530 12180 66536 12192
rect 66588 12180 66594 12232
rect 67560 12220 67588 12260
rect 66732 12192 67588 12220
rect 66732 12152 66760 12192
rect 65260 12124 66760 12152
rect 66800 12155 66858 12161
rect 66800 12121 66812 12155
rect 66846 12152 66858 12155
rect 67174 12152 67180 12164
rect 66846 12124 67180 12152
rect 66846 12121 66858 12124
rect 66800 12115 66858 12121
rect 67174 12112 67180 12124
rect 67232 12112 67238 12164
rect 67266 12112 67272 12164
rect 67324 12152 67330 12164
rect 68554 12152 68560 12164
rect 67324 12124 68560 12152
rect 67324 12112 67330 12124
rect 68554 12112 68560 12124
rect 68612 12112 68618 12164
rect 68664 12152 68692 12260
rect 68756 12260 69612 12288
rect 70723 12260 70768 12288
rect 68756 12229 68784 12260
rect 70762 12248 70768 12260
rect 70820 12248 70826 12300
rect 68741 12223 68799 12229
rect 68741 12189 68753 12223
rect 68787 12189 68799 12223
rect 68922 12220 68928 12232
rect 68883 12192 68928 12220
rect 68741 12183 68799 12189
rect 68922 12180 68928 12192
rect 68980 12180 68986 12232
rect 69308 12192 69612 12220
rect 69308 12161 69336 12192
rect 69293 12155 69351 12161
rect 69293 12152 69305 12155
rect 68664 12124 69305 12152
rect 69293 12121 69305 12124
rect 69339 12121 69351 12155
rect 69293 12115 69351 12121
rect 69382 12112 69388 12164
rect 69440 12152 69446 12164
rect 69493 12155 69551 12161
rect 69493 12152 69505 12155
rect 69440 12124 69505 12152
rect 69440 12112 69446 12124
rect 69493 12121 69505 12124
rect 69539 12121 69551 12155
rect 69584 12152 69612 12192
rect 69658 12180 69664 12232
rect 69716 12220 69722 12232
rect 70302 12220 70308 12232
rect 69716 12192 70164 12220
rect 70263 12192 70308 12220
rect 69716 12180 69722 12192
rect 70136 12164 70164 12192
rect 70302 12180 70308 12192
rect 70360 12180 70366 12232
rect 71314 12180 71320 12232
rect 71372 12220 71378 12232
rect 72697 12223 72755 12229
rect 72697 12220 72709 12223
rect 71372 12192 72709 12220
rect 71372 12180 71378 12192
rect 72697 12189 72709 12192
rect 72743 12189 72755 12223
rect 72697 12183 72755 12189
rect 70026 12152 70032 12164
rect 69584 12124 70032 12152
rect 69493 12115 69551 12121
rect 70026 12112 70032 12124
rect 70084 12112 70090 12164
rect 70118 12112 70124 12164
rect 70176 12152 70182 12164
rect 70213 12155 70271 12161
rect 70213 12152 70225 12155
rect 70176 12124 70225 12152
rect 70176 12112 70182 12124
rect 70213 12121 70225 12124
rect 70259 12121 70271 12155
rect 70213 12115 70271 12121
rect 71032 12155 71090 12161
rect 71032 12121 71044 12155
rect 71078 12152 71090 12155
rect 72804 12152 72832 12328
rect 71078 12124 72832 12152
rect 80026 12328 87144 12356
rect 71078 12121 71090 12124
rect 71032 12115 71090 12121
rect 47912 12056 47957 12084
rect 48286 12056 52224 12084
rect 47912 12044 47918 12056
rect 52822 12044 52828 12096
rect 52880 12084 52886 12096
rect 53561 12087 53619 12093
rect 53561 12084 53573 12087
rect 52880 12056 53573 12084
rect 52880 12044 52886 12056
rect 53561 12053 53573 12056
rect 53607 12084 53619 12087
rect 53650 12084 53656 12096
rect 53607 12056 53656 12084
rect 53607 12053 53619 12056
rect 53561 12047 53619 12053
rect 53650 12044 53656 12056
rect 53708 12044 53714 12096
rect 53926 12044 53932 12096
rect 53984 12084 53990 12096
rect 54205 12087 54263 12093
rect 54205 12084 54217 12087
rect 53984 12056 54217 12084
rect 53984 12044 53990 12056
rect 54205 12053 54217 12056
rect 54251 12084 54263 12087
rect 54754 12084 54760 12096
rect 54251 12056 54760 12084
rect 54251 12053 54263 12056
rect 54205 12047 54263 12053
rect 54754 12044 54760 12056
rect 54812 12044 54818 12096
rect 54846 12044 54852 12096
rect 54904 12084 54910 12096
rect 56594 12084 56600 12096
rect 54904 12056 56600 12084
rect 54904 12044 54910 12056
rect 56594 12044 56600 12056
rect 56652 12044 56658 12096
rect 56873 12087 56931 12093
rect 56873 12053 56885 12087
rect 56919 12084 56931 12087
rect 57609 12087 57667 12093
rect 57609 12084 57621 12087
rect 56919 12056 57621 12084
rect 56919 12053 56931 12056
rect 56873 12047 56931 12053
rect 57609 12053 57621 12056
rect 57655 12053 57667 12087
rect 57609 12047 57667 12053
rect 57790 12044 57796 12096
rect 57848 12084 57854 12096
rect 58618 12084 58624 12096
rect 57848 12056 58624 12084
rect 57848 12044 57854 12056
rect 58618 12044 58624 12056
rect 58676 12044 58682 12096
rect 58713 12087 58771 12093
rect 58713 12053 58725 12087
rect 58759 12084 58771 12087
rect 60366 12084 60372 12096
rect 58759 12056 60372 12084
rect 58759 12053 58771 12056
rect 58713 12047 58771 12053
rect 60366 12044 60372 12056
rect 60424 12044 60430 12096
rect 60642 12044 60648 12096
rect 60700 12044 60706 12096
rect 62758 12044 62764 12096
rect 62816 12084 62822 12096
rect 65061 12087 65119 12093
rect 65061 12084 65073 12087
rect 62816 12056 65073 12084
rect 62816 12044 62822 12056
rect 65061 12053 65073 12056
rect 65107 12084 65119 12087
rect 68094 12084 68100 12096
rect 65107 12056 68100 12084
rect 65107 12053 65119 12056
rect 65061 12047 65119 12053
rect 68094 12044 68100 12056
rect 68152 12044 68158 12096
rect 68830 12084 68836 12096
rect 68791 12056 68836 12084
rect 68830 12044 68836 12056
rect 68888 12044 68894 12096
rect 68922 12044 68928 12096
rect 68980 12084 68986 12096
rect 69661 12087 69719 12093
rect 69661 12084 69673 12087
rect 68980 12056 69673 12084
rect 68980 12044 68986 12056
rect 69661 12053 69673 12056
rect 69707 12053 69719 12087
rect 69661 12047 69719 12053
rect 69750 12044 69756 12096
rect 69808 12084 69814 12096
rect 80026 12084 80054 12328
rect 87138 12316 87144 12328
rect 87196 12316 87202 12368
rect 69808 12056 80054 12084
rect 69808 12044 69814 12056
rect 1104 11994 88872 12016
rect 1104 11942 22898 11994
rect 22950 11942 22962 11994
rect 23014 11942 23026 11994
rect 23078 11942 23090 11994
rect 23142 11942 23154 11994
rect 23206 11942 44846 11994
rect 44898 11942 44910 11994
rect 44962 11942 44974 11994
rect 45026 11942 45038 11994
rect 45090 11942 45102 11994
rect 45154 11942 66794 11994
rect 66846 11942 66858 11994
rect 66910 11942 66922 11994
rect 66974 11942 66986 11994
rect 67038 11942 67050 11994
rect 67102 11942 88872 11994
rect 1104 11920 88872 11942
rect 23566 11880 23572 11892
rect 6886 11852 23572 11880
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 6886 11744 6914 11852
rect 23566 11840 23572 11852
rect 23624 11840 23630 11892
rect 23750 11840 23756 11892
rect 23808 11880 23814 11892
rect 24581 11883 24639 11889
rect 24581 11880 24593 11883
rect 23808 11852 24593 11880
rect 23808 11840 23814 11852
rect 24581 11849 24593 11852
rect 24627 11849 24639 11883
rect 24581 11843 24639 11849
rect 25409 11883 25467 11889
rect 25409 11849 25421 11883
rect 25455 11880 25467 11883
rect 26050 11880 26056 11892
rect 25455 11852 26056 11880
rect 25455 11849 25467 11852
rect 25409 11843 25467 11849
rect 26050 11840 26056 11852
rect 26108 11840 26114 11892
rect 26418 11880 26424 11892
rect 26379 11852 26424 11880
rect 26418 11840 26424 11852
rect 26476 11840 26482 11892
rect 26786 11840 26792 11892
rect 26844 11880 26850 11892
rect 28442 11880 28448 11892
rect 26844 11852 28448 11880
rect 26844 11840 26850 11852
rect 28442 11840 28448 11852
rect 28500 11840 28506 11892
rect 29641 11883 29699 11889
rect 29641 11849 29653 11883
rect 29687 11880 29699 11883
rect 30006 11880 30012 11892
rect 29687 11852 30012 11880
rect 29687 11849 29699 11852
rect 29641 11843 29699 11849
rect 30006 11840 30012 11852
rect 30064 11840 30070 11892
rect 30098 11840 30104 11892
rect 30156 11880 30162 11892
rect 30837 11883 30895 11889
rect 30837 11880 30849 11883
rect 30156 11852 30849 11880
rect 30156 11840 30162 11852
rect 30837 11849 30849 11852
rect 30883 11849 30895 11883
rect 35805 11883 35863 11889
rect 35805 11880 35817 11883
rect 30837 11843 30895 11849
rect 31036 11852 35817 11880
rect 16574 11772 16580 11824
rect 16632 11812 16638 11824
rect 20073 11815 20131 11821
rect 20073 11812 20085 11815
rect 16632 11784 20085 11812
rect 16632 11772 16638 11784
rect 20073 11781 20085 11784
rect 20119 11781 20131 11815
rect 20073 11775 20131 11781
rect 20162 11772 20168 11824
rect 20220 11812 20226 11824
rect 21358 11812 21364 11824
rect 20220 11784 21364 11812
rect 20220 11772 20226 11784
rect 21358 11772 21364 11784
rect 21416 11772 21422 11824
rect 25314 11772 25320 11824
rect 25372 11812 25378 11824
rect 26145 11815 26203 11821
rect 26145 11812 26157 11815
rect 25372 11784 26157 11812
rect 25372 11772 25378 11784
rect 26145 11781 26157 11784
rect 26191 11781 26203 11815
rect 26145 11775 26203 11781
rect 27982 11772 27988 11824
rect 28040 11812 28046 11824
rect 29733 11815 29791 11821
rect 29733 11812 29745 11815
rect 28040 11784 29745 11812
rect 28040 11772 28046 11784
rect 29733 11781 29745 11784
rect 29779 11812 29791 11815
rect 29822 11812 29828 11824
rect 29779 11784 29828 11812
rect 29779 11781 29791 11784
rect 29733 11775 29791 11781
rect 29822 11772 29828 11784
rect 29880 11772 29886 11824
rect 18782 11744 18788 11756
rect 1627 11716 6914 11744
rect 18743 11716 18788 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 18966 11744 18972 11756
rect 18927 11716 18972 11744
rect 18966 11704 18972 11716
rect 19024 11704 19030 11756
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11744 19119 11747
rect 19702 11744 19708 11756
rect 19107 11716 19708 11744
rect 19107 11713 19119 11716
rect 19061 11707 19119 11713
rect 19702 11704 19708 11716
rect 19760 11704 19766 11756
rect 19797 11747 19855 11753
rect 19797 11713 19809 11747
rect 19843 11713 19855 11747
rect 19797 11707 19855 11713
rect 19889 11747 19947 11753
rect 19889 11713 19901 11747
rect 19935 11744 19947 11747
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 19935 11716 20729 11744
rect 19935 11713 19947 11716
rect 19889 11707 19947 11713
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 2648 11648 18828 11676
rect 2648 11636 2654 11648
rect 1394 11608 1400 11620
rect 1355 11580 1400 11608
rect 1394 11568 1400 11580
rect 1452 11568 1458 11620
rect 18598 11540 18604 11552
rect 18559 11512 18604 11540
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 18800 11540 18828 11648
rect 18874 11568 18880 11620
rect 18932 11608 18938 11620
rect 19337 11611 19395 11617
rect 19337 11608 19349 11611
rect 18932 11580 19349 11608
rect 18932 11568 18938 11580
rect 19337 11577 19349 11580
rect 19383 11608 19395 11611
rect 19812 11608 19840 11707
rect 20088 11688 20116 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11744 24179 11747
rect 24302 11744 24308 11756
rect 24167 11716 24308 11744
rect 24167 11713 24179 11716
rect 24121 11707 24179 11713
rect 24302 11704 24308 11716
rect 24360 11744 24366 11756
rect 24578 11744 24584 11756
rect 24360 11716 24584 11744
rect 24360 11704 24366 11716
rect 24578 11704 24584 11716
rect 24636 11704 24642 11756
rect 25774 11744 25780 11756
rect 25735 11716 25780 11744
rect 25774 11704 25780 11716
rect 25832 11704 25838 11756
rect 25866 11704 25872 11756
rect 25924 11744 25930 11756
rect 25924 11716 25969 11744
rect 25924 11704 25930 11716
rect 26050 11704 26056 11756
rect 26108 11744 26114 11756
rect 26326 11753 26332 11756
rect 26283 11747 26332 11753
rect 26108 11716 26153 11744
rect 26108 11704 26114 11716
rect 26283 11713 26295 11747
rect 26329 11713 26332 11747
rect 26283 11707 26332 11713
rect 26326 11704 26332 11707
rect 26384 11704 26390 11756
rect 26510 11704 26516 11756
rect 26568 11744 26574 11756
rect 28994 11744 29000 11756
rect 26568 11716 29000 11744
rect 26568 11704 26574 11716
rect 28994 11704 29000 11716
rect 29052 11704 29058 11756
rect 30834 11744 30840 11756
rect 29748 11716 30840 11744
rect 20070 11636 20076 11688
rect 20128 11636 20134 11688
rect 20990 11636 20996 11688
rect 21048 11676 21054 11688
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 21048 11648 21189 11676
rect 21048 11636 21054 11648
rect 21177 11645 21189 11648
rect 21223 11645 21235 11679
rect 21177 11639 21235 11645
rect 24210 11636 24216 11688
rect 24268 11676 24274 11688
rect 24949 11679 25007 11685
rect 24949 11676 24961 11679
rect 24268 11648 24961 11676
rect 24268 11636 24274 11648
rect 24949 11645 24961 11648
rect 24995 11676 25007 11679
rect 25682 11676 25688 11688
rect 24995 11648 25688 11676
rect 24995 11645 25007 11648
rect 24949 11639 25007 11645
rect 25682 11636 25688 11648
rect 25740 11636 25746 11688
rect 25958 11636 25964 11688
rect 26016 11676 26022 11688
rect 26973 11679 27031 11685
rect 26973 11676 26985 11679
rect 26016 11648 26985 11676
rect 26016 11636 26022 11648
rect 26973 11645 26985 11648
rect 27019 11645 27031 11679
rect 26973 11639 27031 11645
rect 27249 11679 27307 11685
rect 27249 11645 27261 11679
rect 27295 11676 27307 11679
rect 27614 11676 27620 11688
rect 27295 11648 27620 11676
rect 27295 11645 27307 11648
rect 27249 11639 27307 11645
rect 27614 11636 27620 11648
rect 27672 11636 27678 11688
rect 28166 11636 28172 11688
rect 28224 11676 28230 11688
rect 28353 11679 28411 11685
rect 28353 11676 28365 11679
rect 28224 11648 28365 11676
rect 28224 11636 28230 11648
rect 28353 11645 28365 11648
rect 28399 11676 28411 11679
rect 29748 11676 29776 11716
rect 30834 11704 30840 11716
rect 30892 11704 30898 11756
rect 31036 11753 31064 11852
rect 35805 11849 35817 11852
rect 35851 11880 35863 11883
rect 35851 11852 37136 11880
rect 35851 11849 35863 11852
rect 35805 11843 35863 11849
rect 31110 11772 31116 11824
rect 31168 11812 31174 11824
rect 32493 11815 32551 11821
rect 31168 11784 32444 11812
rect 31168 11772 31174 11784
rect 31021 11747 31079 11753
rect 31021 11713 31033 11747
rect 31067 11713 31079 11747
rect 31478 11744 31484 11756
rect 31439 11716 31484 11744
rect 31021 11707 31079 11713
rect 31478 11704 31484 11716
rect 31536 11704 31542 11756
rect 32416 11744 32444 11784
rect 32493 11781 32505 11815
rect 32539 11812 32551 11815
rect 33042 11812 33048 11824
rect 32539 11784 33048 11812
rect 32539 11781 32551 11784
rect 32493 11775 32551 11781
rect 33042 11772 33048 11784
rect 33100 11772 33106 11824
rect 33152 11784 33824 11812
rect 32858 11744 32864 11756
rect 32416 11716 32864 11744
rect 32858 11704 32864 11716
rect 32916 11704 32922 11756
rect 28399 11648 29776 11676
rect 28399 11645 28411 11648
rect 28353 11639 28411 11645
rect 29822 11636 29828 11688
rect 29880 11676 29886 11688
rect 29880 11648 29925 11676
rect 29880 11636 29886 11648
rect 25317 11611 25375 11617
rect 19383 11580 22094 11608
rect 19383 11577 19395 11580
rect 19337 11571 19395 11577
rect 20162 11540 20168 11552
rect 18800 11512 20168 11540
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 20714 11500 20720 11552
rect 20772 11540 20778 11552
rect 20990 11540 20996 11552
rect 20772 11512 20996 11540
rect 20772 11500 20778 11512
rect 20990 11500 20996 11512
rect 21048 11500 21054 11552
rect 22066 11540 22094 11580
rect 25317 11577 25329 11611
rect 25363 11608 25375 11611
rect 26786 11608 26792 11620
rect 25363 11580 26792 11608
rect 25363 11577 25375 11580
rect 25317 11571 25375 11577
rect 26786 11568 26792 11580
rect 26844 11568 26850 11620
rect 31110 11608 31116 11620
rect 29104 11580 31116 11608
rect 24302 11540 24308 11552
rect 22066 11512 24308 11540
rect 24302 11500 24308 11512
rect 24360 11500 24366 11552
rect 24397 11543 24455 11549
rect 24397 11509 24409 11543
rect 24443 11540 24455 11543
rect 25590 11540 25596 11552
rect 24443 11512 25596 11540
rect 24443 11509 24455 11512
rect 24397 11503 24455 11509
rect 25590 11500 25596 11512
rect 25648 11500 25654 11552
rect 25774 11500 25780 11552
rect 25832 11540 25838 11552
rect 29104 11540 29132 11580
rect 31110 11568 31116 11580
rect 31168 11568 31174 11620
rect 31662 11608 31668 11620
rect 31575 11580 31668 11608
rect 31662 11568 31668 11580
rect 31720 11608 31726 11620
rect 33152 11608 33180 11784
rect 33594 11753 33600 11756
rect 33588 11707 33600 11753
rect 33594 11704 33600 11707
rect 33652 11704 33658 11756
rect 33796 11744 33824 11784
rect 33870 11772 33876 11824
rect 33928 11812 33934 11824
rect 33928 11784 36584 11812
rect 33928 11772 33934 11784
rect 35621 11747 35679 11753
rect 35621 11744 35633 11747
rect 33796 11716 35633 11744
rect 35621 11713 35633 11716
rect 35667 11744 35679 11747
rect 35802 11744 35808 11756
rect 35667 11716 35808 11744
rect 35667 11713 35679 11716
rect 35621 11707 35679 11713
rect 35802 11704 35808 11716
rect 35860 11704 35866 11756
rect 35897 11748 35955 11753
rect 35897 11747 36032 11748
rect 35897 11713 35909 11747
rect 35943 11720 36032 11747
rect 36446 11744 36452 11756
rect 35943 11713 35955 11720
rect 35897 11707 35955 11713
rect 33318 11636 33324 11688
rect 33376 11676 33382 11688
rect 36004 11676 36032 11720
rect 36407 11716 36452 11744
rect 36446 11704 36452 11716
rect 36504 11704 36510 11756
rect 36556 11753 36584 11784
rect 36541 11747 36599 11753
rect 36541 11713 36553 11747
rect 36587 11713 36599 11747
rect 36541 11707 36599 11713
rect 36722 11704 36728 11756
rect 36780 11744 36786 11756
rect 37108 11744 37136 11852
rect 37366 11840 37372 11892
rect 37424 11880 37430 11892
rect 37461 11883 37519 11889
rect 37461 11880 37473 11883
rect 37424 11852 37473 11880
rect 37424 11840 37430 11852
rect 37461 11849 37473 11852
rect 37507 11849 37519 11883
rect 43806 11880 43812 11892
rect 37461 11843 37519 11849
rect 37548 11852 43812 11880
rect 37274 11812 37280 11824
rect 37235 11784 37280 11812
rect 37274 11772 37280 11784
rect 37332 11772 37338 11824
rect 37548 11812 37576 11852
rect 43806 11840 43812 11852
rect 43864 11840 43870 11892
rect 44634 11880 44640 11892
rect 43916 11852 44640 11880
rect 37476 11784 37576 11812
rect 37476 11744 37504 11784
rect 38378 11772 38384 11824
rect 38436 11812 38442 11824
rect 38436 11784 41552 11812
rect 38436 11772 38442 11784
rect 36780 11716 36825 11744
rect 37108 11716 37504 11744
rect 37553 11747 37611 11753
rect 36780 11704 36786 11716
rect 37553 11713 37565 11747
rect 37599 11713 37611 11747
rect 39485 11747 39543 11753
rect 39485 11744 39497 11747
rect 37553 11707 37611 11713
rect 38626 11716 39497 11744
rect 36262 11676 36268 11688
rect 33376 11648 33421 11676
rect 34348 11648 36032 11676
rect 36223 11648 36268 11676
rect 33376 11636 33382 11648
rect 31720 11580 33180 11608
rect 31720 11568 31726 11580
rect 25832 11512 29132 11540
rect 25832 11500 25838 11512
rect 29178 11500 29184 11552
rect 29236 11540 29242 11552
rect 29273 11543 29331 11549
rect 29273 11540 29285 11543
rect 29236 11512 29285 11540
rect 29236 11500 29242 11512
rect 29273 11509 29285 11512
rect 29319 11509 29331 11543
rect 32582 11540 32588 11552
rect 32543 11512 32588 11540
rect 29273 11503 29331 11509
rect 32582 11500 32588 11512
rect 32640 11500 32646 11552
rect 32766 11500 32772 11552
rect 32824 11540 32830 11552
rect 34348 11540 34376 11648
rect 36262 11636 36268 11648
rect 36320 11636 36326 11688
rect 36630 11636 36636 11688
rect 36688 11676 36694 11688
rect 36688 11648 36733 11676
rect 36688 11636 36694 11648
rect 36998 11636 37004 11688
rect 37056 11676 37062 11688
rect 37568 11676 37596 11707
rect 37056 11648 37596 11676
rect 37921 11679 37979 11685
rect 37056 11636 37062 11648
rect 37921 11645 37933 11679
rect 37967 11676 37979 11679
rect 38194 11676 38200 11688
rect 37967 11648 38200 11676
rect 37967 11645 37979 11648
rect 37921 11639 37979 11645
rect 38194 11636 38200 11648
rect 38252 11676 38258 11688
rect 38470 11676 38476 11688
rect 38252 11648 38476 11676
rect 38252 11636 38258 11648
rect 38470 11636 38476 11648
rect 38528 11676 38534 11688
rect 38626 11676 38654 11716
rect 39485 11713 39497 11716
rect 39531 11713 39543 11747
rect 39485 11707 39543 11713
rect 39666 11704 39672 11756
rect 39724 11744 39730 11756
rect 40037 11747 40095 11753
rect 40037 11744 40049 11747
rect 39724 11716 40049 11744
rect 39724 11704 39730 11716
rect 40037 11713 40049 11716
rect 40083 11713 40095 11747
rect 40218 11744 40224 11756
rect 40179 11716 40224 11744
rect 40037 11707 40095 11713
rect 40218 11704 40224 11716
rect 40276 11704 40282 11756
rect 40402 11704 40408 11756
rect 40460 11744 40466 11756
rect 41141 11747 41199 11753
rect 41141 11744 41153 11747
rect 40460 11716 41153 11744
rect 40460 11704 40466 11716
rect 41141 11713 41153 11716
rect 41187 11713 41199 11747
rect 41524 11744 41552 11784
rect 41598 11772 41604 11824
rect 41656 11812 41662 11824
rect 43714 11812 43720 11824
rect 41656 11784 43720 11812
rect 41656 11772 41662 11784
rect 43714 11772 43720 11784
rect 43772 11772 43778 11824
rect 43916 11753 43944 11852
rect 44634 11840 44640 11852
rect 44692 11840 44698 11892
rect 44726 11840 44732 11892
rect 44784 11880 44790 11892
rect 46106 11880 46112 11892
rect 44784 11852 46112 11880
rect 44784 11840 44790 11852
rect 46106 11840 46112 11852
rect 46164 11840 46170 11892
rect 46201 11883 46259 11889
rect 46201 11849 46213 11883
rect 46247 11880 46259 11883
rect 46937 11883 46995 11889
rect 46937 11880 46949 11883
rect 46247 11852 46949 11880
rect 46247 11849 46259 11852
rect 46201 11843 46259 11849
rect 46937 11849 46949 11852
rect 46983 11849 46995 11883
rect 47578 11880 47584 11892
rect 47539 11852 47584 11880
rect 46937 11843 46995 11849
rect 47578 11840 47584 11852
rect 47636 11840 47642 11892
rect 47670 11840 47676 11892
rect 47728 11880 47734 11892
rect 47949 11883 48007 11889
rect 47949 11880 47961 11883
rect 47728 11852 47961 11880
rect 47728 11840 47734 11852
rect 47949 11849 47961 11852
rect 47995 11880 48007 11883
rect 48130 11880 48136 11892
rect 47995 11852 48136 11880
rect 47995 11849 48007 11852
rect 47949 11843 48007 11849
rect 48130 11840 48136 11852
rect 48188 11840 48194 11892
rect 48590 11840 48596 11892
rect 48648 11880 48654 11892
rect 49602 11880 49608 11892
rect 48648 11852 49608 11880
rect 48648 11840 48654 11852
rect 49602 11840 49608 11852
rect 49660 11840 49666 11892
rect 49789 11883 49847 11889
rect 49789 11849 49801 11883
rect 49835 11849 49847 11883
rect 49789 11843 49847 11849
rect 44085 11815 44143 11821
rect 44085 11781 44097 11815
rect 44131 11812 44143 11815
rect 44818 11812 44824 11824
rect 44131 11784 44824 11812
rect 44131 11781 44143 11784
rect 44085 11775 44143 11781
rect 44818 11772 44824 11784
rect 44876 11772 44882 11824
rect 45094 11821 45100 11824
rect 45088 11812 45100 11821
rect 45055 11784 45100 11812
rect 45088 11775 45100 11784
rect 45094 11772 45100 11775
rect 45152 11772 45158 11824
rect 45554 11772 45560 11824
rect 45612 11812 45618 11824
rect 45612 11784 47808 11812
rect 45612 11772 45618 11784
rect 43901 11747 43959 11753
rect 41524 11716 43760 11744
rect 41141 11707 41199 11713
rect 38528 11648 38654 11676
rect 38528 11636 38534 11648
rect 38930 11636 38936 11688
rect 38988 11676 38994 11688
rect 39301 11679 39359 11685
rect 39301 11676 39313 11679
rect 38988 11648 39313 11676
rect 38988 11636 38994 11648
rect 39301 11645 39313 11648
rect 39347 11645 39359 11679
rect 39301 11639 39359 11645
rect 39390 11636 39396 11688
rect 39448 11676 39454 11688
rect 39577 11679 39635 11685
rect 39448 11648 39493 11676
rect 39448 11636 39454 11648
rect 39577 11645 39589 11679
rect 39623 11676 39635 11679
rect 39850 11676 39856 11688
rect 39623 11648 39856 11676
rect 39623 11645 39635 11648
rect 39577 11639 39635 11645
rect 39850 11636 39856 11648
rect 39908 11636 39914 11688
rect 40586 11636 40592 11688
rect 40644 11676 40650 11688
rect 40770 11676 40776 11688
rect 40644 11648 40776 11676
rect 40644 11636 40650 11648
rect 40770 11636 40776 11648
rect 40828 11676 40834 11688
rect 40954 11676 40960 11688
rect 40828 11648 40960 11676
rect 40828 11636 40834 11648
rect 40954 11636 40960 11648
rect 41012 11636 41018 11688
rect 41156 11676 41184 11707
rect 43622 11676 43628 11688
rect 41156 11648 43628 11676
rect 43622 11636 43628 11648
rect 43680 11636 43686 11688
rect 43732 11676 43760 11716
rect 43901 11713 43913 11747
rect 43947 11713 43959 11747
rect 44174 11744 44180 11756
rect 44135 11716 44180 11744
rect 43901 11707 43959 11713
rect 44174 11704 44180 11716
rect 44232 11704 44238 11756
rect 44269 11748 44327 11753
rect 44358 11748 44364 11756
rect 44269 11747 44364 11748
rect 44269 11713 44281 11747
rect 44315 11720 44364 11747
rect 44315 11713 44327 11720
rect 44269 11707 44327 11713
rect 44358 11704 44364 11720
rect 44416 11704 44422 11756
rect 44468 11716 45876 11744
rect 44468 11676 44496 11716
rect 43732 11648 44496 11676
rect 44821 11679 44879 11685
rect 44821 11645 44833 11679
rect 44867 11645 44879 11679
rect 45848 11676 45876 11716
rect 46106 11704 46112 11756
rect 46164 11744 46170 11756
rect 46750 11744 46756 11756
rect 46164 11716 46756 11744
rect 46164 11704 46170 11716
rect 46750 11704 46756 11716
rect 46808 11704 46814 11756
rect 47029 11747 47087 11753
rect 47029 11713 47041 11747
rect 47075 11744 47087 11747
rect 47210 11744 47216 11756
rect 47075 11716 47216 11744
rect 47075 11713 47087 11716
rect 47029 11707 47087 11713
rect 47210 11704 47216 11716
rect 47268 11704 47274 11756
rect 47780 11753 47808 11784
rect 47854 11772 47860 11824
rect 47912 11812 47918 11824
rect 48222 11812 48228 11824
rect 47912 11784 48228 11812
rect 47912 11772 47918 11784
rect 48222 11772 48228 11784
rect 48280 11772 48286 11824
rect 49804 11812 49832 11843
rect 49878 11840 49884 11892
rect 49936 11880 49942 11892
rect 51721 11883 51779 11889
rect 49936 11852 50752 11880
rect 49936 11840 49942 11852
rect 50586 11815 50644 11821
rect 50586 11812 50598 11815
rect 49804 11784 50598 11812
rect 50586 11781 50598 11784
rect 50632 11781 50644 11815
rect 50586 11775 50644 11781
rect 47765 11747 47823 11753
rect 47765 11713 47777 11747
rect 47811 11713 47823 11747
rect 47765 11707 47823 11713
rect 48041 11747 48099 11753
rect 48041 11713 48053 11747
rect 48087 11744 48099 11747
rect 49712 11744 49832 11748
rect 48087 11720 49924 11744
rect 48087 11716 49740 11720
rect 49804 11716 49924 11720
rect 48087 11713 48099 11716
rect 48041 11707 48099 11713
rect 49510 11676 49516 11688
rect 45848 11648 49516 11676
rect 44821 11639 44879 11645
rect 35434 11608 35440 11620
rect 35395 11580 35440 11608
rect 35434 11568 35440 11580
rect 35492 11568 35498 11620
rect 36722 11568 36728 11620
rect 36780 11608 36786 11620
rect 36780 11580 37136 11608
rect 36780 11568 36786 11580
rect 32824 11512 34376 11540
rect 34701 11543 34759 11549
rect 32824 11500 32830 11512
rect 34701 11509 34713 11543
rect 34747 11540 34759 11543
rect 35986 11540 35992 11552
rect 34747 11512 35992 11540
rect 34747 11509 34759 11512
rect 34701 11503 34759 11509
rect 35986 11500 35992 11512
rect 36044 11500 36050 11552
rect 36170 11500 36176 11552
rect 36228 11540 36234 11552
rect 36906 11540 36912 11552
rect 36228 11512 36912 11540
rect 36228 11500 36234 11512
rect 36906 11500 36912 11512
rect 36964 11500 36970 11552
rect 37108 11540 37136 11580
rect 37182 11568 37188 11620
rect 37240 11608 37246 11620
rect 37277 11611 37335 11617
rect 37277 11608 37289 11611
rect 37240 11580 37289 11608
rect 37240 11568 37246 11580
rect 37277 11577 37289 11580
rect 37323 11577 37335 11611
rect 37277 11571 37335 11577
rect 37366 11568 37372 11620
rect 37424 11608 37430 11620
rect 37550 11608 37556 11620
rect 37424 11580 37556 11608
rect 37424 11568 37430 11580
rect 37550 11568 37556 11580
rect 37608 11608 37614 11620
rect 38286 11608 38292 11620
rect 37608 11580 38292 11608
rect 37608 11568 37614 11580
rect 38286 11568 38292 11580
rect 38344 11568 38350 11620
rect 38746 11568 38752 11620
rect 38804 11608 38810 11620
rect 44082 11608 44088 11620
rect 38804 11580 44088 11608
rect 38804 11568 38810 11580
rect 44082 11568 44088 11580
rect 44140 11568 44146 11620
rect 38151 11543 38209 11549
rect 38151 11540 38163 11543
rect 37108 11512 38163 11540
rect 38151 11509 38163 11512
rect 38197 11540 38209 11543
rect 39022 11540 39028 11552
rect 38197 11512 39028 11540
rect 38197 11509 38209 11512
rect 38151 11503 38209 11509
rect 39022 11500 39028 11512
rect 39080 11500 39086 11552
rect 39117 11543 39175 11549
rect 39117 11509 39129 11543
rect 39163 11540 39175 11543
rect 40310 11540 40316 11552
rect 39163 11512 40316 11540
rect 39163 11509 39175 11512
rect 39117 11503 39175 11509
rect 40310 11500 40316 11512
rect 40368 11500 40374 11552
rect 40405 11543 40463 11549
rect 40405 11509 40417 11543
rect 40451 11540 40463 11543
rect 40770 11540 40776 11552
rect 40451 11512 40776 11540
rect 40451 11509 40463 11512
rect 40405 11503 40463 11509
rect 40770 11500 40776 11512
rect 40828 11500 40834 11552
rect 41138 11500 41144 11552
rect 41196 11540 41202 11552
rect 41371 11543 41429 11549
rect 41371 11540 41383 11543
rect 41196 11512 41383 11540
rect 41196 11500 41202 11512
rect 41371 11509 41383 11512
rect 41417 11540 41429 11543
rect 44174 11540 44180 11552
rect 41417 11512 44180 11540
rect 41417 11509 41429 11512
rect 41371 11503 41429 11509
rect 44174 11500 44180 11512
rect 44232 11500 44238 11552
rect 44450 11540 44456 11552
rect 44411 11512 44456 11540
rect 44450 11500 44456 11512
rect 44508 11500 44514 11552
rect 44836 11540 44864 11639
rect 49510 11636 49516 11648
rect 49568 11636 49574 11688
rect 49896 11676 49924 11716
rect 49970 11704 49976 11756
rect 50028 11744 50034 11756
rect 50338 11744 50344 11756
rect 50028 11716 50073 11744
rect 50299 11716 50344 11744
rect 50028 11704 50034 11716
rect 50338 11704 50344 11716
rect 50396 11704 50402 11756
rect 50724 11744 50752 11852
rect 51721 11849 51733 11883
rect 51767 11849 51779 11883
rect 52086 11880 52092 11892
rect 52047 11852 52092 11880
rect 51721 11843 51779 11849
rect 51074 11772 51080 11824
rect 51132 11812 51138 11824
rect 51736 11812 51764 11843
rect 52086 11840 52092 11852
rect 52144 11840 52150 11892
rect 52730 11880 52736 11892
rect 52196 11852 52500 11880
rect 52691 11852 52736 11880
rect 52196 11812 52224 11852
rect 51132 11784 51479 11812
rect 51736 11784 52224 11812
rect 52472 11812 52500 11852
rect 52730 11840 52736 11852
rect 52788 11840 52794 11892
rect 53190 11840 53196 11892
rect 53248 11840 53254 11892
rect 53374 11840 53380 11892
rect 53432 11880 53438 11892
rect 54662 11880 54668 11892
rect 53432 11852 54668 11880
rect 53432 11840 53438 11852
rect 54662 11840 54668 11852
rect 54720 11840 54726 11892
rect 54754 11840 54760 11892
rect 54812 11880 54818 11892
rect 55401 11883 55459 11889
rect 55401 11880 55413 11883
rect 54812 11852 55413 11880
rect 54812 11840 54818 11852
rect 55401 11849 55413 11852
rect 55447 11849 55459 11883
rect 55401 11843 55459 11849
rect 55861 11883 55919 11889
rect 55861 11849 55873 11883
rect 55907 11880 55919 11883
rect 56502 11880 56508 11892
rect 55907 11852 56508 11880
rect 55907 11849 55919 11852
rect 55861 11843 55919 11849
rect 56502 11840 56508 11852
rect 56560 11840 56566 11892
rect 56842 11852 60504 11880
rect 53101 11815 53159 11821
rect 53101 11812 53113 11815
rect 52472 11784 53113 11812
rect 51132 11772 51138 11784
rect 51350 11744 51356 11756
rect 50724 11716 51356 11744
rect 51350 11704 51356 11716
rect 51408 11704 51414 11756
rect 51451 11676 51479 11784
rect 53101 11781 53113 11784
rect 53147 11781 53159 11815
rect 53101 11775 53159 11781
rect 53218 11812 53246 11840
rect 53218 11784 54064 11812
rect 51994 11704 52000 11756
rect 52052 11744 52058 11756
rect 52265 11747 52323 11753
rect 52265 11744 52277 11747
rect 52052 11716 52277 11744
rect 52052 11704 52058 11716
rect 52265 11713 52277 11716
rect 52311 11713 52323 11747
rect 52265 11707 52323 11713
rect 52822 11704 52828 11756
rect 52880 11744 52886 11756
rect 53218 11753 53246 11784
rect 52917 11747 52975 11753
rect 52917 11744 52929 11747
rect 52880 11716 52929 11744
rect 52880 11704 52886 11716
rect 52917 11713 52929 11716
rect 52963 11713 52975 11747
rect 52917 11707 52975 11713
rect 53203 11747 53261 11753
rect 53203 11713 53215 11747
rect 53249 11713 53261 11747
rect 53742 11744 53748 11756
rect 53703 11716 53748 11744
rect 53203 11707 53261 11713
rect 53742 11704 53748 11716
rect 53800 11704 53806 11756
rect 53926 11744 53932 11756
rect 53887 11716 53932 11744
rect 53926 11704 53932 11716
rect 53984 11704 53990 11756
rect 54036 11753 54064 11784
rect 54202 11772 54208 11824
rect 54260 11812 54266 11824
rect 54573 11815 54631 11821
rect 54573 11812 54585 11815
rect 54260 11784 54585 11812
rect 54260 11772 54266 11784
rect 54573 11781 54585 11784
rect 54619 11781 54631 11815
rect 56842 11812 56870 11852
rect 56962 11812 56968 11824
rect 54573 11775 54631 11781
rect 54660 11784 56870 11812
rect 56923 11784 56968 11812
rect 54021 11747 54079 11753
rect 54021 11713 54033 11747
rect 54067 11744 54079 11747
rect 54110 11744 54116 11756
rect 54067 11716 54116 11744
rect 54067 11713 54079 11716
rect 54021 11707 54079 11713
rect 54110 11704 54116 11716
rect 54168 11704 54174 11756
rect 54660 11744 54688 11784
rect 56962 11772 56968 11784
rect 57020 11772 57026 11824
rect 57054 11772 57060 11824
rect 57112 11812 57118 11824
rect 57425 11815 57483 11821
rect 57425 11812 57437 11815
rect 57112 11784 57437 11812
rect 57112 11772 57118 11784
rect 57425 11781 57437 11784
rect 57471 11781 57483 11815
rect 57425 11775 57483 11781
rect 57514 11772 57520 11824
rect 57572 11812 57578 11824
rect 58894 11812 58900 11824
rect 57572 11784 58664 11812
rect 58855 11784 58900 11812
rect 57572 11772 57578 11784
rect 54220 11716 54688 11744
rect 54849 11747 54907 11753
rect 54220 11676 54248 11716
rect 54849 11713 54861 11747
rect 54895 11744 54907 11747
rect 55214 11744 55220 11756
rect 54895 11716 54984 11744
rect 55175 11716 55220 11744
rect 54895 11713 54907 11716
rect 54849 11707 54907 11713
rect 49896 11648 50108 11676
rect 51451 11648 54248 11676
rect 54645 11679 54703 11685
rect 46106 11568 46112 11620
rect 46164 11608 46170 11620
rect 49878 11608 49884 11620
rect 46164 11580 49884 11608
rect 46164 11568 46170 11580
rect 49878 11568 49884 11580
rect 49936 11568 49942 11620
rect 50080 11608 50108 11648
rect 54645 11645 54657 11679
rect 54691 11676 54703 11679
rect 54754 11676 54760 11688
rect 54691 11648 54760 11676
rect 54691 11645 54703 11648
rect 54645 11639 54703 11645
rect 54754 11636 54760 11648
rect 54812 11636 54818 11688
rect 54956 11676 54984 11716
rect 55214 11704 55220 11716
rect 55272 11704 55278 11756
rect 55493 11747 55551 11753
rect 55493 11713 55505 11747
rect 55539 11713 55551 11747
rect 55493 11707 55551 11713
rect 55122 11676 55128 11688
rect 54956 11648 55128 11676
rect 55122 11636 55128 11648
rect 55180 11636 55186 11688
rect 55508 11676 55536 11707
rect 55766 11704 55772 11756
rect 55824 11744 55830 11756
rect 56045 11747 56103 11753
rect 56045 11744 56057 11747
rect 55824 11716 56057 11744
rect 55824 11704 55830 11716
rect 56045 11713 56057 11716
rect 56091 11713 56103 11747
rect 57146 11744 57152 11756
rect 57107 11716 57152 11744
rect 56045 11707 56103 11713
rect 57146 11704 57152 11716
rect 57204 11704 57210 11756
rect 57333 11747 57391 11753
rect 57333 11713 57345 11747
rect 57379 11713 57391 11747
rect 57882 11744 57888 11756
rect 57843 11716 57888 11744
rect 57333 11707 57391 11713
rect 56502 11676 56508 11688
rect 55508 11648 56508 11676
rect 56502 11636 56508 11648
rect 56560 11636 56566 11688
rect 57348 11676 57376 11707
rect 57882 11704 57888 11716
rect 57940 11704 57946 11756
rect 58069 11747 58127 11753
rect 58069 11713 58081 11747
rect 58115 11744 58127 11747
rect 58342 11744 58348 11756
rect 58115 11716 58348 11744
rect 58115 11713 58127 11716
rect 58069 11707 58127 11713
rect 58342 11704 58348 11716
rect 58400 11704 58406 11756
rect 58636 11753 58664 11784
rect 58894 11772 58900 11784
rect 58952 11772 58958 11824
rect 59170 11772 59176 11824
rect 59228 11812 59234 11824
rect 60476 11812 60504 11852
rect 60550 11840 60556 11892
rect 60608 11880 60614 11892
rect 61102 11880 61108 11892
rect 60608 11852 61108 11880
rect 60608 11840 60614 11852
rect 61102 11840 61108 11852
rect 61160 11840 61166 11892
rect 61194 11840 61200 11892
rect 61252 11880 61258 11892
rect 64601 11883 64659 11889
rect 64601 11880 64613 11883
rect 61252 11852 63724 11880
rect 61252 11840 61258 11852
rect 59228 11784 60228 11812
rect 60476 11784 62896 11812
rect 59228 11772 59234 11784
rect 59078 11753 59084 11756
rect 58621 11747 58679 11753
rect 58621 11713 58633 11747
rect 58667 11713 58679 11747
rect 58621 11707 58679 11713
rect 58805 11747 58863 11753
rect 58805 11713 58817 11747
rect 58851 11713 58863 11747
rect 58805 11707 58863 11713
rect 59041 11747 59084 11753
rect 59041 11713 59053 11747
rect 59041 11707 59084 11713
rect 58526 11676 58532 11688
rect 57348 11648 58532 11676
rect 58526 11636 58532 11648
rect 58584 11636 58590 11688
rect 58820 11676 58848 11707
rect 59078 11704 59084 11707
rect 59136 11704 59142 11756
rect 59354 11704 59360 11756
rect 59412 11744 59418 11756
rect 59817 11747 59875 11753
rect 59817 11744 59829 11747
rect 59412 11716 59829 11744
rect 59412 11704 59418 11716
rect 59817 11713 59829 11716
rect 59863 11713 59875 11747
rect 59998 11744 60004 11756
rect 59959 11716 60004 11744
rect 59817 11707 59875 11713
rect 59998 11704 60004 11716
rect 60056 11704 60062 11756
rect 60093 11748 60151 11753
rect 60200 11748 60228 11784
rect 60093 11747 60228 11748
rect 60093 11713 60105 11747
rect 60139 11720 60228 11747
rect 61096 11747 61154 11753
rect 60139 11713 60151 11720
rect 60093 11707 60151 11713
rect 61096 11713 61108 11747
rect 61142 11744 61154 11747
rect 62868 11744 62896 11784
rect 62942 11772 62948 11824
rect 63000 11812 63006 11824
rect 63037 11815 63095 11821
rect 63037 11812 63049 11815
rect 63000 11784 63049 11812
rect 63000 11772 63006 11784
rect 63037 11781 63049 11784
rect 63083 11812 63095 11815
rect 63586 11812 63592 11824
rect 63083 11784 63592 11812
rect 63083 11781 63095 11784
rect 63037 11775 63095 11781
rect 63586 11772 63592 11784
rect 63644 11772 63650 11824
rect 63402 11744 63408 11756
rect 61142 11716 62068 11744
rect 62868 11716 63408 11744
rect 61142 11713 61154 11716
rect 61096 11707 61154 11713
rect 59633 11679 59691 11685
rect 59633 11676 59645 11679
rect 58820 11648 59645 11676
rect 59633 11645 59645 11648
rect 59679 11645 59691 11679
rect 60826 11676 60832 11688
rect 60787 11648 60832 11676
rect 59633 11639 59691 11645
rect 60826 11636 60832 11648
rect 60884 11636 60890 11688
rect 62040 11676 62068 11716
rect 63402 11704 63408 11716
rect 63460 11704 63466 11756
rect 62114 11676 62120 11688
rect 62040 11648 62120 11676
rect 62114 11636 62120 11648
rect 62172 11636 62178 11688
rect 63586 11676 63592 11688
rect 63547 11648 63592 11676
rect 63586 11636 63592 11648
rect 63644 11636 63650 11688
rect 63696 11676 63724 11852
rect 63880 11852 64613 11880
rect 63880 11753 63908 11852
rect 64601 11849 64613 11852
rect 64647 11880 64659 11883
rect 64782 11880 64788 11892
rect 64647 11852 64788 11880
rect 64647 11849 64659 11852
rect 64601 11843 64659 11849
rect 64782 11840 64788 11852
rect 64840 11840 64846 11892
rect 64874 11840 64880 11892
rect 64932 11880 64938 11892
rect 66806 11880 66812 11892
rect 64932 11852 66812 11880
rect 64932 11840 64938 11852
rect 66806 11840 66812 11852
rect 66864 11840 66870 11892
rect 66901 11883 66959 11889
rect 66901 11849 66913 11883
rect 66947 11880 66959 11883
rect 67174 11880 67180 11892
rect 66947 11852 67180 11880
rect 66947 11849 66959 11852
rect 66901 11843 66959 11849
rect 67174 11840 67180 11852
rect 67232 11840 67238 11892
rect 67266 11840 67272 11892
rect 67324 11840 67330 11892
rect 67542 11840 67548 11892
rect 67600 11880 67606 11892
rect 69106 11880 69112 11892
rect 67600 11852 69112 11880
rect 67600 11840 67606 11852
rect 69106 11840 69112 11852
rect 69164 11840 69170 11892
rect 69198 11840 69204 11892
rect 69256 11880 69262 11892
rect 69842 11880 69848 11892
rect 69256 11852 69848 11880
rect 69256 11840 69262 11852
rect 69842 11840 69848 11852
rect 69900 11840 69906 11892
rect 70026 11840 70032 11892
rect 70084 11880 70090 11892
rect 70581 11883 70639 11889
rect 70581 11880 70593 11883
rect 70084 11852 70593 11880
rect 70084 11840 70090 11852
rect 70581 11849 70593 11852
rect 70627 11849 70639 11883
rect 70581 11843 70639 11849
rect 71225 11883 71283 11889
rect 71225 11849 71237 11883
rect 71271 11880 71283 11883
rect 71314 11880 71320 11892
rect 71271 11852 71320 11880
rect 71271 11849 71283 11852
rect 71225 11843 71283 11849
rect 71314 11840 71320 11852
rect 71372 11840 71378 11892
rect 71593 11883 71651 11889
rect 71593 11849 71605 11883
rect 71639 11880 71651 11883
rect 72326 11880 72332 11892
rect 71639 11852 72332 11880
rect 71639 11849 71651 11852
rect 71593 11843 71651 11849
rect 72326 11840 72332 11852
rect 72384 11840 72390 11892
rect 64417 11815 64475 11821
rect 64417 11781 64429 11815
rect 64463 11812 64475 11815
rect 65150 11812 65156 11824
rect 64463 11784 65156 11812
rect 64463 11781 64475 11784
rect 64417 11775 64475 11781
rect 65150 11772 65156 11784
rect 65208 11772 65214 11824
rect 66990 11812 66996 11824
rect 65260 11784 66996 11812
rect 63865 11747 63923 11753
rect 63865 11713 63877 11747
rect 63911 11713 63923 11747
rect 64046 11744 64052 11756
rect 64007 11716 64052 11744
rect 63865 11707 63923 11713
rect 64046 11704 64052 11716
rect 64104 11704 64110 11756
rect 64690 11744 64696 11756
rect 64651 11716 64696 11744
rect 64690 11704 64696 11716
rect 64748 11704 64754 11756
rect 65260 11676 65288 11784
rect 66990 11772 66996 11784
rect 67048 11772 67054 11824
rect 66162 11744 66168 11756
rect 66123 11716 66168 11744
rect 66162 11704 66168 11716
rect 66220 11704 66226 11756
rect 66254 11704 66260 11756
rect 66312 11744 66318 11756
rect 66349 11747 66407 11753
rect 66349 11744 66361 11747
rect 66312 11716 66361 11744
rect 66312 11704 66318 11716
rect 66349 11713 66361 11716
rect 66395 11713 66407 11747
rect 66349 11707 66407 11713
rect 66533 11747 66591 11753
rect 66533 11713 66545 11747
rect 66579 11744 66591 11747
rect 67085 11747 67143 11753
rect 67085 11744 67097 11747
rect 66579 11716 67097 11744
rect 66579 11713 66591 11716
rect 66533 11707 66591 11713
rect 67085 11713 67097 11716
rect 67131 11713 67143 11747
rect 67085 11707 67143 11713
rect 63696 11648 65288 11676
rect 66180 11676 66208 11704
rect 67284 11676 67312 11840
rect 68830 11772 68836 11824
rect 68888 11812 68894 11824
rect 69446 11815 69504 11821
rect 69446 11812 69458 11815
rect 68888 11784 69458 11812
rect 68888 11772 68894 11784
rect 69446 11781 69458 11784
rect 69492 11781 69504 11815
rect 70854 11812 70860 11824
rect 70815 11784 70860 11812
rect 69446 11775 69504 11781
rect 70854 11772 70860 11784
rect 70912 11772 70918 11824
rect 67358 11704 67364 11756
rect 67416 11744 67422 11756
rect 68373 11747 68431 11753
rect 67416 11716 68324 11744
rect 67416 11704 67422 11716
rect 66180 11648 67312 11676
rect 67542 11636 67548 11688
rect 67600 11676 67606 11688
rect 68189 11679 68247 11685
rect 68189 11676 68201 11679
rect 67600 11648 68201 11676
rect 67600 11636 67606 11648
rect 68189 11645 68201 11648
rect 68235 11645 68247 11679
rect 68296 11676 68324 11716
rect 68373 11713 68385 11747
rect 68419 11744 68431 11747
rect 68922 11744 68928 11756
rect 68419 11716 68928 11744
rect 68419 11713 68431 11716
rect 68373 11707 68431 11713
rect 68922 11704 68928 11716
rect 68980 11704 68986 11756
rect 69106 11744 69112 11756
rect 69067 11716 69112 11744
rect 69106 11704 69112 11716
rect 69164 11704 69170 11756
rect 69198 11704 69204 11756
rect 69256 11744 69262 11756
rect 70872 11744 70900 11772
rect 71498 11744 71504 11756
rect 69256 11716 69301 11744
rect 70872 11716 71504 11744
rect 69256 11704 69262 11716
rect 71498 11704 71504 11716
rect 71556 11744 71562 11756
rect 88242 11744 88248 11756
rect 71556 11716 71820 11744
rect 88203 11716 88248 11744
rect 71556 11704 71562 11716
rect 68296 11648 69060 11676
rect 68189 11639 68247 11645
rect 50246 11608 50252 11620
rect 50080 11580 50252 11608
rect 50246 11568 50252 11580
rect 50304 11568 50310 11620
rect 51276 11580 56732 11608
rect 51276 11552 51304 11580
rect 45738 11540 45744 11552
rect 44836 11512 45744 11540
rect 45738 11500 45744 11512
rect 45796 11500 45802 11552
rect 45830 11500 45836 11552
rect 45888 11540 45894 11552
rect 46569 11543 46627 11549
rect 46569 11540 46581 11543
rect 45888 11512 46581 11540
rect 45888 11500 45894 11512
rect 46569 11509 46581 11512
rect 46615 11509 46627 11543
rect 46569 11503 46627 11509
rect 47578 11500 47584 11552
rect 47636 11540 47642 11552
rect 51074 11540 51080 11552
rect 47636 11512 51080 11540
rect 47636 11500 47642 11512
rect 51074 11500 51080 11512
rect 51132 11500 51138 11552
rect 51258 11500 51264 11552
rect 51316 11500 51322 11552
rect 51350 11500 51356 11552
rect 51408 11540 51414 11552
rect 52914 11540 52920 11552
rect 51408 11512 52920 11540
rect 51408 11500 51414 11512
rect 52914 11500 52920 11512
rect 52972 11500 52978 11552
rect 53098 11500 53104 11552
rect 53156 11540 53162 11552
rect 53561 11543 53619 11549
rect 53561 11540 53573 11543
rect 53156 11512 53573 11540
rect 53156 11500 53162 11512
rect 53561 11509 53573 11512
rect 53607 11509 53619 11543
rect 53561 11503 53619 11509
rect 54110 11500 54116 11552
rect 54168 11540 54174 11552
rect 54846 11540 54852 11552
rect 54168 11512 54852 11540
rect 54168 11500 54174 11512
rect 54846 11500 54852 11512
rect 54904 11500 54910 11552
rect 55217 11543 55275 11549
rect 55217 11509 55229 11543
rect 55263 11540 55275 11543
rect 56594 11540 56600 11552
rect 55263 11512 56600 11540
rect 55263 11509 55275 11512
rect 55217 11503 55275 11509
rect 56594 11500 56600 11512
rect 56652 11500 56658 11552
rect 56704 11540 56732 11580
rect 57146 11568 57152 11620
rect 57204 11608 57210 11620
rect 58066 11608 58072 11620
rect 57204 11580 58072 11608
rect 57204 11568 57210 11580
rect 58066 11568 58072 11580
rect 58124 11568 58130 11620
rect 58253 11611 58311 11617
rect 58253 11577 58265 11611
rect 58299 11608 58311 11611
rect 60550 11608 60556 11620
rect 58299 11580 60556 11608
rect 58299 11577 58311 11580
rect 58253 11571 58311 11577
rect 60550 11568 60556 11580
rect 60608 11568 60614 11620
rect 61930 11568 61936 11620
rect 61988 11608 61994 11620
rect 67174 11608 67180 11620
rect 61988 11580 67180 11608
rect 61988 11568 61994 11580
rect 67174 11568 67180 11580
rect 67232 11568 67238 11620
rect 67266 11568 67272 11620
rect 67324 11608 67330 11620
rect 68925 11611 68983 11617
rect 68925 11608 68937 11611
rect 67324 11580 68937 11608
rect 67324 11568 67330 11580
rect 68925 11577 68937 11580
rect 68971 11577 68983 11611
rect 68925 11571 68983 11577
rect 58894 11540 58900 11552
rect 56704 11512 58900 11540
rect 58894 11500 58900 11512
rect 58952 11500 58958 11552
rect 59170 11540 59176 11552
rect 59131 11512 59176 11540
rect 59170 11500 59176 11512
rect 59228 11500 59234 11552
rect 59262 11500 59268 11552
rect 59320 11540 59326 11552
rect 61194 11540 61200 11552
rect 59320 11512 61200 11540
rect 59320 11500 59326 11512
rect 61194 11500 61200 11512
rect 61252 11500 61258 11552
rect 61470 11500 61476 11552
rect 61528 11540 61534 11552
rect 62209 11543 62267 11549
rect 62209 11540 62221 11543
rect 61528 11512 62221 11540
rect 61528 11500 61534 11512
rect 62209 11509 62221 11512
rect 62255 11540 62267 11543
rect 62298 11540 62304 11552
rect 62255 11512 62304 11540
rect 62255 11509 62267 11512
rect 62209 11503 62267 11509
rect 62298 11500 62304 11512
rect 62356 11500 62362 11552
rect 63218 11500 63224 11552
rect 63276 11540 63282 11552
rect 64417 11543 64475 11549
rect 64417 11540 64429 11543
rect 63276 11512 64429 11540
rect 63276 11500 63282 11512
rect 64417 11509 64429 11512
rect 64463 11509 64475 11543
rect 64417 11503 64475 11509
rect 64690 11500 64696 11552
rect 64748 11540 64754 11552
rect 67082 11540 67088 11552
rect 64748 11512 67088 11540
rect 64748 11500 64754 11512
rect 67082 11500 67088 11512
rect 67140 11540 67146 11552
rect 68557 11543 68615 11549
rect 68557 11540 68569 11543
rect 67140 11512 68569 11540
rect 67140 11500 67146 11512
rect 68557 11509 68569 11512
rect 68603 11509 68615 11543
rect 69032 11540 69060 11648
rect 71406 11636 71412 11688
rect 71464 11676 71470 11688
rect 71792 11685 71820 11716
rect 88242 11704 88248 11716
rect 88300 11704 88306 11756
rect 71685 11679 71743 11685
rect 71685 11676 71697 11679
rect 71464 11648 71697 11676
rect 71464 11636 71470 11648
rect 71685 11645 71697 11648
rect 71731 11645 71743 11679
rect 71685 11639 71743 11645
rect 71777 11679 71835 11685
rect 71777 11645 71789 11679
rect 71823 11645 71835 11679
rect 71777 11639 71835 11645
rect 88058 11608 88064 11620
rect 88019 11580 88064 11608
rect 88058 11568 88064 11580
rect 88116 11568 88122 11620
rect 70394 11540 70400 11552
rect 69032 11512 70400 11540
rect 68557 11503 68615 11509
rect 70394 11500 70400 11512
rect 70452 11500 70458 11552
rect 1104 11450 88872 11472
rect 1104 11398 11924 11450
rect 11976 11398 11988 11450
rect 12040 11398 12052 11450
rect 12104 11398 12116 11450
rect 12168 11398 12180 11450
rect 12232 11398 33872 11450
rect 33924 11398 33936 11450
rect 33988 11398 34000 11450
rect 34052 11398 34064 11450
rect 34116 11398 34128 11450
rect 34180 11398 55820 11450
rect 55872 11398 55884 11450
rect 55936 11398 55948 11450
rect 56000 11398 56012 11450
rect 56064 11398 56076 11450
rect 56128 11398 77768 11450
rect 77820 11398 77832 11450
rect 77884 11398 77896 11450
rect 77948 11398 77960 11450
rect 78012 11398 78024 11450
rect 78076 11398 88872 11450
rect 1104 11376 88872 11398
rect 4798 11296 4804 11348
rect 4856 11336 4862 11348
rect 14458 11336 14464 11348
rect 4856 11308 14464 11336
rect 4856 11296 4862 11308
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 15565 11339 15623 11345
rect 15565 11336 15577 11339
rect 14792 11308 15577 11336
rect 14792 11296 14798 11308
rect 15565 11305 15577 11308
rect 15611 11305 15623 11339
rect 24486 11336 24492 11348
rect 15565 11299 15623 11305
rect 19306 11308 24492 11336
rect 19306 11268 19334 11308
rect 24486 11296 24492 11308
rect 24544 11296 24550 11348
rect 24854 11336 24860 11348
rect 24815 11308 24860 11336
rect 24854 11296 24860 11308
rect 24912 11296 24918 11348
rect 27614 11336 27620 11348
rect 27575 11308 27620 11336
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 34238 11336 34244 11348
rect 27724 11308 34100 11336
rect 34199 11308 34244 11336
rect 25314 11268 25320 11280
rect 6886 11240 19334 11268
rect 25275 11240 25320 11268
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 6886 11132 6914 11240
rect 25314 11228 25320 11240
rect 25372 11228 25378 11280
rect 26878 11228 26884 11280
rect 26936 11268 26942 11280
rect 27724 11268 27752 11308
rect 29546 11268 29552 11280
rect 26936 11240 27752 11268
rect 27816 11240 29552 11268
rect 26936 11228 26942 11240
rect 18782 11160 18788 11212
rect 18840 11200 18846 11212
rect 23474 11200 23480 11212
rect 18840 11172 23480 11200
rect 18840 11160 18846 11172
rect 23474 11160 23480 11172
rect 23532 11160 23538 11212
rect 23566 11160 23572 11212
rect 23624 11200 23630 11212
rect 27816 11200 27844 11240
rect 29546 11228 29552 11240
rect 29604 11228 29610 11280
rect 31018 11228 31024 11280
rect 31076 11268 31082 11280
rect 32125 11271 32183 11277
rect 32125 11268 32137 11271
rect 31076 11240 32137 11268
rect 31076 11228 31082 11240
rect 32125 11237 32137 11240
rect 32171 11237 32183 11271
rect 34072 11268 34100 11308
rect 34238 11296 34244 11308
rect 34296 11296 34302 11348
rect 35621 11339 35679 11345
rect 35621 11305 35633 11339
rect 35667 11336 35679 11339
rect 35710 11336 35716 11348
rect 35667 11308 35716 11336
rect 35667 11305 35679 11308
rect 35621 11299 35679 11305
rect 35710 11296 35716 11308
rect 35768 11296 35774 11348
rect 35802 11296 35808 11348
rect 35860 11336 35866 11348
rect 38562 11336 38568 11348
rect 35860 11308 38568 11336
rect 35860 11296 35866 11308
rect 38562 11296 38568 11308
rect 38620 11296 38626 11348
rect 38746 11336 38752 11348
rect 38707 11308 38752 11336
rect 38746 11296 38752 11308
rect 38804 11296 38810 11348
rect 38838 11296 38844 11348
rect 38896 11296 38902 11348
rect 39850 11336 39856 11348
rect 39811 11308 39856 11336
rect 39850 11296 39856 11308
rect 39908 11296 39914 11348
rect 40126 11296 40132 11348
rect 40184 11336 40190 11348
rect 41138 11336 41144 11348
rect 40184 11308 41144 11336
rect 40184 11296 40190 11308
rect 41138 11296 41144 11308
rect 41196 11296 41202 11348
rect 41230 11296 41236 11348
rect 41288 11336 41294 11348
rect 42337 11339 42395 11345
rect 42337 11336 42349 11339
rect 41288 11308 42349 11336
rect 41288 11296 41294 11308
rect 42337 11305 42349 11308
rect 42383 11305 42395 11339
rect 44726 11336 44732 11348
rect 42337 11299 42395 11305
rect 44013 11308 44732 11336
rect 38856 11268 38884 11296
rect 34072 11240 38884 11268
rect 32125 11231 32183 11237
rect 39022 11228 39028 11280
rect 39080 11268 39086 11280
rect 39080 11240 39160 11268
rect 39080 11228 39086 11240
rect 29454 11200 29460 11212
rect 23624 11172 25912 11200
rect 23624 11160 23630 11172
rect 1627 11104 6914 11132
rect 15289 11135 15347 11141
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 15289 11101 15301 11135
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 15304 11064 15332 11095
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 15436 11104 15481 11132
rect 15436 11092 15442 11104
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 24210 11132 24216 11144
rect 15896 11104 24216 11132
rect 15896 11092 15902 11104
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 24397 11135 24455 11141
rect 24397 11101 24409 11135
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24302 11064 24308 11076
rect 15304 11036 24308 11064
rect 24302 11024 24308 11036
rect 24360 11024 24366 11076
rect 24412 11064 24440 11095
rect 24578 11092 24584 11144
rect 24636 11132 24642 11144
rect 25225 11135 25283 11141
rect 25225 11132 25237 11135
rect 24636 11104 25237 11132
rect 24636 11092 24642 11104
rect 25225 11101 25237 11104
rect 25271 11101 25283 11135
rect 25774 11132 25780 11144
rect 25735 11104 25780 11132
rect 25225 11095 25283 11101
rect 25774 11092 25780 11104
rect 25832 11092 25838 11144
rect 25884 11132 25912 11172
rect 26896 11172 27844 11200
rect 29012 11172 29460 11200
rect 26896 11132 26924 11172
rect 25884 11104 26924 11132
rect 27154 11092 27160 11144
rect 27212 11132 27218 11144
rect 27801 11135 27859 11141
rect 27801 11132 27813 11135
rect 27212 11104 27813 11132
rect 27212 11092 27218 11104
rect 27801 11101 27813 11104
rect 27847 11101 27859 11135
rect 29012 11132 29040 11172
rect 29454 11160 29460 11172
rect 29512 11160 29518 11212
rect 34701 11203 34759 11209
rect 34701 11169 34713 11203
rect 34747 11200 34759 11203
rect 34974 11200 34980 11212
rect 34747 11172 34980 11200
rect 34747 11169 34759 11172
rect 34701 11163 34759 11169
rect 34974 11160 34980 11172
rect 35032 11160 35038 11212
rect 36538 11200 36544 11212
rect 35820 11172 36544 11200
rect 27801 11095 27859 11101
rect 28828 11104 29040 11132
rect 29089 11135 29147 11141
rect 24412 11036 24900 11064
rect 1394 10996 1400 11008
rect 1355 10968 1400 10996
rect 1394 10956 1400 10968
rect 1452 10956 1458 11008
rect 24872 10996 24900 11036
rect 25038 11024 25044 11076
rect 25096 11064 25102 11076
rect 26022 11067 26080 11073
rect 26022 11064 26034 11067
rect 25096 11036 26034 11064
rect 25096 11024 25102 11036
rect 26022 11033 26034 11036
rect 26068 11033 26080 11067
rect 26022 11027 26080 11033
rect 26234 11024 26240 11076
rect 26292 11064 26298 11076
rect 28828 11064 28856 11104
rect 29089 11101 29101 11135
rect 29135 11132 29147 11135
rect 29178 11132 29184 11144
rect 29135 11104 29184 11132
rect 29135 11101 29147 11104
rect 29089 11095 29147 11101
rect 29178 11092 29184 11104
rect 29236 11092 29242 11144
rect 29546 11132 29552 11144
rect 29507 11104 29552 11132
rect 29546 11092 29552 11104
rect 29604 11092 29610 11144
rect 30742 11092 30748 11144
rect 30800 11132 30806 11144
rect 31754 11132 31760 11144
rect 30800 11104 31760 11132
rect 30800 11092 30806 11104
rect 31754 11092 31760 11104
rect 31812 11132 31818 11144
rect 31941 11135 31999 11141
rect 31812 11104 31857 11132
rect 31812 11092 31818 11104
rect 31941 11101 31953 11135
rect 31987 11132 31999 11135
rect 32490 11132 32496 11144
rect 31987 11104 32496 11132
rect 31987 11101 31999 11104
rect 31941 11095 31999 11101
rect 32490 11092 32496 11104
rect 32548 11092 32554 11144
rect 32861 11135 32919 11141
rect 32861 11101 32873 11135
rect 32907 11132 32919 11135
rect 34885 11135 34943 11141
rect 32907 11104 33272 11132
rect 32907 11101 32919 11104
rect 32861 11095 32919 11101
rect 33244 11076 33272 11104
rect 34885 11101 34897 11135
rect 34931 11132 34943 11135
rect 35710 11132 35716 11144
rect 34931 11104 35716 11132
rect 34931 11101 34943 11104
rect 34885 11095 34943 11101
rect 35710 11092 35716 11104
rect 35768 11092 35774 11144
rect 35820 11141 35848 11172
rect 36538 11160 36544 11172
rect 36596 11160 36602 11212
rect 36633 11203 36691 11209
rect 36633 11169 36645 11203
rect 36679 11200 36691 11203
rect 37734 11200 37740 11212
rect 36679 11172 37740 11200
rect 36679 11169 36691 11172
rect 36633 11163 36691 11169
rect 37734 11160 37740 11172
rect 37792 11160 37798 11212
rect 38194 11160 38200 11212
rect 38252 11200 38258 11212
rect 38252 11172 38297 11200
rect 38252 11160 38258 11172
rect 38470 11160 38476 11212
rect 38528 11200 38534 11212
rect 38838 11200 38844 11212
rect 38528 11172 38844 11200
rect 38528 11160 38534 11172
rect 38838 11160 38844 11172
rect 38896 11160 38902 11212
rect 39132 11209 39160 11240
rect 41690 11228 41696 11280
rect 41748 11268 41754 11280
rect 41748 11240 41793 11268
rect 41748 11228 41754 11240
rect 41874 11228 41880 11280
rect 41932 11268 41938 11280
rect 44013 11268 44041 11308
rect 44726 11296 44732 11308
rect 44784 11296 44790 11348
rect 45005 11339 45063 11345
rect 45005 11305 45017 11339
rect 45051 11336 45063 11339
rect 45094 11336 45100 11348
rect 45051 11308 45100 11336
rect 45051 11305 45063 11308
rect 45005 11299 45063 11305
rect 45094 11296 45100 11308
rect 45152 11296 45158 11348
rect 45649 11339 45707 11345
rect 45649 11305 45661 11339
rect 45695 11336 45707 11339
rect 45695 11308 46336 11336
rect 45695 11305 45707 11308
rect 45649 11299 45707 11305
rect 41932 11240 44041 11268
rect 41932 11228 41938 11240
rect 44082 11228 44088 11280
rect 44140 11268 44146 11280
rect 46106 11268 46112 11280
rect 44140 11240 46112 11268
rect 44140 11228 44146 11240
rect 46106 11228 46112 11240
rect 46164 11228 46170 11280
rect 46308 11268 46336 11308
rect 46382 11296 46388 11348
rect 46440 11336 46446 11348
rect 51166 11336 51172 11348
rect 46440 11308 51172 11336
rect 46440 11296 46446 11308
rect 51166 11296 51172 11308
rect 51224 11296 51230 11348
rect 51350 11296 51356 11348
rect 51408 11336 51414 11348
rect 53469 11339 53527 11345
rect 53469 11336 53481 11339
rect 51408 11308 53481 11336
rect 51408 11296 51414 11308
rect 53469 11305 53481 11308
rect 53515 11305 53527 11339
rect 53469 11299 53527 11305
rect 55122 11296 55128 11348
rect 55180 11336 55186 11348
rect 55401 11339 55459 11345
rect 55401 11336 55413 11339
rect 55180 11308 55413 11336
rect 55180 11296 55186 11308
rect 55401 11305 55413 11308
rect 55447 11305 55459 11339
rect 55401 11299 55459 11305
rect 55582 11296 55588 11348
rect 55640 11336 55646 11348
rect 55953 11339 56011 11345
rect 55953 11336 55965 11339
rect 55640 11308 55965 11336
rect 55640 11296 55646 11308
rect 55953 11305 55965 11308
rect 55999 11305 56011 11339
rect 59725 11339 59783 11345
rect 55953 11299 56011 11305
rect 56060 11308 59308 11336
rect 47578 11268 47584 11280
rect 46308 11240 47440 11268
rect 47539 11240 47584 11268
rect 39117 11203 39175 11209
rect 39117 11169 39129 11203
rect 39163 11169 39175 11203
rect 39117 11163 39175 11169
rect 41049 11203 41107 11209
rect 41049 11169 41061 11203
rect 41095 11200 41107 11203
rect 41138 11200 41144 11212
rect 41095 11172 41144 11200
rect 41095 11169 41107 11172
rect 41049 11163 41107 11169
rect 41138 11160 41144 11172
rect 41196 11160 41202 11212
rect 41322 11200 41328 11212
rect 41283 11172 41328 11200
rect 41322 11160 41328 11172
rect 41380 11160 41386 11212
rect 42242 11160 42248 11212
rect 42300 11200 42306 11212
rect 43070 11200 43076 11212
rect 42300 11172 43076 11200
rect 42300 11160 42306 11172
rect 43070 11160 43076 11172
rect 43128 11200 43134 11212
rect 47412 11200 47440 11240
rect 47578 11228 47584 11240
rect 47636 11228 47642 11280
rect 49421 11271 49479 11277
rect 49421 11237 49433 11271
rect 49467 11237 49479 11271
rect 49421 11231 49479 11237
rect 49234 11200 49240 11212
rect 43128 11172 47348 11200
rect 47412 11172 49240 11200
rect 43128 11160 43134 11172
rect 46109 11169 46167 11172
rect 35805 11135 35863 11141
rect 35805 11101 35817 11135
rect 35851 11101 35863 11135
rect 35986 11132 35992 11144
rect 35947 11104 35992 11132
rect 35805 11095 35863 11101
rect 35986 11092 35992 11104
rect 36044 11092 36050 11144
rect 36078 11092 36084 11144
rect 36136 11132 36142 11144
rect 36136 11104 36181 11132
rect 36136 11092 36142 11104
rect 36446 11092 36452 11144
rect 36504 11132 36510 11144
rect 36909 11135 36967 11141
rect 36909 11132 36921 11135
rect 36504 11104 36921 11132
rect 36504 11092 36510 11104
rect 36909 11101 36921 11104
rect 36955 11132 36967 11135
rect 37090 11132 37096 11144
rect 36955 11104 37096 11132
rect 36955 11101 36967 11104
rect 36909 11095 36967 11101
rect 37090 11092 37096 11104
rect 37148 11132 37154 11144
rect 37987 11135 38045 11141
rect 37148 11128 37872 11132
rect 37987 11128 37999 11135
rect 37148 11104 37999 11128
rect 37148 11092 37154 11104
rect 37844 11101 37999 11104
rect 38033 11101 38045 11135
rect 37844 11100 38045 11101
rect 37987 11095 38045 11100
rect 38102 11092 38108 11144
rect 38160 11132 38166 11144
rect 38160 11104 38205 11132
rect 38160 11092 38166 11104
rect 38286 11092 38292 11144
rect 38344 11132 38350 11144
rect 38930 11132 38936 11144
rect 38344 11104 38389 11132
rect 38891 11104 38936 11132
rect 38344 11092 38350 11104
rect 38930 11092 38936 11104
rect 38988 11092 38994 11144
rect 39022 11092 39028 11144
rect 39080 11132 39086 11144
rect 39080 11104 39125 11132
rect 39080 11092 39086 11104
rect 39206 11092 39212 11144
rect 39264 11132 39270 11144
rect 40034 11132 40040 11144
rect 39264 11104 39309 11132
rect 39995 11104 40040 11132
rect 39264 11092 39270 11104
rect 40034 11092 40040 11104
rect 40092 11092 40098 11144
rect 40218 11092 40224 11144
rect 40276 11132 40282 11144
rect 40313 11135 40371 11141
rect 40313 11132 40325 11135
rect 40276 11104 40325 11132
rect 40276 11092 40282 11104
rect 40313 11101 40325 11104
rect 40359 11101 40371 11135
rect 40313 11095 40371 11101
rect 40862 11092 40868 11144
rect 40920 11132 40926 11144
rect 40957 11135 41015 11141
rect 40957 11132 40969 11135
rect 40920 11104 40969 11132
rect 40920 11092 40926 11104
rect 40957 11101 40969 11104
rect 41003 11101 41015 11135
rect 40957 11095 41015 11101
rect 41693 11135 41751 11141
rect 41693 11101 41705 11135
rect 41739 11132 41751 11135
rect 41782 11132 41788 11144
rect 41739 11104 41788 11132
rect 41739 11101 41751 11104
rect 41693 11095 41751 11101
rect 41782 11092 41788 11104
rect 41840 11092 41846 11144
rect 41966 11092 41972 11144
rect 42024 11132 42030 11144
rect 42024 11104 42069 11132
rect 42024 11092 42030 11104
rect 42334 11092 42340 11144
rect 42392 11132 42398 11144
rect 42521 11135 42579 11141
rect 42521 11132 42533 11135
rect 42392 11104 42533 11132
rect 42392 11092 42398 11104
rect 42521 11101 42533 11104
rect 42567 11101 42579 11135
rect 44266 11132 44272 11144
rect 44227 11104 44272 11132
rect 42521 11095 42579 11101
rect 44266 11092 44272 11104
rect 44324 11092 44330 11144
rect 44358 11092 44364 11144
rect 44416 11132 44422 11144
rect 44545 11135 44603 11141
rect 44416 11104 44461 11132
rect 44416 11092 44422 11104
rect 44545 11101 44557 11135
rect 44591 11132 44603 11135
rect 45189 11135 45247 11141
rect 45189 11132 45201 11135
rect 44591 11104 45201 11132
rect 44591 11101 44603 11104
rect 44545 11095 44603 11101
rect 45189 11101 45201 11104
rect 45235 11101 45247 11135
rect 45189 11095 45247 11101
rect 45554 11092 45560 11144
rect 45612 11132 45618 11144
rect 45833 11135 45891 11141
rect 45833 11132 45845 11135
rect 45612 11104 45845 11132
rect 45612 11092 45618 11104
rect 45833 11101 45845 11104
rect 45879 11101 45891 11135
rect 46014 11132 46020 11144
rect 45975 11104 46020 11132
rect 45833 11095 45891 11101
rect 46014 11092 46020 11104
rect 46072 11092 46078 11144
rect 46109 11135 46121 11169
rect 46155 11135 46167 11169
rect 46109 11129 46167 11135
rect 46198 11092 46204 11144
rect 46256 11132 46262 11144
rect 46658 11132 46664 11144
rect 46256 11104 46664 11132
rect 46256 11092 46262 11104
rect 46658 11092 46664 11104
rect 46716 11092 46722 11144
rect 46750 11092 46756 11144
rect 46808 11132 46814 11144
rect 46845 11135 46903 11141
rect 46845 11132 46857 11135
rect 46808 11104 46857 11132
rect 46808 11092 46814 11104
rect 46845 11101 46857 11104
rect 46891 11101 46903 11135
rect 46845 11095 46903 11101
rect 46937 11135 46995 11141
rect 46937 11101 46949 11135
rect 46983 11132 46995 11135
rect 47210 11132 47216 11144
rect 46983 11104 47216 11132
rect 46983 11101 46995 11104
rect 46937 11095 46995 11101
rect 47210 11092 47216 11104
rect 47268 11092 47274 11144
rect 47320 11132 47348 11172
rect 49234 11160 49240 11172
rect 49292 11160 49298 11212
rect 49436 11200 49464 11231
rect 49970 11228 49976 11280
rect 50028 11268 50034 11280
rect 50801 11271 50859 11277
rect 50801 11268 50813 11271
rect 50028 11240 50813 11268
rect 50028 11228 50034 11240
rect 50801 11237 50813 11240
rect 50847 11237 50859 11271
rect 50801 11231 50859 11237
rect 52549 11271 52607 11277
rect 52549 11237 52561 11271
rect 52595 11268 52607 11271
rect 53926 11268 53932 11280
rect 52595 11240 53932 11268
rect 52595 11237 52607 11240
rect 52549 11231 52607 11237
rect 53926 11228 53932 11240
rect 53984 11228 53990 11280
rect 56060 11268 56088 11308
rect 54036 11240 56088 11268
rect 49436 11172 50108 11200
rect 47397 11135 47455 11141
rect 47397 11132 47409 11135
rect 47320 11104 47409 11132
rect 47397 11101 47409 11104
rect 47443 11101 47455 11135
rect 49418 11132 49424 11144
rect 49379 11104 49424 11132
rect 47397 11095 47455 11101
rect 49418 11092 49424 11104
rect 49476 11092 49482 11144
rect 49697 11135 49755 11141
rect 49697 11101 49709 11135
rect 49743 11132 49755 11135
rect 49786 11132 49792 11144
rect 49743 11104 49792 11132
rect 49743 11101 49755 11104
rect 49697 11095 49755 11101
rect 49786 11092 49792 11104
rect 49844 11092 49850 11144
rect 33134 11073 33140 11076
rect 29794 11067 29852 11073
rect 29794 11064 29806 11067
rect 26292 11036 28856 11064
rect 28920 11036 29806 11064
rect 26292 11024 26298 11036
rect 25866 10996 25872 11008
rect 24872 10968 25872 10996
rect 25866 10956 25872 10968
rect 25924 10956 25930 11008
rect 27154 10996 27160 11008
rect 27115 10968 27160 10996
rect 27154 10956 27160 10968
rect 27212 10996 27218 11008
rect 27338 10996 27344 11008
rect 27212 10968 27344 10996
rect 27212 10956 27218 10968
rect 27338 10956 27344 10968
rect 27396 10956 27402 11008
rect 28920 11005 28948 11036
rect 29794 11033 29806 11036
rect 29840 11033 29852 11067
rect 33128 11064 33140 11073
rect 33095 11036 33140 11064
rect 29794 11027 29852 11033
rect 33128 11027 33140 11036
rect 33134 11024 33140 11027
rect 33192 11024 33198 11076
rect 33226 11024 33232 11076
rect 33284 11024 33290 11076
rect 37550 11024 37556 11076
rect 37608 11064 37614 11076
rect 37608 11036 37872 11064
rect 37608 11024 37614 11036
rect 28905 10999 28963 11005
rect 28905 10965 28917 10999
rect 28951 10965 28963 10999
rect 28905 10959 28963 10965
rect 30006 10956 30012 11008
rect 30064 10996 30070 11008
rect 30929 10999 30987 11005
rect 30929 10996 30941 10999
rect 30064 10968 30941 10996
rect 30064 10956 30070 10968
rect 30929 10965 30941 10968
rect 30975 10996 30987 10999
rect 32766 10996 32772 11008
rect 30975 10968 32772 10996
rect 30975 10965 30987 10968
rect 30929 10959 30987 10965
rect 32766 10956 32772 10968
rect 32824 10956 32830 11008
rect 35066 10996 35072 11008
rect 35027 10968 35072 10996
rect 35066 10956 35072 10968
rect 35124 10956 35130 11008
rect 35158 10956 35164 11008
rect 35216 10996 35222 11008
rect 37734 10996 37740 11008
rect 35216 10968 37740 10996
rect 35216 10956 35222 10968
rect 37734 10956 37740 10968
rect 37792 10956 37798 11008
rect 37844 11005 37872 11036
rect 38562 11024 38568 11076
rect 38620 11064 38626 11076
rect 41322 11064 41328 11076
rect 38620 11036 41328 11064
rect 38620 11024 38626 11036
rect 41322 11024 41328 11036
rect 41380 11024 41386 11076
rect 41874 11024 41880 11076
rect 41932 11064 41938 11076
rect 41932 11036 41977 11064
rect 41932 11024 41938 11036
rect 44634 11024 44640 11076
rect 44692 11064 44698 11076
rect 46477 11067 46535 11073
rect 46477 11064 46489 11067
rect 44692 11036 46489 11064
rect 44692 11024 44698 11036
rect 46477 11033 46489 11036
rect 46523 11033 46535 11067
rect 46477 11027 46535 11033
rect 49605 11067 49663 11073
rect 49605 11033 49617 11067
rect 49651 11064 49663 11067
rect 49970 11064 49976 11076
rect 49651 11036 49976 11064
rect 49651 11033 49663 11036
rect 49605 11027 49663 11033
rect 49970 11024 49976 11036
rect 50028 11024 50034 11076
rect 50080 11064 50108 11172
rect 50154 11160 50160 11212
rect 50212 11200 50218 11212
rect 50338 11200 50344 11212
rect 50212 11172 50344 11200
rect 50212 11160 50218 11172
rect 50338 11160 50344 11172
rect 50396 11200 50402 11212
rect 51169 11203 51227 11209
rect 51169 11200 51181 11203
rect 50396 11172 51181 11200
rect 50396 11160 50402 11172
rect 51169 11169 51181 11172
rect 51215 11169 51227 11203
rect 51169 11163 51227 11169
rect 52270 11160 52276 11212
rect 52328 11200 52334 11212
rect 54036 11200 54064 11240
rect 57790 11228 57796 11280
rect 57848 11268 57854 11280
rect 57977 11271 58035 11277
rect 57977 11268 57989 11271
rect 57848 11240 57989 11268
rect 57848 11228 57854 11240
rect 57977 11237 57989 11240
rect 58023 11237 58035 11271
rect 59280 11268 59308 11308
rect 59725 11305 59737 11339
rect 59771 11336 59783 11339
rect 59998 11336 60004 11348
rect 59771 11308 60004 11336
rect 59771 11305 59783 11308
rect 59725 11299 59783 11305
rect 59998 11296 60004 11308
rect 60056 11296 60062 11348
rect 60461 11339 60519 11345
rect 60461 11305 60473 11339
rect 60507 11336 60519 11339
rect 60734 11336 60740 11348
rect 60507 11308 60740 11336
rect 60507 11305 60519 11308
rect 60461 11299 60519 11305
rect 60734 11296 60740 11308
rect 60792 11296 60798 11348
rect 61930 11336 61936 11348
rect 60936 11308 61936 11336
rect 60936 11268 60964 11308
rect 61930 11296 61936 11308
rect 61988 11296 61994 11348
rect 62301 11339 62359 11345
rect 62301 11305 62313 11339
rect 62347 11336 62359 11339
rect 62574 11336 62580 11348
rect 62347 11308 62580 11336
rect 62347 11305 62359 11308
rect 62301 11299 62359 11305
rect 62574 11296 62580 11308
rect 62632 11296 62638 11348
rect 62666 11296 62672 11348
rect 62724 11336 62730 11348
rect 67726 11336 67732 11348
rect 62724 11308 67732 11336
rect 62724 11296 62730 11308
rect 67726 11296 67732 11308
rect 67784 11296 67790 11348
rect 69290 11296 69296 11348
rect 69348 11336 69354 11348
rect 73798 11336 73804 11348
rect 69348 11308 73804 11336
rect 69348 11296 69354 11308
rect 73798 11296 73804 11308
rect 73856 11296 73862 11348
rect 59280 11240 60964 11268
rect 61013 11271 61071 11277
rect 57977 11231 58035 11237
rect 61013 11237 61025 11271
rect 61059 11268 61071 11271
rect 62206 11268 62212 11280
rect 61059 11240 62212 11268
rect 61059 11237 61071 11240
rect 61013 11231 61071 11237
rect 62206 11228 62212 11240
rect 62264 11228 62270 11280
rect 67269 11271 67327 11277
rect 62960 11240 65288 11268
rect 52328 11172 54064 11200
rect 52328 11160 52334 11172
rect 55490 11160 55496 11212
rect 55548 11200 55554 11212
rect 56597 11203 56655 11209
rect 56597 11200 56609 11203
rect 55548 11172 56609 11200
rect 55548 11160 55554 11172
rect 56597 11169 56609 11172
rect 56643 11169 56655 11203
rect 60550 11200 60556 11212
rect 56597 11163 56655 11169
rect 59556 11172 60556 11200
rect 50522 11132 50528 11144
rect 50483 11104 50528 11132
rect 50522 11092 50528 11104
rect 50580 11092 50586 11144
rect 50614 11092 50620 11144
rect 50672 11132 50678 11144
rect 52917 11135 52975 11141
rect 52917 11132 52929 11135
rect 50672 11104 50717 11132
rect 51046 11104 52929 11132
rect 50672 11092 50678 11104
rect 51046 11064 51074 11104
rect 52917 11101 52929 11104
rect 52963 11101 52975 11135
rect 53098 11132 53104 11144
rect 53059 11104 53104 11132
rect 52917 11095 52975 11101
rect 53098 11092 53104 11104
rect 53156 11092 53162 11144
rect 53285 11135 53343 11141
rect 53285 11101 53297 11135
rect 53331 11132 53343 11135
rect 55214 11132 55220 11144
rect 53331 11104 55220 11132
rect 53331 11101 53343 11104
rect 53285 11095 53343 11101
rect 55214 11092 55220 11104
rect 55272 11092 55278 11144
rect 55309 11135 55367 11141
rect 55309 11101 55321 11135
rect 55355 11132 55367 11135
rect 56042 11132 56048 11144
rect 55355 11104 56048 11132
rect 55355 11101 55367 11104
rect 55309 11095 55367 11101
rect 56042 11092 56048 11104
rect 56100 11092 56106 11144
rect 56137 11135 56195 11141
rect 56137 11101 56149 11135
rect 56183 11132 56195 11135
rect 56226 11132 56232 11144
rect 56183 11104 56232 11132
rect 56183 11101 56195 11104
rect 56137 11095 56195 11101
rect 56226 11092 56232 11104
rect 56284 11092 56290 11144
rect 58345 11135 58403 11141
rect 58345 11101 58357 11135
rect 58391 11132 58403 11135
rect 58434 11132 58440 11144
rect 58391 11104 58440 11132
rect 58391 11101 58403 11104
rect 58345 11095 58403 11101
rect 58434 11092 58440 11104
rect 58492 11132 58498 11144
rect 59446 11132 59452 11144
rect 58492 11104 59452 11132
rect 58492 11092 58498 11104
rect 59446 11092 59452 11104
rect 59504 11092 59510 11144
rect 50080 11036 51074 11064
rect 51436 11067 51494 11073
rect 51436 11033 51448 11067
rect 51482 11064 51494 11067
rect 52730 11064 52736 11076
rect 51482 11036 52736 11064
rect 51482 11033 51494 11036
rect 51436 11027 51494 11033
rect 52730 11024 52736 11036
rect 52788 11024 52794 11076
rect 52822 11024 52828 11076
rect 52880 11064 52886 11076
rect 53193 11067 53251 11073
rect 53193 11064 53205 11067
rect 52880 11036 53205 11064
rect 52880 11024 52886 11036
rect 53193 11033 53205 11036
rect 53239 11064 53251 11067
rect 54570 11064 54576 11076
rect 53239 11036 54576 11064
rect 53239 11033 53251 11036
rect 53193 11027 53251 11033
rect 54570 11024 54576 11036
rect 54628 11024 54634 11076
rect 54754 11024 54760 11076
rect 54812 11064 54818 11076
rect 56686 11064 56692 11076
rect 54812 11036 56692 11064
rect 54812 11024 54818 11036
rect 56686 11024 56692 11036
rect 56744 11024 56750 11076
rect 56864 11067 56922 11073
rect 56864 11033 56876 11067
rect 56910 11064 56922 11067
rect 57054 11064 57060 11076
rect 56910 11036 57060 11064
rect 56910 11033 56922 11036
rect 56864 11027 56922 11033
rect 57054 11024 57060 11036
rect 57112 11024 57118 11076
rect 58066 11024 58072 11076
rect 58124 11064 58130 11076
rect 58590 11067 58648 11073
rect 58590 11064 58602 11067
rect 58124 11036 58602 11064
rect 58124 11024 58130 11036
rect 58590 11033 58602 11036
rect 58636 11033 58648 11067
rect 58590 11027 58648 11033
rect 58894 11024 58900 11076
rect 58952 11064 58958 11076
rect 59556 11064 59584 11172
rect 60550 11160 60556 11172
rect 60608 11160 60614 11212
rect 61565 11203 61623 11209
rect 61565 11200 61577 11203
rect 61120 11172 61577 11200
rect 60642 11132 60648 11144
rect 60603 11104 60648 11132
rect 60642 11092 60648 11104
rect 60700 11092 60706 11144
rect 58952 11036 59584 11064
rect 58952 11024 58958 11036
rect 59630 11024 59636 11076
rect 59688 11064 59694 11076
rect 61120 11064 61148 11172
rect 61565 11169 61577 11172
rect 61611 11169 61623 11203
rect 62960 11200 62988 11240
rect 61565 11163 61623 11169
rect 62132 11172 62988 11200
rect 61378 11132 61384 11144
rect 61339 11104 61384 11132
rect 61378 11092 61384 11104
rect 61436 11092 61442 11144
rect 61473 11135 61531 11141
rect 61473 11101 61485 11135
rect 61519 11132 61531 11135
rect 62132 11132 62160 11172
rect 63034 11160 63040 11212
rect 63092 11200 63098 11212
rect 63589 11203 63647 11209
rect 63589 11200 63601 11203
rect 63092 11172 63601 11200
rect 63092 11160 63098 11172
rect 63589 11169 63601 11172
rect 63635 11169 63647 11203
rect 63589 11163 63647 11169
rect 63773 11203 63831 11209
rect 63773 11169 63785 11203
rect 63819 11200 63831 11203
rect 65150 11200 65156 11212
rect 63819 11172 65156 11200
rect 63819 11169 63831 11172
rect 63773 11163 63831 11169
rect 65150 11160 65156 11172
rect 65208 11160 65214 11212
rect 62301 11135 62359 11141
rect 62301 11132 62313 11135
rect 61519 11104 62160 11132
rect 62224 11104 62313 11132
rect 61519 11101 61531 11104
rect 61473 11095 61531 11101
rect 59688 11036 61148 11064
rect 59688 11024 59694 11036
rect 61194 11024 61200 11076
rect 61252 11064 61258 11076
rect 62224 11064 62252 11104
rect 62301 11101 62313 11104
rect 62347 11132 62359 11135
rect 62482 11132 62488 11144
rect 62347 11104 62488 11132
rect 62347 11101 62359 11104
rect 62301 11095 62359 11101
rect 62482 11092 62488 11104
rect 62540 11092 62546 11144
rect 62577 11135 62635 11141
rect 62577 11101 62589 11135
rect 62623 11101 62635 11135
rect 62577 11095 62635 11101
rect 62592 11064 62620 11095
rect 62850 11092 62856 11144
rect 62908 11132 62914 11144
rect 63865 11135 63923 11141
rect 62908 11104 63540 11132
rect 62908 11092 62914 11104
rect 61252 11036 62252 11064
rect 62316 11036 62620 11064
rect 61252 11024 61258 11036
rect 37829 10999 37887 11005
rect 37829 10965 37841 10999
rect 37875 10965 37887 10999
rect 37829 10959 37887 10965
rect 40126 10956 40132 11008
rect 40184 10996 40190 11008
rect 40221 10999 40279 11005
rect 40221 10996 40233 10999
rect 40184 10968 40233 10996
rect 40184 10956 40190 10968
rect 40221 10965 40233 10968
rect 40267 10965 40279 10999
rect 40221 10959 40279 10965
rect 40310 10956 40316 11008
rect 40368 10996 40374 11008
rect 41046 10996 41052 11008
rect 40368 10968 41052 10996
rect 40368 10956 40374 10968
rect 41046 10956 41052 10968
rect 41104 10956 41110 11008
rect 41138 10956 41144 11008
rect 41196 10996 41202 11008
rect 61838 10996 61844 11008
rect 41196 10968 61844 10996
rect 41196 10956 41202 10968
rect 61838 10956 61844 10968
rect 61896 10956 61902 11008
rect 61930 10956 61936 11008
rect 61988 10996 61994 11008
rect 62316 10996 62344 11036
rect 63310 11024 63316 11076
rect 63368 11064 63374 11076
rect 63405 11067 63463 11073
rect 63405 11064 63417 11067
rect 63368 11036 63417 11064
rect 63368 11024 63374 11036
rect 63405 11033 63417 11036
rect 63451 11033 63463 11067
rect 63512 11064 63540 11104
rect 63865 11101 63877 11135
rect 63911 11132 63923 11135
rect 64046 11132 64052 11144
rect 63911 11104 64052 11132
rect 63911 11101 63923 11104
rect 63865 11095 63923 11101
rect 64046 11092 64052 11104
rect 64104 11092 64110 11144
rect 64230 11132 64236 11144
rect 64191 11104 64236 11132
rect 64230 11092 64236 11104
rect 64288 11092 64294 11144
rect 64322 11092 64328 11144
rect 64380 11132 64386 11144
rect 64417 11135 64475 11141
rect 64417 11132 64429 11135
rect 64380 11104 64429 11132
rect 64380 11092 64386 11104
rect 64417 11101 64429 11104
rect 64463 11101 64475 11135
rect 64417 11095 64475 11101
rect 64506 11092 64512 11144
rect 64564 11132 64570 11144
rect 64693 11135 64751 11141
rect 64693 11132 64705 11135
rect 64564 11104 64705 11132
rect 64564 11092 64570 11104
rect 64693 11101 64705 11104
rect 64739 11101 64751 11135
rect 64693 11095 64751 11101
rect 65260 11064 65288 11240
rect 67269 11237 67281 11271
rect 67315 11268 67327 11271
rect 67450 11268 67456 11280
rect 67315 11240 67456 11268
rect 67315 11237 67327 11240
rect 67269 11231 67327 11237
rect 67450 11228 67456 11240
rect 67508 11228 67514 11280
rect 67542 11228 67548 11280
rect 67600 11228 67606 11280
rect 69106 11228 69112 11280
rect 69164 11268 69170 11280
rect 69201 11271 69259 11277
rect 69201 11268 69213 11271
rect 69164 11240 69213 11268
rect 69164 11228 69170 11240
rect 69201 11237 69213 11240
rect 69247 11237 69259 11271
rect 69201 11231 69259 11237
rect 69382 11228 69388 11280
rect 69440 11268 69446 11280
rect 73982 11268 73988 11280
rect 69440 11240 73988 11268
rect 69440 11228 69446 11240
rect 73982 11228 73988 11240
rect 74040 11228 74046 11280
rect 75886 11240 87736 11268
rect 67082 11160 67088 11212
rect 67140 11200 67146 11212
rect 67560 11200 67588 11228
rect 67818 11200 67824 11212
rect 67140 11172 67404 11200
rect 67560 11172 67824 11200
rect 67140 11160 67146 11172
rect 67266 11132 67272 11144
rect 67227 11104 67272 11132
rect 67266 11092 67272 11104
rect 67324 11092 67330 11144
rect 67376 11126 67404 11172
rect 67818 11160 67824 11172
rect 67876 11160 67882 11212
rect 67453 11135 67511 11141
rect 67453 11126 67465 11135
rect 67376 11101 67465 11126
rect 67499 11101 67511 11135
rect 75886 11132 75914 11240
rect 87506 11200 87512 11212
rect 67376 11098 67511 11101
rect 67453 11095 67511 11098
rect 67560 11104 75914 11132
rect 80026 11172 87512 11200
rect 67560 11064 67588 11104
rect 63512 11036 63908 11064
rect 65260 11036 67588 11064
rect 63405 11027 63463 11033
rect 61988 10968 62344 10996
rect 62485 10999 62543 11005
rect 61988 10956 61994 10968
rect 62485 10965 62497 10999
rect 62531 10996 62543 10999
rect 62758 10996 62764 11008
rect 62531 10968 62764 10996
rect 62531 10965 62543 10968
rect 62485 10959 62543 10965
rect 62758 10956 62764 10968
rect 62816 10956 62822 11008
rect 63880 10996 63908 11036
rect 67634 11024 67640 11076
rect 67692 11064 67698 11076
rect 68066 11067 68124 11073
rect 68066 11064 68078 11067
rect 67692 11036 68078 11064
rect 67692 11024 67698 11036
rect 68066 11033 68078 11036
rect 68112 11033 68124 11067
rect 68066 11027 68124 11033
rect 69106 11024 69112 11076
rect 69164 11064 69170 11076
rect 80026 11064 80054 11172
rect 87506 11160 87512 11172
rect 87564 11160 87570 11212
rect 87708 11209 87736 11240
rect 87693 11203 87751 11209
rect 87693 11169 87705 11203
rect 87739 11169 87751 11203
rect 87693 11163 87751 11169
rect 87414 11132 87420 11144
rect 87375 11104 87420 11132
rect 87414 11092 87420 11104
rect 87472 11092 87478 11144
rect 69164 11036 80054 11064
rect 69164 11024 69170 11036
rect 64601 10999 64659 11005
rect 64601 10996 64613 10999
rect 63880 10968 64613 10996
rect 64601 10965 64613 10968
rect 64647 10965 64659 10999
rect 64601 10959 64659 10965
rect 67450 10956 67456 11008
rect 67508 10996 67514 11008
rect 87690 10996 87696 11008
rect 67508 10968 87696 10996
rect 67508 10956 67514 10968
rect 87690 10956 87696 10968
rect 87748 10956 87754 11008
rect 1104 10906 88872 10928
rect 1104 10854 22898 10906
rect 22950 10854 22962 10906
rect 23014 10854 23026 10906
rect 23078 10854 23090 10906
rect 23142 10854 23154 10906
rect 23206 10854 44846 10906
rect 44898 10854 44910 10906
rect 44962 10854 44974 10906
rect 45026 10854 45038 10906
rect 45090 10854 45102 10906
rect 45154 10854 66794 10906
rect 66846 10854 66858 10906
rect 66910 10854 66922 10906
rect 66974 10854 66986 10906
rect 67038 10854 67050 10906
rect 67102 10854 88872 10906
rect 1104 10832 88872 10854
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 24765 10795 24823 10801
rect 24765 10792 24777 10795
rect 20956 10764 24777 10792
rect 20956 10752 20962 10764
rect 24765 10761 24777 10764
rect 24811 10792 24823 10795
rect 26142 10792 26148 10804
rect 24811 10764 26004 10792
rect 26103 10764 26148 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 25976 10724 26004 10764
rect 26142 10752 26148 10764
rect 26200 10752 26206 10804
rect 29089 10795 29147 10801
rect 29089 10761 29101 10795
rect 29135 10792 29147 10795
rect 29730 10792 29736 10804
rect 29135 10764 29736 10792
rect 29135 10761 29147 10764
rect 29089 10755 29147 10761
rect 29730 10752 29736 10764
rect 29788 10752 29794 10804
rect 30742 10752 30748 10804
rect 30800 10792 30806 10804
rect 31478 10792 31484 10804
rect 30800 10764 31484 10792
rect 30800 10752 30806 10764
rect 31478 10752 31484 10764
rect 31536 10752 31542 10804
rect 33045 10795 33103 10801
rect 33045 10761 33057 10795
rect 33091 10792 33103 10795
rect 33134 10792 33140 10804
rect 33091 10764 33140 10792
rect 33091 10761 33103 10764
rect 33045 10755 33103 10761
rect 33134 10752 33140 10764
rect 33192 10752 33198 10804
rect 33594 10752 33600 10804
rect 33652 10792 33658 10804
rect 33689 10795 33747 10801
rect 33689 10792 33701 10795
rect 33652 10764 33701 10792
rect 33652 10752 33658 10764
rect 33689 10761 33701 10764
rect 33735 10761 33747 10795
rect 33689 10755 33747 10761
rect 33870 10752 33876 10804
rect 33928 10792 33934 10804
rect 35158 10792 35164 10804
rect 33928 10764 35164 10792
rect 33928 10752 33934 10764
rect 35158 10752 35164 10764
rect 35216 10752 35222 10804
rect 35805 10795 35863 10801
rect 35805 10761 35817 10795
rect 35851 10792 35863 10795
rect 36998 10792 37004 10804
rect 35851 10764 37004 10792
rect 35851 10761 35863 10764
rect 35805 10755 35863 10761
rect 36998 10752 37004 10764
rect 37056 10752 37062 10804
rect 37550 10752 37556 10804
rect 37608 10792 37614 10804
rect 38470 10792 38476 10804
rect 37608 10764 38476 10792
rect 37608 10752 37614 10764
rect 38470 10752 38476 10764
rect 38528 10752 38534 10804
rect 39025 10795 39083 10801
rect 39025 10761 39037 10795
rect 39071 10792 39083 10795
rect 40218 10792 40224 10804
rect 39071 10764 40224 10792
rect 39071 10761 39083 10764
rect 39025 10755 39083 10761
rect 40218 10752 40224 10764
rect 40276 10752 40282 10804
rect 40865 10795 40923 10801
rect 40865 10761 40877 10795
rect 40911 10792 40923 10795
rect 87690 10792 87696 10804
rect 40911 10764 66668 10792
rect 40911 10761 40923 10764
rect 40865 10755 40923 10761
rect 27154 10724 27160 10736
rect 25976 10696 27160 10724
rect 27154 10684 27160 10696
rect 27212 10684 27218 10736
rect 29822 10724 29828 10736
rect 29196 10696 29828 10724
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 27062 10656 27068 10668
rect 25056 10628 27068 10656
rect 23382 10548 23388 10600
rect 23440 10588 23446 10600
rect 25056 10597 25084 10628
rect 27062 10616 27068 10628
rect 27120 10616 27126 10668
rect 28261 10659 28319 10665
rect 28261 10625 28273 10659
rect 28307 10656 28319 10659
rect 28994 10656 29000 10668
rect 28307 10628 28672 10656
rect 28955 10628 29000 10656
rect 28307 10625 28319 10628
rect 28261 10619 28319 10625
rect 24857 10591 24915 10597
rect 24857 10588 24869 10591
rect 23440 10560 24869 10588
rect 23440 10548 23446 10560
rect 24857 10557 24869 10560
rect 24903 10557 24915 10591
rect 24857 10551 24915 10557
rect 25041 10591 25099 10597
rect 25041 10557 25053 10591
rect 25087 10557 25099 10591
rect 25041 10551 25099 10557
rect 25685 10591 25743 10597
rect 25685 10557 25697 10591
rect 25731 10588 25743 10591
rect 25866 10588 25872 10600
rect 25731 10560 25872 10588
rect 25731 10557 25743 10560
rect 25685 10551 25743 10557
rect 25866 10548 25872 10560
rect 25924 10548 25930 10600
rect 24486 10480 24492 10532
rect 24544 10520 24550 10532
rect 25961 10523 26019 10529
rect 25961 10520 25973 10523
rect 24544 10492 25973 10520
rect 24544 10480 24550 10492
rect 25961 10489 25973 10492
rect 26007 10520 26019 10523
rect 26418 10520 26424 10532
rect 26007 10492 26424 10520
rect 26007 10489 26019 10492
rect 25961 10483 26019 10489
rect 26418 10480 26424 10492
rect 26476 10480 26482 10532
rect 28644 10529 28672 10628
rect 28994 10616 29000 10628
rect 29052 10616 29058 10668
rect 29196 10597 29224 10696
rect 29822 10684 29828 10696
rect 29880 10724 29886 10736
rect 30282 10724 30288 10736
rect 29880 10696 30288 10724
rect 29880 10684 29886 10696
rect 30282 10684 30288 10696
rect 30340 10684 30346 10736
rect 32490 10684 32496 10736
rect 32548 10724 32554 10736
rect 33778 10724 33784 10736
rect 32548 10696 33784 10724
rect 32548 10684 32554 10696
rect 33778 10684 33784 10696
rect 33836 10684 33842 10736
rect 35066 10724 35072 10736
rect 33888 10696 35072 10724
rect 29270 10616 29276 10668
rect 29328 10656 29334 10668
rect 29989 10659 30047 10665
rect 29989 10656 30001 10659
rect 29328 10628 30001 10656
rect 29328 10616 29334 10628
rect 29989 10625 30001 10628
rect 30035 10625 30047 10659
rect 29989 10619 30047 10625
rect 33229 10659 33287 10665
rect 33229 10625 33241 10659
rect 33275 10656 33287 10659
rect 33502 10656 33508 10668
rect 33275 10628 33508 10656
rect 33275 10625 33287 10628
rect 33229 10619 33287 10625
rect 33502 10616 33508 10628
rect 33560 10616 33566 10668
rect 33888 10665 33916 10696
rect 35066 10684 35072 10696
rect 35124 10684 35130 10736
rect 38194 10724 38200 10736
rect 36648 10696 38200 10724
rect 33873 10659 33931 10665
rect 33873 10625 33885 10659
rect 33919 10625 33931 10659
rect 34238 10656 34244 10668
rect 34199 10628 34244 10656
rect 33873 10619 33931 10625
rect 34238 10616 34244 10628
rect 34296 10616 34302 10668
rect 35713 10659 35771 10665
rect 35713 10625 35725 10659
rect 35759 10656 35771 10659
rect 36262 10656 36268 10668
rect 35759 10628 36268 10656
rect 35759 10625 35771 10628
rect 35713 10619 35771 10625
rect 36262 10616 36268 10628
rect 36320 10616 36326 10668
rect 36446 10656 36452 10668
rect 36407 10628 36452 10656
rect 36446 10616 36452 10628
rect 36504 10616 36510 10668
rect 36648 10665 36676 10696
rect 38194 10684 38200 10696
rect 38252 10684 38258 10736
rect 39114 10684 39120 10736
rect 39172 10724 39178 10736
rect 50433 10727 50491 10733
rect 50433 10724 50445 10727
rect 39172 10696 50445 10724
rect 39172 10684 39178 10696
rect 50433 10693 50445 10696
rect 50479 10724 50491 10727
rect 51350 10724 51356 10736
rect 50479 10696 51356 10724
rect 50479 10693 50491 10696
rect 50433 10687 50491 10693
rect 51350 10684 51356 10696
rect 51408 10684 51414 10736
rect 51905 10727 51963 10733
rect 51905 10693 51917 10727
rect 51951 10724 51963 10727
rect 54294 10724 54300 10736
rect 51951 10696 54300 10724
rect 51951 10693 51963 10696
rect 51905 10687 51963 10693
rect 54294 10684 54300 10696
rect 54352 10684 54358 10736
rect 56229 10727 56287 10733
rect 56229 10693 56241 10727
rect 56275 10724 56287 10727
rect 56318 10724 56324 10736
rect 56275 10696 56324 10724
rect 56275 10693 56287 10696
rect 56229 10687 56287 10693
rect 56318 10684 56324 10696
rect 56376 10684 56382 10736
rect 56502 10684 56508 10736
rect 56560 10724 56566 10736
rect 56781 10727 56839 10733
rect 56781 10724 56793 10727
rect 56560 10696 56793 10724
rect 56560 10684 56566 10696
rect 56781 10693 56793 10696
rect 56827 10693 56839 10727
rect 56781 10687 56839 10693
rect 58526 10684 58532 10736
rect 58584 10724 58590 10736
rect 58805 10727 58863 10733
rect 58805 10724 58817 10727
rect 58584 10696 58817 10724
rect 58584 10684 58590 10696
rect 58805 10693 58817 10696
rect 58851 10724 58863 10727
rect 59814 10724 59820 10736
rect 58851 10696 59676 10724
rect 59775 10696 59820 10724
rect 58851 10693 58863 10696
rect 58805 10687 58863 10693
rect 36633 10659 36691 10665
rect 36633 10625 36645 10659
rect 36679 10625 36691 10659
rect 37366 10656 37372 10668
rect 36633 10619 36691 10625
rect 37016 10628 37372 10656
rect 29181 10591 29239 10597
rect 29181 10557 29193 10591
rect 29227 10557 29239 10591
rect 29181 10551 29239 10557
rect 29546 10548 29552 10600
rect 29604 10588 29610 10600
rect 29733 10591 29791 10597
rect 29733 10588 29745 10591
rect 29604 10560 29745 10588
rect 29604 10548 29610 10560
rect 29733 10557 29745 10560
rect 29779 10557 29791 10591
rect 29733 10551 29791 10557
rect 36541 10591 36599 10597
rect 36541 10557 36553 10591
rect 36587 10557 36599 10591
rect 36541 10551 36599 10557
rect 36725 10591 36783 10597
rect 36725 10557 36737 10591
rect 36771 10588 36783 10591
rect 37016 10588 37044 10628
rect 37366 10616 37372 10628
rect 37424 10616 37430 10668
rect 37642 10616 37648 10668
rect 37700 10656 37706 10668
rect 38562 10656 38568 10668
rect 37700 10628 38568 10656
rect 37700 10616 37706 10628
rect 38562 10616 38568 10628
rect 38620 10616 38626 10668
rect 39390 10656 39396 10668
rect 39132 10628 39396 10656
rect 36771 10560 37044 10588
rect 36771 10557 36783 10560
rect 36725 10551 36783 10557
rect 28629 10523 28687 10529
rect 28629 10489 28641 10523
rect 28675 10489 28687 10523
rect 36556 10520 36584 10551
rect 37090 10548 37096 10600
rect 37148 10588 37154 10600
rect 37277 10591 37335 10597
rect 37277 10588 37289 10591
rect 37148 10560 37289 10588
rect 37148 10548 37154 10560
rect 37277 10557 37289 10560
rect 37323 10557 37335 10591
rect 37550 10588 37556 10600
rect 37511 10560 37556 10588
rect 37277 10551 37335 10557
rect 28629 10483 28687 10489
rect 30668 10492 36584 10520
rect 37292 10520 37320 10551
rect 37550 10548 37556 10560
rect 37608 10548 37614 10600
rect 38378 10588 38384 10600
rect 37660 10560 38384 10588
rect 37660 10520 37688 10560
rect 38378 10548 38384 10560
rect 38436 10548 38442 10600
rect 39132 10597 39160 10628
rect 39390 10616 39396 10628
rect 39448 10616 39454 10668
rect 39482 10616 39488 10668
rect 39540 10656 39546 10668
rect 40037 10659 40095 10665
rect 40037 10656 40049 10659
rect 39540 10628 40049 10656
rect 39540 10616 39546 10628
rect 40037 10625 40049 10628
rect 40083 10625 40095 10659
rect 40310 10656 40316 10668
rect 40271 10628 40316 10656
rect 40037 10619 40095 10625
rect 40310 10616 40316 10628
rect 40368 10616 40374 10668
rect 40770 10656 40776 10668
rect 40731 10628 40776 10656
rect 40770 10616 40776 10628
rect 40828 10616 40834 10668
rect 41414 10616 41420 10668
rect 41472 10656 41478 10668
rect 42981 10659 43039 10665
rect 41472 10628 42840 10656
rect 41472 10616 41478 10628
rect 39117 10591 39175 10597
rect 39117 10557 39129 10591
rect 39163 10557 39175 10591
rect 39298 10588 39304 10600
rect 39259 10560 39304 10588
rect 39117 10551 39175 10557
rect 39298 10548 39304 10560
rect 39356 10548 39362 10600
rect 40221 10591 40279 10597
rect 40221 10557 40233 10591
rect 40267 10588 40279 10591
rect 42610 10588 42616 10600
rect 40267 10560 42616 10588
rect 40267 10557 40279 10560
rect 40221 10551 40279 10557
rect 42610 10548 42616 10560
rect 42668 10548 42674 10600
rect 42705 10591 42763 10597
rect 42705 10557 42717 10591
rect 42751 10557 42763 10591
rect 42812 10588 42840 10628
rect 42981 10625 42993 10659
rect 43027 10656 43039 10659
rect 43070 10656 43076 10668
rect 43027 10628 43076 10656
rect 43027 10625 43039 10628
rect 42981 10619 43039 10625
rect 43070 10616 43076 10628
rect 43128 10616 43134 10668
rect 43349 10659 43407 10665
rect 43349 10625 43361 10659
rect 43395 10625 43407 10659
rect 45005 10659 45063 10665
rect 45005 10656 45017 10659
rect 43349 10619 43407 10625
rect 43824 10628 45017 10656
rect 43364 10588 43392 10619
rect 42812 10560 43392 10588
rect 42705 10551 42763 10557
rect 37292 10492 37688 10520
rect 38304 10492 41000 10520
rect 1394 10452 1400 10464
rect 1355 10424 1400 10452
rect 1394 10412 1400 10424
rect 1452 10412 1458 10464
rect 24397 10455 24455 10461
rect 24397 10421 24409 10455
rect 24443 10452 24455 10455
rect 25222 10452 25228 10464
rect 24443 10424 25228 10452
rect 24443 10421 24455 10424
rect 24397 10415 24455 10421
rect 25222 10412 25228 10424
rect 25280 10412 25286 10464
rect 28074 10452 28080 10464
rect 28035 10424 28080 10452
rect 28074 10412 28080 10424
rect 28132 10412 28138 10464
rect 30098 10412 30104 10464
rect 30156 10452 30162 10464
rect 30668 10452 30696 10492
rect 31110 10452 31116 10464
rect 30156 10424 30696 10452
rect 31071 10424 31116 10452
rect 30156 10412 30162 10424
rect 31110 10412 31116 10424
rect 31168 10412 31174 10464
rect 32306 10412 32312 10464
rect 32364 10452 32370 10464
rect 33870 10452 33876 10464
rect 32364 10424 33876 10452
rect 32364 10412 32370 10424
rect 33870 10412 33876 10424
rect 33928 10412 33934 10464
rect 34330 10452 34336 10464
rect 34291 10424 34336 10452
rect 34330 10412 34336 10424
rect 34388 10412 34394 10464
rect 36265 10455 36323 10461
rect 36265 10421 36277 10455
rect 36311 10452 36323 10455
rect 38304 10452 38332 10492
rect 36311 10424 38332 10452
rect 38657 10455 38715 10461
rect 36311 10421 36323 10424
rect 36265 10415 36323 10421
rect 38657 10421 38669 10455
rect 38703 10452 38715 10455
rect 38746 10452 38752 10464
rect 38703 10424 38752 10452
rect 38703 10421 38715 10424
rect 38657 10415 38715 10421
rect 38746 10412 38752 10424
rect 38804 10412 38810 10464
rect 38930 10412 38936 10464
rect 38988 10452 38994 10464
rect 39758 10452 39764 10464
rect 38988 10424 39764 10452
rect 38988 10412 38994 10424
rect 39758 10412 39764 10424
rect 39816 10452 39822 10464
rect 39853 10455 39911 10461
rect 39853 10452 39865 10455
rect 39816 10424 39865 10452
rect 39816 10412 39822 10424
rect 39853 10421 39865 10424
rect 39899 10421 39911 10455
rect 40972 10452 41000 10492
rect 41046 10480 41052 10532
rect 41104 10520 41110 10532
rect 42720 10520 42748 10551
rect 42886 10520 42892 10532
rect 41104 10492 42748 10520
rect 42847 10492 42892 10520
rect 41104 10480 41110 10492
rect 42886 10480 42892 10492
rect 42944 10480 42950 10532
rect 42978 10480 42984 10532
rect 43036 10520 43042 10532
rect 43824 10520 43852 10628
rect 45005 10625 45017 10628
rect 45051 10656 45063 10659
rect 45278 10656 45284 10668
rect 45051 10628 45284 10656
rect 45051 10625 45063 10628
rect 45005 10619 45063 10625
rect 45278 10616 45284 10628
rect 45336 10616 45342 10668
rect 45997 10659 46055 10665
rect 45997 10656 46009 10659
rect 45388 10628 46009 10656
rect 43990 10588 43996 10600
rect 43903 10560 43996 10588
rect 43990 10548 43996 10560
rect 44048 10588 44054 10600
rect 45097 10591 45155 10597
rect 44048 10560 44772 10588
rect 44048 10548 44054 10560
rect 43036 10492 43852 10520
rect 44361 10523 44419 10529
rect 43036 10480 43042 10492
rect 44361 10489 44373 10523
rect 44407 10520 44419 10523
rect 44634 10520 44640 10532
rect 44407 10492 44640 10520
rect 44407 10489 44419 10492
rect 44361 10483 44419 10489
rect 44634 10480 44640 10492
rect 44692 10480 44698 10532
rect 44744 10520 44772 10560
rect 45097 10557 45109 10591
rect 45143 10588 45155 10591
rect 45186 10588 45192 10600
rect 45143 10560 45192 10588
rect 45143 10557 45155 10560
rect 45097 10551 45155 10557
rect 45186 10548 45192 10560
rect 45244 10548 45250 10600
rect 45388 10597 45416 10628
rect 45997 10625 46009 10628
rect 46043 10625 46055 10659
rect 45997 10619 46055 10625
rect 46290 10616 46296 10668
rect 46348 10656 46354 10668
rect 46348 10628 46796 10656
rect 46348 10616 46354 10628
rect 45373 10591 45431 10597
rect 45373 10557 45385 10591
rect 45419 10557 45431 10591
rect 45738 10588 45744 10600
rect 45699 10560 45744 10588
rect 45373 10551 45431 10557
rect 45738 10548 45744 10560
rect 45796 10548 45802 10600
rect 46768 10588 46796 10628
rect 47118 10616 47124 10668
rect 47176 10656 47182 10668
rect 47765 10659 47823 10665
rect 47765 10656 47777 10659
rect 47176 10628 47777 10656
rect 47176 10616 47182 10628
rect 47765 10625 47777 10628
rect 47811 10625 47823 10659
rect 48682 10656 48688 10668
rect 48643 10628 48688 10656
rect 47765 10619 47823 10625
rect 48682 10616 48688 10628
rect 48740 10616 48746 10668
rect 50522 10616 50528 10668
rect 50580 10656 50586 10668
rect 50801 10659 50859 10665
rect 50801 10656 50813 10659
rect 50580 10628 50813 10656
rect 50580 10616 50586 10628
rect 50801 10625 50813 10628
rect 50847 10625 50859 10659
rect 50801 10619 50859 10625
rect 50890 10616 50896 10668
rect 50948 10656 50954 10668
rect 50985 10659 51043 10665
rect 50985 10656 50997 10659
rect 50948 10628 50997 10656
rect 50948 10616 50954 10628
rect 50985 10625 50997 10628
rect 51031 10625 51043 10659
rect 50985 10619 51043 10625
rect 51169 10659 51227 10665
rect 51169 10625 51181 10659
rect 51215 10656 51227 10659
rect 52917 10659 52975 10665
rect 52917 10656 52929 10659
rect 51215 10628 52929 10656
rect 51215 10625 51227 10628
rect 51169 10619 51227 10625
rect 52917 10625 52929 10628
rect 52963 10625 52975 10659
rect 52917 10619 52975 10625
rect 53098 10616 53104 10668
rect 53156 10656 53162 10668
rect 53469 10659 53527 10665
rect 53469 10656 53481 10659
rect 53156 10628 53481 10656
rect 53156 10616 53162 10628
rect 53469 10625 53481 10628
rect 53515 10625 53527 10659
rect 53469 10619 53527 10625
rect 54478 10616 54484 10668
rect 54536 10656 54542 10668
rect 54645 10659 54703 10665
rect 54645 10656 54657 10659
rect 54536 10628 54657 10656
rect 54536 10616 54542 10628
rect 54645 10625 54657 10628
rect 54691 10625 54703 10659
rect 54645 10619 54703 10625
rect 56137 10659 56195 10665
rect 56137 10625 56149 10659
rect 56183 10656 56195 10659
rect 56594 10656 56600 10668
rect 56183 10628 56600 10656
rect 56183 10625 56195 10628
rect 56137 10619 56195 10625
rect 56594 10616 56600 10628
rect 56652 10616 56658 10668
rect 56689 10659 56747 10665
rect 56689 10625 56701 10659
rect 56735 10625 56747 10659
rect 57422 10656 57428 10668
rect 57383 10628 57428 10656
rect 56689 10619 56747 10625
rect 51997 10591 52055 10597
rect 51997 10588 52009 10591
rect 46768 10560 52009 10588
rect 51997 10557 52009 10560
rect 52043 10557 52055 10591
rect 51997 10551 52055 10557
rect 52086 10548 52092 10600
rect 52144 10588 52150 10600
rect 52181 10591 52239 10597
rect 52181 10588 52193 10591
rect 52144 10560 52193 10588
rect 52144 10548 52150 10560
rect 52181 10557 52193 10560
rect 52227 10588 52239 10591
rect 52227 10560 53420 10588
rect 52227 10557 52239 10560
rect 52181 10551 52239 10557
rect 45646 10520 45652 10532
rect 44744 10492 45652 10520
rect 45646 10480 45652 10492
rect 45704 10480 45710 10532
rect 47581 10523 47639 10529
rect 47581 10520 47593 10523
rect 46676 10492 47593 10520
rect 42426 10452 42432 10464
rect 40972 10424 42432 10452
rect 39853 10415 39911 10421
rect 42426 10412 42432 10424
rect 42484 10412 42490 10464
rect 42521 10455 42579 10461
rect 42521 10421 42533 10455
rect 42567 10452 42579 10455
rect 43438 10452 43444 10464
rect 42567 10424 43444 10452
rect 42567 10421 42579 10424
rect 42521 10415 42579 10421
rect 43438 10412 43444 10424
rect 43496 10412 43502 10464
rect 43530 10412 43536 10464
rect 43588 10452 43594 10464
rect 44450 10452 44456 10464
rect 43588 10424 43633 10452
rect 44411 10424 44456 10452
rect 43588 10412 43594 10424
rect 44450 10412 44456 10424
rect 44508 10412 44514 10464
rect 45554 10412 45560 10464
rect 45612 10452 45618 10464
rect 46676 10452 46704 10492
rect 47581 10489 47593 10492
rect 47627 10489 47639 10523
rect 52546 10520 52552 10532
rect 47581 10483 47639 10489
rect 47688 10492 52552 10520
rect 45612 10424 46704 10452
rect 45612 10412 45618 10424
rect 46750 10412 46756 10464
rect 46808 10452 46814 10464
rect 47121 10455 47179 10461
rect 47121 10452 47133 10455
rect 46808 10424 47133 10452
rect 46808 10412 46814 10424
rect 47121 10421 47133 10424
rect 47167 10421 47179 10455
rect 47121 10415 47179 10421
rect 47210 10412 47216 10464
rect 47268 10452 47274 10464
rect 47688 10452 47716 10492
rect 52546 10480 52552 10492
rect 52604 10480 52610 10532
rect 52730 10520 52736 10532
rect 52691 10492 52736 10520
rect 52730 10480 52736 10492
rect 52788 10480 52794 10532
rect 47268 10424 47716 10452
rect 47268 10412 47274 10424
rect 48038 10412 48044 10464
rect 48096 10452 48102 10464
rect 49970 10452 49976 10464
rect 48096 10424 49976 10452
rect 48096 10412 48102 10424
rect 49970 10412 49976 10424
rect 50028 10412 50034 10464
rect 51537 10455 51595 10461
rect 51537 10421 51549 10455
rect 51583 10452 51595 10455
rect 53098 10452 53104 10464
rect 51583 10424 53104 10452
rect 51583 10421 51595 10424
rect 51537 10415 51595 10421
rect 53098 10412 53104 10424
rect 53156 10412 53162 10464
rect 53282 10452 53288 10464
rect 53243 10424 53288 10452
rect 53282 10412 53288 10424
rect 53340 10412 53346 10464
rect 53392 10452 53420 10560
rect 53742 10548 53748 10600
rect 53800 10588 53806 10600
rect 54389 10591 54447 10597
rect 54389 10588 54401 10591
rect 53800 10560 54401 10588
rect 53800 10548 53806 10560
rect 54389 10557 54401 10560
rect 54435 10557 54447 10591
rect 54389 10551 54447 10557
rect 55674 10548 55680 10600
rect 55732 10588 55738 10600
rect 56704 10588 56732 10619
rect 57422 10616 57428 10628
rect 57480 10616 57486 10668
rect 58621 10659 58679 10665
rect 58621 10625 58633 10659
rect 58667 10656 58679 10659
rect 58710 10656 58716 10668
rect 58667 10628 58716 10656
rect 58667 10625 58679 10628
rect 58621 10619 58679 10625
rect 58710 10616 58716 10628
rect 58768 10616 58774 10668
rect 58894 10656 58900 10668
rect 58855 10628 58900 10656
rect 58894 10616 58900 10628
rect 58952 10656 58958 10668
rect 59078 10656 59084 10668
rect 58952 10628 59084 10656
rect 58952 10616 58958 10628
rect 59078 10616 59084 10628
rect 59136 10616 59142 10668
rect 59648 10656 59676 10696
rect 59814 10684 59820 10696
rect 59872 10684 59878 10736
rect 60642 10724 60648 10736
rect 60108 10696 60648 10724
rect 60108 10656 60136 10696
rect 60642 10684 60648 10696
rect 60700 10684 60706 10736
rect 60826 10684 60832 10736
rect 60884 10724 60890 10736
rect 61565 10727 61623 10733
rect 61565 10724 61577 10727
rect 60884 10696 61577 10724
rect 60884 10684 60890 10696
rect 61565 10693 61577 10696
rect 61611 10724 61623 10727
rect 63678 10724 63684 10736
rect 61611 10696 63684 10724
rect 61611 10693 61623 10696
rect 61565 10687 61623 10693
rect 63678 10684 63684 10696
rect 63736 10724 63742 10736
rect 66640 10724 66668 10764
rect 67606 10764 70394 10792
rect 87651 10764 87696 10792
rect 67606 10724 67634 10764
rect 63736 10696 66116 10724
rect 66640 10696 67634 10724
rect 70366 10724 70394 10764
rect 87690 10752 87696 10764
rect 87748 10752 87754 10804
rect 87046 10724 87052 10736
rect 70366 10696 87052 10724
rect 63736 10684 63742 10696
rect 59648 10628 60136 10656
rect 60182 10616 60188 10668
rect 60240 10656 60246 10668
rect 60734 10656 60740 10668
rect 60240 10628 60740 10656
rect 60240 10616 60246 10628
rect 60734 10616 60740 10628
rect 60792 10616 60798 10668
rect 62206 10616 62212 10668
rect 62264 10656 62270 10668
rect 62301 10659 62359 10665
rect 62301 10656 62313 10659
rect 62264 10628 62313 10656
rect 62264 10616 62270 10628
rect 62301 10625 62313 10628
rect 62347 10625 62359 10659
rect 63218 10656 63224 10668
rect 63179 10628 63224 10656
rect 62301 10619 62359 10625
rect 63218 10616 63224 10628
rect 63276 10616 63282 10668
rect 63402 10656 63408 10668
rect 63363 10628 63408 10656
rect 63402 10616 63408 10628
rect 63460 10616 63466 10668
rect 63788 10665 63816 10696
rect 65536 10665 65564 10696
rect 63773 10659 63831 10665
rect 63773 10625 63785 10659
rect 63819 10625 63831 10659
rect 64029 10659 64087 10665
rect 64029 10656 64041 10659
rect 63773 10619 63831 10625
rect 63880 10628 64041 10656
rect 63034 10588 63040 10600
rect 55732 10560 56732 10588
rect 56796 10560 63040 10588
rect 55732 10548 55738 10560
rect 55398 10480 55404 10532
rect 55456 10520 55462 10532
rect 56796 10520 56824 10560
rect 63034 10548 63040 10560
rect 63092 10548 63098 10600
rect 63313 10591 63371 10597
rect 63313 10557 63325 10591
rect 63359 10588 63371 10591
rect 63880 10588 63908 10628
rect 64029 10625 64041 10628
rect 64075 10625 64087 10659
rect 64029 10619 64087 10625
rect 65521 10659 65579 10665
rect 65521 10625 65533 10659
rect 65567 10625 65579 10659
rect 65521 10619 65579 10625
rect 65610 10616 65616 10668
rect 65668 10656 65674 10668
rect 65777 10659 65835 10665
rect 65777 10656 65789 10659
rect 65668 10628 65789 10656
rect 65668 10616 65674 10628
rect 65777 10625 65789 10628
rect 65823 10625 65835 10659
rect 66088 10656 66116 10696
rect 87046 10684 87052 10696
rect 87104 10684 87110 10736
rect 66530 10656 66536 10668
rect 66088 10628 66536 10656
rect 65777 10619 65835 10625
rect 66530 10616 66536 10628
rect 66588 10656 66594 10668
rect 67542 10656 67548 10668
rect 66588 10628 67548 10656
rect 66588 10616 66594 10628
rect 67542 10616 67548 10628
rect 67600 10616 67606 10668
rect 87708 10656 87736 10752
rect 88245 10659 88303 10665
rect 88245 10656 88257 10659
rect 87708 10628 88257 10656
rect 88245 10625 88257 10628
rect 88291 10625 88303 10659
rect 88245 10619 88303 10625
rect 63359 10560 63908 10588
rect 63359 10557 63371 10560
rect 63313 10551 63371 10557
rect 55456 10492 56824 10520
rect 57241 10523 57299 10529
rect 55456 10480 55462 10492
rect 57241 10489 57253 10523
rect 57287 10520 57299 10523
rect 58066 10520 58072 10532
rect 57287 10492 58072 10520
rect 57287 10489 57299 10492
rect 57241 10483 57299 10489
rect 58066 10480 58072 10492
rect 58124 10480 58130 10532
rect 59170 10480 59176 10532
rect 59228 10520 59234 10532
rect 61930 10520 61936 10532
rect 59228 10492 61936 10520
rect 59228 10480 59234 10492
rect 61930 10480 61936 10492
rect 61988 10480 61994 10532
rect 62114 10520 62120 10532
rect 62075 10492 62120 10520
rect 62114 10480 62120 10492
rect 62172 10480 62178 10532
rect 64782 10480 64788 10532
rect 64840 10520 64846 10532
rect 64840 10492 65288 10520
rect 64840 10480 64846 10492
rect 55490 10452 55496 10464
rect 53392 10424 55496 10452
rect 55490 10412 55496 10424
rect 55548 10412 55554 10464
rect 55674 10412 55680 10464
rect 55732 10452 55738 10464
rect 55769 10455 55827 10461
rect 55769 10452 55781 10455
rect 55732 10424 55781 10452
rect 55732 10412 55738 10424
rect 55769 10421 55781 10424
rect 55815 10421 55827 10455
rect 55769 10415 55827 10421
rect 56594 10412 56600 10464
rect 56652 10452 56658 10464
rect 57790 10452 57796 10464
rect 56652 10424 57796 10452
rect 56652 10412 56658 10424
rect 57790 10412 57796 10424
rect 57848 10412 57854 10464
rect 58434 10452 58440 10464
rect 58395 10424 58440 10452
rect 58434 10412 58440 10424
rect 58492 10412 58498 10464
rect 58894 10412 58900 10464
rect 58952 10452 58958 10464
rect 64874 10452 64880 10464
rect 58952 10424 64880 10452
rect 58952 10412 58958 10424
rect 64874 10412 64880 10424
rect 64932 10412 64938 10464
rect 65150 10452 65156 10464
rect 65111 10424 65156 10452
rect 65150 10412 65156 10424
rect 65208 10412 65214 10464
rect 65260 10452 65288 10492
rect 66901 10455 66959 10461
rect 66901 10452 66913 10455
rect 65260 10424 66913 10452
rect 66901 10421 66913 10424
rect 66947 10421 66959 10455
rect 88058 10452 88064 10464
rect 88019 10424 88064 10452
rect 66901 10415 66959 10421
rect 88058 10412 88064 10424
rect 88116 10412 88122 10464
rect 1104 10362 88872 10384
rect 1104 10310 11924 10362
rect 11976 10310 11988 10362
rect 12040 10310 12052 10362
rect 12104 10310 12116 10362
rect 12168 10310 12180 10362
rect 12232 10310 33872 10362
rect 33924 10310 33936 10362
rect 33988 10310 34000 10362
rect 34052 10310 34064 10362
rect 34116 10310 34128 10362
rect 34180 10310 55820 10362
rect 55872 10310 55884 10362
rect 55936 10310 55948 10362
rect 56000 10310 56012 10362
rect 56064 10310 56076 10362
rect 56128 10310 77768 10362
rect 77820 10310 77832 10362
rect 77884 10310 77896 10362
rect 77948 10310 77960 10362
rect 78012 10310 78024 10362
rect 78076 10310 88872 10362
rect 1104 10288 88872 10310
rect 25038 10248 25044 10260
rect 24999 10220 25044 10248
rect 25038 10208 25044 10220
rect 25096 10208 25102 10260
rect 28905 10251 28963 10257
rect 28905 10217 28917 10251
rect 28951 10248 28963 10251
rect 29270 10248 29276 10260
rect 28951 10220 29276 10248
rect 28951 10217 28963 10220
rect 28905 10211 28963 10217
rect 29270 10208 29276 10220
rect 29328 10208 29334 10260
rect 32490 10208 32496 10260
rect 32548 10248 32554 10260
rect 32548 10220 33456 10248
rect 32548 10208 32554 10220
rect 33428 10180 33456 10220
rect 33502 10208 33508 10260
rect 33560 10248 33566 10260
rect 33873 10251 33931 10257
rect 33873 10248 33885 10251
rect 33560 10220 33885 10248
rect 33560 10208 33566 10220
rect 33873 10217 33885 10220
rect 33919 10248 33931 10251
rect 34238 10248 34244 10260
rect 33919 10220 34244 10248
rect 33919 10217 33931 10220
rect 33873 10211 33931 10217
rect 34238 10208 34244 10220
rect 34296 10208 34302 10260
rect 34330 10208 34336 10260
rect 34388 10248 34394 10260
rect 34388 10220 37872 10248
rect 34388 10208 34394 10220
rect 33428 10152 35112 10180
rect 33778 10072 33784 10124
rect 33836 10112 33842 10124
rect 35084 10112 35112 10152
rect 35158 10140 35164 10192
rect 35216 10180 35222 10192
rect 37737 10183 37795 10189
rect 37737 10180 37749 10183
rect 35216 10152 37749 10180
rect 35216 10140 35222 10152
rect 37737 10149 37749 10152
rect 37783 10149 37795 10183
rect 37844 10180 37872 10220
rect 38102 10208 38108 10260
rect 38160 10248 38166 10260
rect 38838 10248 38844 10260
rect 38160 10220 38844 10248
rect 38160 10208 38166 10220
rect 38838 10208 38844 10220
rect 38896 10208 38902 10260
rect 39206 10208 39212 10260
rect 39264 10248 39270 10260
rect 39853 10251 39911 10257
rect 39853 10248 39865 10251
rect 39264 10220 39865 10248
rect 39264 10208 39270 10220
rect 39853 10217 39865 10220
rect 39899 10217 39911 10251
rect 39853 10211 39911 10217
rect 40310 10208 40316 10260
rect 40368 10248 40374 10260
rect 40773 10251 40831 10257
rect 40773 10248 40785 10251
rect 40368 10220 40785 10248
rect 40368 10208 40374 10220
rect 40773 10217 40785 10220
rect 40819 10248 40831 10251
rect 42242 10248 42248 10260
rect 40819 10220 42248 10248
rect 40819 10217 40831 10220
rect 40773 10211 40831 10217
rect 42242 10208 42248 10220
rect 42300 10208 42306 10260
rect 42886 10208 42892 10260
rect 42944 10248 42950 10260
rect 43625 10251 43683 10257
rect 43625 10248 43637 10251
rect 42944 10220 43637 10248
rect 42944 10208 42950 10220
rect 43625 10217 43637 10220
rect 43671 10217 43683 10251
rect 43625 10211 43683 10217
rect 44450 10208 44456 10260
rect 44508 10248 44514 10260
rect 47118 10248 47124 10260
rect 44508 10220 47124 10248
rect 44508 10208 44514 10220
rect 47118 10208 47124 10220
rect 47176 10208 47182 10260
rect 47213 10251 47271 10257
rect 47213 10217 47225 10251
rect 47259 10217 47271 10251
rect 47213 10211 47271 10217
rect 49605 10251 49663 10257
rect 49605 10217 49617 10251
rect 49651 10248 49663 10251
rect 49694 10248 49700 10260
rect 49651 10220 49700 10248
rect 49651 10217 49663 10220
rect 49605 10211 49663 10217
rect 41966 10180 41972 10192
rect 37844 10152 41972 10180
rect 37737 10143 37795 10149
rect 41966 10140 41972 10152
rect 42024 10140 42030 10192
rect 45278 10180 45284 10192
rect 43272 10152 45284 10180
rect 39117 10115 39175 10121
rect 39117 10112 39129 10115
rect 33836 10084 35020 10112
rect 35084 10084 39129 10112
rect 33836 10072 33842 10084
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 21542 10044 21548 10056
rect 1627 10016 21548 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 21542 10004 21548 10016
rect 21600 10004 21606 10056
rect 25222 10044 25228 10056
rect 25183 10016 25228 10044
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 29086 10044 29092 10056
rect 29047 10016 29092 10044
rect 29086 10004 29092 10016
rect 29144 10004 29150 10056
rect 29546 10044 29552 10056
rect 29459 10016 29552 10044
rect 29546 10004 29552 10016
rect 29604 10044 29610 10056
rect 31754 10044 31760 10056
rect 29604 10016 31760 10044
rect 29604 10004 29610 10016
rect 31754 10004 31760 10016
rect 31812 10044 31818 10056
rect 32493 10047 32551 10053
rect 32493 10044 32505 10047
rect 31812 10016 32505 10044
rect 31812 10004 31818 10016
rect 32493 10013 32505 10016
rect 32539 10044 32551 10047
rect 33226 10044 33232 10056
rect 32539 10016 33232 10044
rect 32539 10013 32551 10016
rect 32493 10007 32551 10013
rect 33226 10004 33232 10016
rect 33284 10044 33290 10056
rect 34514 10044 34520 10056
rect 33284 10016 34520 10044
rect 33284 10004 33290 10016
rect 34514 10004 34520 10016
rect 34572 10004 34578 10056
rect 34882 10044 34888 10056
rect 34843 10016 34888 10044
rect 34882 10004 34888 10016
rect 34940 10004 34946 10056
rect 28074 9936 28080 9988
rect 28132 9976 28138 9988
rect 29794 9979 29852 9985
rect 29794 9976 29806 9979
rect 28132 9948 29806 9976
rect 28132 9936 28138 9948
rect 29794 9945 29806 9948
rect 29840 9945 29852 9979
rect 29794 9939 29852 9945
rect 32760 9979 32818 9985
rect 32760 9945 32772 9979
rect 32806 9976 32818 9979
rect 34992 9976 35020 10084
rect 39117 10081 39129 10084
rect 39163 10112 39175 10115
rect 39298 10112 39304 10124
rect 39163 10084 39304 10112
rect 39163 10081 39175 10084
rect 39117 10075 39175 10081
rect 39298 10072 39304 10084
rect 39356 10072 39362 10124
rect 40052 10084 40724 10112
rect 40052 10056 40080 10084
rect 35986 10044 35992 10056
rect 35947 10016 35992 10044
rect 35986 10004 35992 10016
rect 36044 10004 36050 10056
rect 37550 10004 37556 10056
rect 37608 10044 37614 10056
rect 40034 10044 40040 10056
rect 37608 10016 40040 10044
rect 37608 10004 37614 10016
rect 40034 10004 40040 10016
rect 40092 10004 40098 10056
rect 40126 10004 40132 10056
rect 40184 10044 40190 10056
rect 40696 10053 40724 10084
rect 40221 10047 40279 10053
rect 40221 10044 40233 10047
rect 40184 10016 40233 10044
rect 40184 10004 40190 10016
rect 40221 10013 40233 10016
rect 40267 10013 40279 10047
rect 40221 10007 40279 10013
rect 40313 10047 40371 10053
rect 40313 10013 40325 10047
rect 40359 10013 40371 10047
rect 40313 10007 40371 10013
rect 40681 10047 40739 10053
rect 40681 10013 40693 10047
rect 40727 10013 40739 10047
rect 40681 10007 40739 10013
rect 42245 10047 42303 10053
rect 42245 10013 42257 10047
rect 42291 10044 42303 10047
rect 42291 10016 42748 10044
rect 42291 10013 42303 10016
rect 42245 10007 42303 10013
rect 36449 9979 36507 9985
rect 32806 9948 34744 9976
rect 34992 9948 36400 9976
rect 32806 9945 32818 9948
rect 32760 9939 32818 9945
rect 1394 9908 1400 9920
rect 1355 9880 1400 9908
rect 1394 9868 1400 9880
rect 1452 9868 1458 9920
rect 28994 9868 29000 9920
rect 29052 9908 29058 9920
rect 30929 9911 30987 9917
rect 30929 9908 30941 9911
rect 29052 9880 30941 9908
rect 29052 9868 29058 9880
rect 30929 9877 30941 9880
rect 30975 9908 30987 9911
rect 34606 9908 34612 9920
rect 30975 9880 34612 9908
rect 30975 9877 30987 9880
rect 30929 9871 30987 9877
rect 34606 9868 34612 9880
rect 34664 9868 34670 9920
rect 34716 9917 34744 9948
rect 34701 9911 34759 9917
rect 34701 9877 34713 9911
rect 34747 9877 34759 9911
rect 35802 9908 35808 9920
rect 35763 9880 35808 9908
rect 34701 9871 34759 9877
rect 35802 9868 35808 9880
rect 35860 9868 35866 9920
rect 36372 9908 36400 9948
rect 36449 9945 36461 9979
rect 36495 9976 36507 9979
rect 38654 9976 38660 9988
rect 36495 9948 38660 9976
rect 36495 9945 36507 9948
rect 36449 9939 36507 9945
rect 38654 9936 38660 9948
rect 38712 9936 38718 9988
rect 40328 9976 40356 10007
rect 42720 9988 42748 10016
rect 42794 10004 42800 10056
rect 42852 10044 42858 10056
rect 43272 10044 43300 10152
rect 45278 10140 45284 10152
rect 45336 10140 45342 10192
rect 46658 10180 46664 10192
rect 46619 10152 46664 10180
rect 46658 10140 46664 10152
rect 46716 10180 46722 10192
rect 47228 10180 47256 10211
rect 49694 10208 49700 10220
rect 49752 10208 49758 10260
rect 51353 10251 51411 10257
rect 51353 10217 51365 10251
rect 51399 10248 51411 10251
rect 51902 10248 51908 10260
rect 51399 10220 51908 10248
rect 51399 10217 51411 10220
rect 51353 10211 51411 10217
rect 51902 10208 51908 10220
rect 51960 10208 51966 10260
rect 55490 10208 55496 10260
rect 55548 10248 55554 10260
rect 55548 10220 56272 10248
rect 55548 10208 55554 10220
rect 46716 10152 47256 10180
rect 47397 10183 47455 10189
rect 46716 10140 46722 10152
rect 47397 10149 47409 10183
rect 47443 10149 47455 10183
rect 47397 10143 47455 10149
rect 49053 10183 49111 10189
rect 49053 10149 49065 10183
rect 49099 10180 49111 10183
rect 49786 10180 49792 10192
rect 49099 10152 49792 10180
rect 49099 10149 49111 10152
rect 49053 10143 49111 10149
rect 42852 10016 43300 10044
rect 45281 10047 45339 10053
rect 42852 10004 42858 10016
rect 45281 10013 45293 10047
rect 45327 10044 45339 10047
rect 45370 10044 45376 10056
rect 45327 10016 45376 10044
rect 45327 10013 45339 10016
rect 45281 10007 45339 10013
rect 41690 9976 41696 9988
rect 38948 9948 41696 9976
rect 38102 9908 38108 9920
rect 36372 9880 38108 9908
rect 38102 9868 38108 9880
rect 38160 9868 38166 9920
rect 38194 9868 38200 9920
rect 38252 9908 38258 9920
rect 38565 9911 38623 9917
rect 38565 9908 38577 9911
rect 38252 9880 38577 9908
rect 38252 9868 38258 9880
rect 38565 9877 38577 9880
rect 38611 9877 38623 9911
rect 38565 9871 38623 9877
rect 38838 9868 38844 9920
rect 38896 9908 38902 9920
rect 38948 9917 38976 9948
rect 41690 9936 41696 9948
rect 41748 9936 41754 9988
rect 42512 9979 42570 9985
rect 42512 9945 42524 9979
rect 42558 9976 42570 9979
rect 42558 9948 42656 9976
rect 42558 9945 42570 9948
rect 42512 9939 42570 9945
rect 38933 9911 38991 9917
rect 38933 9908 38945 9911
rect 38896 9880 38945 9908
rect 38896 9868 38902 9880
rect 38933 9877 38945 9880
rect 38979 9877 38991 9911
rect 38933 9871 38991 9877
rect 39025 9911 39083 9917
rect 39025 9877 39037 9911
rect 39071 9908 39083 9911
rect 39298 9908 39304 9920
rect 39071 9880 39304 9908
rect 39071 9877 39083 9880
rect 39025 9871 39083 9877
rect 39298 9868 39304 9880
rect 39356 9868 39362 9920
rect 42628 9908 42656 9948
rect 42702 9936 42708 9988
rect 42760 9976 42766 9988
rect 45296 9976 45324 10007
rect 45370 10004 45376 10016
rect 45428 10004 45434 10056
rect 47412 10044 47440 10143
rect 49786 10140 49792 10152
rect 49844 10140 49850 10192
rect 53098 10180 53104 10192
rect 49896 10152 53104 10180
rect 49896 10112 49924 10152
rect 53098 10140 53104 10152
rect 53156 10140 53162 10192
rect 54113 10183 54171 10189
rect 54113 10149 54125 10183
rect 54159 10180 54171 10183
rect 55214 10180 55220 10192
rect 54159 10152 55220 10180
rect 54159 10149 54171 10152
rect 54113 10143 54171 10149
rect 55214 10140 55220 10152
rect 55272 10140 55278 10192
rect 56244 10180 56272 10220
rect 57422 10208 57428 10260
rect 57480 10248 57486 10260
rect 59449 10251 59507 10257
rect 59449 10248 59461 10251
rect 57480 10220 59461 10248
rect 57480 10208 57486 10220
rect 59449 10217 59461 10220
rect 59495 10217 59507 10251
rect 59449 10211 59507 10217
rect 60734 10208 60740 10260
rect 60792 10248 60798 10260
rect 61657 10251 61715 10257
rect 61657 10248 61669 10251
rect 60792 10220 61669 10248
rect 60792 10208 60798 10220
rect 61657 10217 61669 10220
rect 61703 10217 61715 10251
rect 61657 10211 61715 10217
rect 62209 10251 62267 10257
rect 62209 10217 62221 10251
rect 62255 10248 62267 10251
rect 64598 10248 64604 10260
rect 62255 10220 64604 10248
rect 62255 10217 62267 10220
rect 62209 10211 62267 10217
rect 64598 10208 64604 10220
rect 64656 10208 64662 10260
rect 64877 10251 64935 10257
rect 64877 10217 64889 10251
rect 64923 10248 64935 10251
rect 65610 10248 65616 10260
rect 64923 10220 65616 10248
rect 64923 10217 64935 10220
rect 64877 10211 64935 10217
rect 65610 10208 65616 10220
rect 65668 10208 65674 10260
rect 86586 10248 86592 10260
rect 70366 10220 86592 10248
rect 56244 10152 60734 10180
rect 45848 10016 47440 10044
rect 48286 10084 49924 10112
rect 45554 9985 45560 9988
rect 45548 9976 45560 9985
rect 42760 9948 45324 9976
rect 45515 9948 45560 9976
rect 42760 9936 42766 9948
rect 45548 9939 45560 9948
rect 45554 9936 45560 9939
rect 45612 9936 45618 9988
rect 45646 9936 45652 9988
rect 45704 9976 45710 9988
rect 45848 9976 45876 10016
rect 45704 9948 45876 9976
rect 45704 9936 45710 9948
rect 46750 9936 46756 9988
rect 46808 9976 46814 9988
rect 47029 9979 47087 9985
rect 47029 9976 47041 9979
rect 46808 9948 47041 9976
rect 46808 9936 46814 9948
rect 47029 9945 47041 9948
rect 47075 9945 47087 9979
rect 48286 9976 48314 10084
rect 49970 10072 49976 10124
rect 50028 10112 50034 10124
rect 50617 10115 50675 10121
rect 50617 10112 50629 10115
rect 50028 10084 50629 10112
rect 50028 10072 50034 10084
rect 50617 10081 50629 10084
rect 50663 10081 50675 10115
rect 50617 10075 50675 10081
rect 50709 10115 50767 10121
rect 50709 10081 50721 10115
rect 50755 10081 50767 10115
rect 53742 10112 53748 10124
rect 53703 10084 53748 10112
rect 50709 10075 50767 10081
rect 48958 10044 48964 10056
rect 48919 10016 48964 10044
rect 48958 10004 48964 10016
rect 49016 10004 49022 10056
rect 49513 10047 49571 10053
rect 49513 10013 49525 10047
rect 49559 10013 49571 10047
rect 49513 10007 49571 10013
rect 47029 9939 47087 9945
rect 47136 9948 48314 9976
rect 42978 9908 42984 9920
rect 42628 9880 42984 9908
rect 42978 9868 42984 9880
rect 43036 9868 43042 9920
rect 43438 9868 43444 9920
rect 43496 9908 43502 9920
rect 47136 9908 47164 9948
rect 43496 9880 47164 9908
rect 43496 9868 43502 9880
rect 47210 9868 47216 9920
rect 47268 9917 47274 9920
rect 47268 9911 47287 9917
rect 47275 9877 47287 9911
rect 47268 9871 47287 9877
rect 47268 9868 47274 9871
rect 47486 9868 47492 9920
rect 47544 9908 47550 9920
rect 49528 9908 49556 10007
rect 50062 10004 50068 10056
rect 50120 10044 50126 10056
rect 50724 10044 50752 10075
rect 53742 10072 53748 10084
rect 53800 10072 53806 10124
rect 53834 10072 53840 10124
rect 53892 10112 53898 10124
rect 54665 10115 54723 10121
rect 54665 10112 54677 10115
rect 53892 10084 54677 10112
rect 53892 10072 53898 10084
rect 54665 10081 54677 10084
rect 54711 10112 54723 10115
rect 55030 10112 55036 10124
rect 54711 10084 55036 10112
rect 54711 10081 54723 10084
rect 54665 10075 54723 10081
rect 55030 10072 55036 10084
rect 55088 10072 55094 10124
rect 55306 10112 55312 10124
rect 55267 10084 55312 10112
rect 55306 10072 55312 10084
rect 55364 10072 55370 10124
rect 58084 10121 58112 10152
rect 58069 10115 58127 10121
rect 58069 10081 58081 10115
rect 58115 10081 58127 10115
rect 60706 10112 60734 10152
rect 61930 10140 61936 10192
rect 61988 10180 61994 10192
rect 70366 10180 70394 10220
rect 86586 10208 86592 10220
rect 86644 10208 86650 10260
rect 61988 10152 70394 10180
rect 61988 10140 61994 10152
rect 61013 10115 61071 10121
rect 61013 10112 61025 10115
rect 58069 10075 58127 10081
rect 59004 10084 60596 10112
rect 60706 10084 61025 10112
rect 50120 10016 50752 10044
rect 50120 10004 50126 10016
rect 50982 10004 50988 10056
rect 51040 10044 51046 10056
rect 51261 10047 51319 10053
rect 51261 10044 51273 10047
rect 51040 10016 51273 10044
rect 51040 10004 51046 10016
rect 51261 10013 51273 10016
rect 51307 10013 51319 10047
rect 51261 10007 51319 10013
rect 51350 10004 51356 10056
rect 51408 10044 51414 10056
rect 51997 10047 52055 10053
rect 51997 10044 52009 10047
rect 51408 10016 52009 10044
rect 51408 10004 51414 10016
rect 51997 10013 52009 10016
rect 52043 10044 52055 10047
rect 52178 10044 52184 10056
rect 52043 10016 52184 10044
rect 52043 10013 52055 10016
rect 51997 10007 52055 10013
rect 52178 10004 52184 10016
rect 52236 10004 52242 10056
rect 53098 10004 53104 10056
rect 53156 10044 53162 10056
rect 57790 10044 57796 10056
rect 53156 10016 55720 10044
rect 57751 10016 57796 10044
rect 53156 10004 53162 10016
rect 49602 9936 49608 9988
rect 49660 9976 49666 9988
rect 54481 9979 54539 9985
rect 49660 9948 51074 9976
rect 49660 9936 49666 9948
rect 47544 9880 49556 9908
rect 47544 9868 47550 9880
rect 49694 9868 49700 9920
rect 49752 9908 49758 9920
rect 50157 9911 50215 9917
rect 50157 9908 50169 9911
rect 49752 9880 50169 9908
rect 49752 9868 49758 9880
rect 50157 9877 50169 9880
rect 50203 9877 50215 9911
rect 50522 9908 50528 9920
rect 50483 9880 50528 9908
rect 50157 9871 50215 9877
rect 50522 9868 50528 9880
rect 50580 9868 50586 9920
rect 51046 9908 51074 9948
rect 54481 9945 54493 9979
rect 54527 9976 54539 9979
rect 54527 9948 55352 9976
rect 54527 9945 54539 9948
rect 54481 9939 54539 9945
rect 54386 9908 54392 9920
rect 51046 9880 54392 9908
rect 54386 9868 54392 9880
rect 54444 9868 54450 9920
rect 54570 9908 54576 9920
rect 54531 9880 54576 9908
rect 54570 9868 54576 9880
rect 54628 9868 54634 9920
rect 55324 9908 55352 9948
rect 55398 9936 55404 9988
rect 55456 9976 55462 9988
rect 55554 9979 55612 9985
rect 55554 9976 55566 9979
rect 55456 9948 55566 9976
rect 55456 9936 55462 9948
rect 55554 9945 55566 9948
rect 55600 9945 55612 9979
rect 55692 9976 55720 10016
rect 57790 10004 57796 10016
rect 57848 10004 57854 10056
rect 57885 10047 57943 10053
rect 57885 10013 57897 10047
rect 57931 10044 57943 10047
rect 59004 10044 59032 10084
rect 57931 10016 59032 10044
rect 59081 10047 59139 10053
rect 57931 10013 57943 10016
rect 57885 10007 57943 10013
rect 59081 10013 59093 10047
rect 59127 10013 59139 10047
rect 59081 10007 59139 10013
rect 55692 9948 57974 9976
rect 55554 9939 55612 9945
rect 56226 9908 56232 9920
rect 55324 9880 56232 9908
rect 56226 9868 56232 9880
rect 56284 9908 56290 9920
rect 56689 9911 56747 9917
rect 56689 9908 56701 9911
rect 56284 9880 56701 9908
rect 56284 9868 56290 9880
rect 56689 9877 56701 9880
rect 56735 9877 56747 9911
rect 56689 9871 56747 9877
rect 57238 9868 57244 9920
rect 57296 9908 57302 9920
rect 57425 9911 57483 9917
rect 57425 9908 57437 9911
rect 57296 9880 57437 9908
rect 57296 9868 57302 9880
rect 57425 9877 57437 9880
rect 57471 9877 57483 9911
rect 57946 9908 57974 9948
rect 58158 9936 58164 9988
rect 58216 9976 58222 9988
rect 59096 9976 59124 10007
rect 59170 10004 59176 10056
rect 59228 10044 59234 10056
rect 59265 10047 59323 10053
rect 59265 10044 59277 10047
rect 59228 10016 59277 10044
rect 59228 10004 59234 10016
rect 59265 10013 59277 10016
rect 59311 10013 59323 10047
rect 59265 10007 59323 10013
rect 60001 10047 60059 10053
rect 60001 10013 60013 10047
rect 60047 10044 60059 10047
rect 60047 10016 60504 10044
rect 60047 10013 60059 10016
rect 60001 10007 60059 10013
rect 58216 9948 59124 9976
rect 58216 9936 58222 9948
rect 58618 9908 58624 9920
rect 57946 9880 58624 9908
rect 57425 9871 57483 9877
rect 58618 9868 58624 9880
rect 58676 9868 58682 9920
rect 58805 9911 58863 9917
rect 58805 9877 58817 9911
rect 58851 9908 58863 9911
rect 59188 9908 59216 10004
rect 59814 9908 59820 9920
rect 58851 9880 59216 9908
rect 59775 9880 59820 9908
rect 58851 9877 58863 9880
rect 58805 9871 58863 9877
rect 59814 9868 59820 9880
rect 59872 9868 59878 9920
rect 60476 9917 60504 10016
rect 60568 9976 60596 10084
rect 61013 10081 61025 10084
rect 61059 10081 61071 10115
rect 61013 10075 61071 10081
rect 64601 10115 64659 10121
rect 64601 10081 64613 10115
rect 64647 10112 64659 10115
rect 64690 10112 64696 10124
rect 64647 10084 64696 10112
rect 64647 10081 64659 10084
rect 64601 10075 64659 10081
rect 64690 10072 64696 10084
rect 64748 10072 64754 10124
rect 60826 10044 60832 10056
rect 60739 10016 60832 10044
rect 60826 10004 60832 10016
rect 60884 10044 60890 10056
rect 61565 10047 61623 10053
rect 61565 10044 61577 10047
rect 60884 10016 61577 10044
rect 60884 10004 60890 10016
rect 61565 10013 61577 10016
rect 61611 10013 61623 10047
rect 61565 10007 61623 10013
rect 62117 10047 62175 10053
rect 62117 10013 62129 10047
rect 62163 10044 62175 10047
rect 62298 10044 62304 10056
rect 62163 10016 62304 10044
rect 62163 10013 62175 10016
rect 62117 10007 62175 10013
rect 62298 10004 62304 10016
rect 62356 10004 62362 10056
rect 64230 10004 64236 10056
rect 64288 10044 64294 10056
rect 64509 10047 64567 10053
rect 64509 10044 64521 10047
rect 64288 10016 64521 10044
rect 64288 10004 64294 10016
rect 64509 10013 64521 10016
rect 64555 10044 64567 10047
rect 64782 10044 64788 10056
rect 64555 10016 64788 10044
rect 64555 10013 64567 10016
rect 64509 10007 64567 10013
rect 64782 10004 64788 10016
rect 64840 10004 64846 10056
rect 69014 9976 69020 9988
rect 60568 9948 69020 9976
rect 69014 9936 69020 9948
rect 69072 9936 69078 9988
rect 60461 9911 60519 9917
rect 60461 9877 60473 9911
rect 60507 9877 60519 9911
rect 60918 9908 60924 9920
rect 60879 9880 60924 9908
rect 60461 9871 60519 9877
rect 60918 9868 60924 9880
rect 60976 9868 60982 9920
rect 1104 9818 88872 9840
rect 1104 9766 22898 9818
rect 22950 9766 22962 9818
rect 23014 9766 23026 9818
rect 23078 9766 23090 9818
rect 23142 9766 23154 9818
rect 23206 9766 44846 9818
rect 44898 9766 44910 9818
rect 44962 9766 44974 9818
rect 45026 9766 45038 9818
rect 45090 9766 45102 9818
rect 45154 9766 66794 9818
rect 66846 9766 66858 9818
rect 66910 9766 66922 9818
rect 66974 9766 66986 9818
rect 67038 9766 67050 9818
rect 67102 9766 88872 9818
rect 1104 9744 88872 9766
rect 29086 9664 29092 9716
rect 29144 9704 29150 9716
rect 29733 9707 29791 9713
rect 29733 9704 29745 9707
rect 29144 9676 29745 9704
rect 29144 9664 29150 9676
rect 29733 9673 29745 9676
rect 29779 9673 29791 9707
rect 29733 9667 29791 9673
rect 30282 9664 30288 9716
rect 30340 9704 30346 9716
rect 32582 9704 32588 9716
rect 30340 9676 32588 9704
rect 30340 9664 30346 9676
rect 32582 9664 32588 9676
rect 32640 9664 32646 9716
rect 34514 9664 34520 9716
rect 34572 9664 34578 9716
rect 36262 9664 36268 9716
rect 36320 9704 36326 9716
rect 36541 9707 36599 9713
rect 36541 9704 36553 9707
rect 36320 9676 36553 9704
rect 36320 9664 36326 9676
rect 36541 9673 36553 9676
rect 36587 9673 36599 9707
rect 37642 9704 37648 9716
rect 37603 9676 37648 9704
rect 36541 9667 36599 9673
rect 37642 9664 37648 9676
rect 37700 9664 37706 9716
rect 38378 9664 38384 9716
rect 38436 9704 38442 9716
rect 49418 9704 49424 9716
rect 38436 9676 49424 9704
rect 38436 9664 38442 9676
rect 49418 9664 49424 9676
rect 49476 9664 49482 9716
rect 49694 9704 49700 9716
rect 49528 9676 49700 9704
rect 33502 9636 33508 9648
rect 33463 9608 33508 9636
rect 33502 9596 33508 9608
rect 33560 9596 33566 9648
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 30101 9571 30159 9577
rect 30101 9568 30113 9571
rect 15436 9540 30113 9568
rect 15436 9528 15442 9540
rect 30101 9537 30113 9540
rect 30147 9568 30159 9571
rect 31110 9568 31116 9580
rect 30147 9540 31116 9568
rect 30147 9537 30159 9540
rect 30101 9531 30159 9537
rect 31110 9528 31116 9540
rect 31168 9528 31174 9580
rect 34532 9568 34560 9664
rect 34606 9596 34612 9648
rect 34664 9636 34670 9648
rect 35428 9639 35486 9645
rect 34664 9608 35296 9636
rect 34664 9596 34670 9608
rect 35158 9568 35164 9580
rect 34532 9540 35164 9568
rect 35158 9528 35164 9540
rect 35216 9528 35222 9580
rect 35268 9568 35296 9608
rect 35428 9605 35440 9639
rect 35474 9636 35486 9639
rect 35802 9636 35808 9648
rect 35474 9608 35808 9636
rect 35474 9605 35486 9608
rect 35428 9599 35486 9605
rect 35802 9596 35808 9608
rect 35860 9596 35866 9648
rect 37277 9639 37335 9645
rect 37277 9605 37289 9639
rect 37323 9636 37335 9639
rect 38286 9636 38292 9648
rect 37323 9608 38292 9636
rect 37323 9605 37335 9608
rect 37277 9599 37335 9605
rect 38286 9596 38292 9608
rect 38344 9596 38350 9648
rect 45189 9639 45247 9645
rect 38580 9608 40356 9636
rect 35710 9568 35716 9580
rect 35268 9540 35716 9568
rect 35710 9528 35716 9540
rect 35768 9568 35774 9580
rect 37461 9571 37519 9577
rect 35768 9540 37412 9568
rect 35768 9528 35774 9540
rect 30190 9500 30196 9512
rect 30151 9472 30196 9500
rect 30190 9460 30196 9472
rect 30248 9460 30254 9512
rect 30282 9460 30288 9512
rect 30340 9500 30346 9512
rect 33597 9503 33655 9509
rect 33597 9500 33609 9503
rect 30340 9472 30385 9500
rect 31726 9472 33609 9500
rect 30340 9460 30346 9472
rect 23566 9392 23572 9444
rect 23624 9432 23630 9444
rect 31726 9432 31754 9472
rect 33597 9469 33609 9472
rect 33643 9469 33655 9503
rect 33778 9500 33784 9512
rect 33739 9472 33784 9500
rect 33597 9463 33655 9469
rect 33778 9460 33784 9472
rect 33836 9460 33842 9512
rect 37384 9500 37412 9540
rect 37461 9537 37473 9571
rect 37507 9568 37519 9571
rect 37550 9568 37556 9580
rect 37507 9540 37556 9568
rect 37507 9537 37519 9540
rect 37461 9531 37519 9537
rect 37550 9528 37556 9540
rect 37608 9528 37614 9580
rect 37737 9571 37795 9577
rect 37737 9537 37749 9571
rect 37783 9537 37795 9571
rect 37737 9531 37795 9537
rect 37752 9500 37780 9531
rect 38010 9528 38016 9580
rect 38068 9568 38074 9580
rect 38580 9577 38608 9608
rect 40328 9580 40356 9608
rect 45189 9605 45201 9639
rect 45235 9636 45247 9639
rect 47394 9636 47400 9648
rect 45235 9608 47400 9636
rect 45235 9605 45247 9608
rect 45189 9599 45247 9605
rect 47394 9596 47400 9608
rect 47452 9596 47458 9648
rect 38838 9577 38844 9580
rect 38565 9571 38623 9577
rect 38565 9568 38577 9571
rect 38068 9540 38577 9568
rect 38068 9528 38074 9540
rect 38565 9537 38577 9540
rect 38611 9537 38623 9571
rect 38565 9531 38623 9537
rect 38832 9531 38844 9577
rect 38896 9568 38902 9580
rect 40310 9568 40316 9580
rect 38896 9540 38932 9568
rect 40223 9540 40316 9568
rect 38838 9528 38844 9531
rect 38896 9528 38902 9540
rect 40310 9528 40316 9540
rect 40368 9528 40374 9580
rect 40402 9528 40408 9580
rect 40460 9568 40466 9580
rect 40569 9571 40627 9577
rect 40569 9568 40581 9571
rect 40460 9540 40581 9568
rect 40460 9528 40466 9540
rect 40569 9537 40581 9540
rect 40615 9537 40627 9571
rect 40569 9531 40627 9537
rect 42613 9571 42671 9577
rect 42613 9537 42625 9571
rect 42659 9568 42671 9571
rect 42886 9568 42892 9580
rect 42659 9540 42892 9568
rect 42659 9537 42671 9540
rect 42613 9531 42671 9537
rect 42886 9528 42892 9540
rect 42944 9528 42950 9580
rect 44082 9528 44088 9580
rect 44140 9568 44146 9580
rect 45097 9571 45155 9577
rect 45097 9568 45109 9571
rect 44140 9540 45109 9568
rect 44140 9528 44146 9540
rect 45097 9537 45109 9540
rect 45143 9537 45155 9571
rect 45097 9531 45155 9537
rect 45830 9528 45836 9580
rect 45888 9568 45894 9580
rect 45997 9571 46055 9577
rect 45997 9568 46009 9571
rect 45888 9540 46009 9568
rect 45888 9528 45894 9540
rect 45997 9537 46009 9540
rect 46043 9537 46055 9571
rect 45997 9531 46055 9537
rect 49237 9571 49295 9577
rect 49237 9537 49249 9571
rect 49283 9568 49295 9571
rect 49528 9568 49556 9676
rect 49694 9664 49700 9676
rect 49752 9664 49758 9716
rect 49786 9664 49792 9716
rect 49844 9704 49850 9716
rect 50798 9704 50804 9716
rect 49844 9676 50804 9704
rect 49844 9664 49850 9676
rect 50798 9664 50804 9676
rect 50856 9664 50862 9716
rect 50982 9704 50988 9716
rect 50895 9676 50988 9704
rect 50982 9664 50988 9676
rect 51040 9664 51046 9716
rect 54113 9707 54171 9713
rect 54113 9673 54125 9707
rect 54159 9704 54171 9707
rect 54294 9704 54300 9716
rect 54159 9676 54300 9704
rect 54159 9673 54171 9676
rect 54113 9667 54171 9673
rect 54294 9664 54300 9676
rect 54352 9664 54358 9716
rect 54478 9704 54484 9716
rect 54439 9676 54484 9704
rect 54478 9664 54484 9676
rect 54536 9664 54542 9716
rect 54570 9664 54576 9716
rect 54628 9704 54634 9716
rect 55401 9707 55459 9713
rect 54628 9676 55352 9704
rect 54628 9664 54634 9676
rect 50154 9636 50160 9648
rect 49620 9608 50160 9636
rect 49620 9577 49648 9608
rect 50154 9596 50160 9608
rect 50212 9596 50218 9648
rect 50522 9596 50528 9648
rect 50580 9636 50586 9648
rect 51000 9636 51028 9664
rect 50580 9608 51028 9636
rect 50580 9596 50586 9608
rect 51166 9596 51172 9648
rect 51224 9636 51230 9648
rect 51445 9639 51503 9645
rect 51445 9636 51457 9639
rect 51224 9608 51457 9636
rect 51224 9596 51230 9608
rect 51445 9605 51457 9608
rect 51491 9605 51503 9639
rect 53742 9636 53748 9648
rect 51445 9599 51503 9605
rect 52748 9608 53748 9636
rect 52748 9580 52776 9608
rect 53742 9596 53748 9608
rect 53800 9596 53806 9648
rect 55030 9596 55036 9648
rect 55088 9636 55094 9648
rect 55324 9636 55352 9676
rect 55401 9673 55413 9707
rect 55447 9704 55459 9707
rect 55674 9704 55680 9716
rect 55447 9676 55680 9704
rect 55447 9673 55459 9676
rect 55401 9667 55459 9673
rect 55674 9664 55680 9676
rect 55732 9664 55738 9716
rect 59262 9704 59268 9716
rect 55784 9676 59268 9704
rect 55784 9636 55812 9676
rect 59262 9664 59268 9676
rect 59320 9664 59326 9716
rect 60826 9704 60832 9716
rect 60787 9676 60832 9704
rect 60826 9664 60832 9676
rect 60884 9664 60890 9716
rect 64443 9707 64501 9713
rect 64443 9673 64455 9707
rect 64489 9704 64501 9707
rect 64690 9704 64696 9716
rect 64489 9676 64696 9704
rect 64489 9673 64501 9676
rect 64443 9667 64501 9673
rect 64690 9664 64696 9676
rect 64748 9664 64754 9716
rect 68189 9707 68247 9713
rect 68189 9673 68201 9707
rect 68235 9673 68247 9707
rect 68189 9667 68247 9673
rect 55088 9608 55260 9636
rect 55324 9608 55812 9636
rect 59716 9639 59774 9645
rect 55088 9596 55094 9608
rect 49283 9540 49556 9568
rect 49605 9571 49663 9577
rect 49283 9537 49295 9540
rect 49237 9531 49295 9537
rect 49605 9537 49617 9571
rect 49651 9537 49663 9571
rect 49861 9571 49919 9577
rect 49861 9568 49873 9571
rect 49605 9531 49663 9537
rect 49712 9540 49873 9568
rect 37384 9472 37780 9500
rect 42705 9503 42763 9509
rect 42705 9469 42717 9503
rect 42751 9469 42763 9503
rect 42978 9500 42984 9512
rect 42939 9472 42984 9500
rect 42705 9463 42763 9469
rect 23624 9404 31754 9432
rect 33137 9435 33195 9441
rect 23624 9392 23630 9404
rect 33137 9401 33149 9435
rect 33183 9432 33195 9435
rect 34882 9432 34888 9444
rect 33183 9404 34888 9432
rect 33183 9401 33195 9404
rect 33137 9395 33195 9401
rect 34882 9392 34888 9404
rect 34940 9392 34946 9444
rect 42720 9432 42748 9463
rect 42978 9460 42984 9472
rect 43036 9460 43042 9512
rect 45554 9460 45560 9512
rect 45612 9500 45618 9512
rect 45741 9503 45799 9509
rect 45741 9500 45753 9503
rect 45612 9472 45753 9500
rect 45612 9460 45618 9472
rect 45741 9469 45753 9472
rect 45787 9469 45799 9503
rect 49712 9500 49740 9540
rect 49861 9537 49873 9540
rect 49907 9537 49919 9571
rect 49861 9531 49919 9537
rect 51353 9571 51411 9577
rect 51353 9537 51365 9571
rect 51399 9537 51411 9571
rect 52730 9568 52736 9580
rect 52643 9540 52736 9568
rect 51353 9531 51411 9537
rect 45741 9463 45799 9469
rect 49068 9472 49740 9500
rect 51368 9500 51396 9531
rect 52730 9528 52736 9540
rect 52788 9528 52794 9580
rect 53000 9571 53058 9577
rect 53000 9537 53012 9571
rect 53046 9568 53058 9571
rect 53282 9568 53288 9580
rect 53046 9540 53288 9568
rect 53046 9537 53058 9540
rect 53000 9531 53058 9537
rect 53282 9528 53288 9540
rect 53340 9528 53346 9580
rect 54665 9571 54723 9577
rect 54665 9537 54677 9571
rect 54711 9568 54723 9571
rect 55232 9568 55260 9608
rect 59716 9605 59728 9639
rect 59762 9636 59774 9639
rect 59814 9636 59820 9648
rect 59762 9608 59820 9636
rect 59762 9605 59774 9608
rect 59716 9599 59774 9605
rect 59814 9596 59820 9608
rect 59872 9596 59878 9648
rect 64230 9636 64236 9648
rect 64191 9608 64236 9636
rect 64230 9596 64236 9608
rect 64288 9596 64294 9648
rect 68204 9636 68232 9667
rect 68204 9608 68692 9636
rect 57238 9568 57244 9580
rect 54711 9540 55076 9568
rect 55232 9540 55628 9568
rect 57199 9540 57244 9568
rect 54711 9537 54723 9540
rect 54665 9531 54723 9537
rect 51368 9472 52776 9500
rect 43990 9432 43996 9444
rect 42720 9404 43996 9432
rect 43990 9392 43996 9404
rect 44048 9392 44054 9444
rect 38562 9324 38568 9376
rect 38620 9364 38626 9376
rect 39298 9364 39304 9376
rect 38620 9336 39304 9364
rect 38620 9324 38626 9336
rect 39298 9324 39304 9336
rect 39356 9324 39362 9376
rect 39945 9367 40003 9373
rect 39945 9333 39957 9367
rect 39991 9364 40003 9367
rect 40218 9364 40224 9376
rect 39991 9336 40224 9364
rect 39991 9333 40003 9336
rect 39945 9327 40003 9333
rect 40218 9324 40224 9336
rect 40276 9324 40282 9376
rect 41690 9364 41696 9376
rect 41651 9336 41696 9364
rect 41690 9324 41696 9336
rect 41748 9324 41754 9376
rect 45756 9364 45784 9463
rect 47121 9435 47179 9441
rect 47121 9401 47133 9435
rect 47167 9432 47179 9435
rect 47486 9432 47492 9444
rect 47167 9404 47492 9432
rect 47167 9401 47179 9404
rect 47121 9395 47179 9401
rect 47486 9392 47492 9404
rect 47544 9392 47550 9444
rect 49068 9441 49096 9472
rect 49053 9435 49111 9441
rect 49053 9401 49065 9435
rect 49099 9401 49111 9435
rect 49053 9395 49111 9401
rect 46382 9364 46388 9376
rect 45756 9336 46388 9364
rect 46382 9324 46388 9336
rect 46440 9324 46446 9376
rect 48590 9324 48596 9376
rect 48648 9364 48654 9376
rect 52638 9364 52644 9376
rect 48648 9336 52644 9364
rect 48648 9324 48654 9336
rect 52638 9324 52644 9336
rect 52696 9324 52702 9376
rect 52748 9364 52776 9472
rect 55048 9441 55076 9540
rect 55600 9509 55628 9540
rect 57238 9528 57244 9540
rect 57296 9528 57302 9580
rect 59446 9568 59452 9580
rect 59407 9540 59452 9568
rect 59446 9528 59452 9540
rect 59504 9528 59510 9580
rect 68186 9528 68192 9580
rect 68244 9568 68250 9580
rect 68373 9571 68431 9577
rect 68373 9568 68385 9571
rect 68244 9540 68385 9568
rect 68244 9528 68250 9540
rect 68373 9537 68385 9540
rect 68419 9537 68431 9571
rect 68664 9568 68692 9608
rect 69017 9571 69075 9577
rect 69017 9568 69029 9571
rect 68664 9540 69029 9568
rect 68373 9531 68431 9537
rect 69017 9537 69029 9540
rect 69063 9537 69075 9571
rect 69017 9531 69075 9537
rect 55493 9503 55551 9509
rect 55493 9500 55505 9503
rect 55416 9472 55505 9500
rect 55033 9435 55091 9441
rect 55033 9401 55045 9435
rect 55079 9401 55091 9435
rect 55033 9395 55091 9401
rect 53098 9364 53104 9376
rect 52748 9336 53104 9364
rect 53098 9324 53104 9336
rect 53156 9324 53162 9376
rect 55416 9364 55444 9472
rect 55493 9469 55505 9472
rect 55539 9469 55551 9503
rect 55493 9463 55551 9469
rect 55585 9503 55643 9509
rect 55585 9469 55597 9503
rect 55631 9469 55643 9503
rect 55585 9463 55643 9469
rect 63402 9460 63408 9512
rect 63460 9500 63466 9512
rect 63460 9472 64644 9500
rect 63460 9460 63466 9472
rect 57054 9432 57060 9444
rect 57015 9404 57060 9432
rect 57054 9392 57060 9404
rect 57112 9392 57118 9444
rect 64616 9441 64644 9472
rect 67542 9460 67548 9512
rect 67600 9500 67606 9512
rect 68741 9503 68799 9509
rect 68741 9500 68753 9503
rect 67600 9472 68753 9500
rect 67600 9460 67606 9472
rect 68741 9469 68753 9472
rect 68787 9469 68799 9503
rect 68741 9463 68799 9469
rect 64601 9435 64659 9441
rect 64601 9401 64613 9435
rect 64647 9401 64659 9435
rect 64601 9395 64659 9401
rect 63402 9364 63408 9376
rect 55416 9336 63408 9364
rect 63402 9324 63408 9336
rect 63460 9324 63466 9376
rect 64417 9367 64475 9373
rect 64417 9333 64429 9367
rect 64463 9364 64475 9367
rect 65150 9364 65156 9376
rect 64463 9336 65156 9364
rect 64463 9333 64475 9336
rect 64417 9327 64475 9333
rect 65150 9324 65156 9336
rect 65208 9324 65214 9376
rect 68278 9324 68284 9376
rect 68336 9364 68342 9376
rect 70121 9367 70179 9373
rect 70121 9364 70133 9367
rect 68336 9336 70133 9364
rect 68336 9324 68342 9336
rect 70121 9333 70133 9336
rect 70167 9333 70179 9367
rect 70121 9327 70179 9333
rect 1104 9274 88872 9296
rect 1104 9222 11924 9274
rect 11976 9222 11988 9274
rect 12040 9222 12052 9274
rect 12104 9222 12116 9274
rect 12168 9222 12180 9274
rect 12232 9222 33872 9274
rect 33924 9222 33936 9274
rect 33988 9222 34000 9274
rect 34052 9222 34064 9274
rect 34116 9222 34128 9274
rect 34180 9222 55820 9274
rect 55872 9222 55884 9274
rect 55936 9222 55948 9274
rect 56000 9222 56012 9274
rect 56064 9222 56076 9274
rect 56128 9222 77768 9274
rect 77820 9222 77832 9274
rect 77884 9222 77896 9274
rect 77948 9222 77960 9274
rect 78012 9222 78024 9274
rect 78076 9222 88872 9274
rect 1104 9200 88872 9222
rect 35986 9120 35992 9172
rect 36044 9160 36050 9172
rect 36265 9163 36323 9169
rect 36265 9160 36277 9163
rect 36044 9132 36277 9160
rect 36044 9120 36050 9132
rect 36265 9129 36277 9132
rect 36311 9129 36323 9163
rect 37366 9160 37372 9172
rect 37327 9132 37372 9160
rect 36265 9123 36323 9129
rect 37366 9120 37372 9132
rect 37424 9120 37430 9172
rect 38657 9163 38715 9169
rect 38657 9129 38669 9163
rect 38703 9160 38715 9163
rect 38838 9160 38844 9172
rect 38703 9132 38844 9160
rect 38703 9129 38715 9132
rect 38657 9123 38715 9129
rect 38838 9120 38844 9132
rect 38896 9120 38902 9172
rect 40862 9120 40868 9172
rect 40920 9160 40926 9172
rect 41322 9160 41328 9172
rect 40920 9132 41328 9160
rect 40920 9120 40926 9132
rect 41322 9120 41328 9132
rect 41380 9160 41386 9172
rect 44082 9160 44088 9172
rect 41380 9132 43944 9160
rect 44043 9132 44088 9160
rect 41380 9120 41386 9132
rect 37734 9092 37740 9104
rect 37660 9064 37740 9092
rect 33778 8984 33784 9036
rect 33836 9024 33842 9036
rect 36817 9027 36875 9033
rect 36817 9024 36829 9027
rect 33836 8996 36829 9024
rect 33836 8984 33842 8996
rect 36817 8993 36829 8996
rect 36863 9024 36875 9027
rect 37660 9024 37688 9064
rect 37734 9052 37740 9064
rect 37792 9052 37798 9104
rect 40126 9024 40132 9036
rect 36863 8996 37688 9024
rect 37752 8996 40132 9024
rect 36863 8993 36875 8996
rect 36817 8987 36875 8993
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 36262 8916 36268 8968
rect 36320 8956 36326 8968
rect 36633 8959 36691 8965
rect 36633 8956 36645 8959
rect 36320 8928 36645 8956
rect 36320 8916 36326 8928
rect 36633 8925 36645 8928
rect 36679 8925 36691 8959
rect 37550 8956 37556 8968
rect 37511 8928 37556 8956
rect 36633 8919 36691 8925
rect 37550 8916 37556 8928
rect 37608 8916 37614 8968
rect 37642 8916 37648 8968
rect 37700 8956 37706 8968
rect 37752 8965 37780 8996
rect 40126 8984 40132 8996
rect 40184 8984 40190 9036
rect 40310 8984 40316 9036
rect 40368 9024 40374 9036
rect 42702 9024 42708 9036
rect 40368 8996 42708 9024
rect 40368 8984 40374 8996
rect 42702 8984 42708 8996
rect 42760 8984 42766 9036
rect 43916 9024 43944 9132
rect 44082 9120 44088 9132
rect 44140 9120 44146 9172
rect 45830 9160 45836 9172
rect 45791 9132 45836 9160
rect 45830 9120 45836 9132
rect 45888 9120 45894 9172
rect 48130 9160 48136 9172
rect 48091 9132 48136 9160
rect 48130 9120 48136 9132
rect 48188 9120 48194 9172
rect 48406 9120 48412 9172
rect 48464 9160 48470 9172
rect 51721 9163 51779 9169
rect 51721 9160 51733 9163
rect 48464 9132 51733 9160
rect 48464 9120 48470 9132
rect 51721 9129 51733 9132
rect 51767 9160 51779 9163
rect 55309 9163 55367 9169
rect 51767 9132 54432 9160
rect 51767 9129 51779 9132
rect 51721 9123 51779 9129
rect 47765 9095 47823 9101
rect 47765 9061 47777 9095
rect 47811 9092 47823 9095
rect 54404 9092 54432 9132
rect 55309 9129 55321 9163
rect 55355 9160 55367 9163
rect 55398 9160 55404 9172
rect 55355 9132 55404 9160
rect 55355 9129 55367 9132
rect 55309 9123 55367 9129
rect 55398 9120 55404 9132
rect 55456 9120 55462 9172
rect 68186 9160 68192 9172
rect 68147 9132 68192 9160
rect 68186 9120 68192 9132
rect 68244 9120 68250 9172
rect 47811 9064 48544 9092
rect 54404 9064 60734 9092
rect 47811 9061 47823 9064
rect 47765 9055 47823 9061
rect 43916 8996 46520 9024
rect 37737 8959 37795 8965
rect 37737 8956 37749 8959
rect 37700 8928 37749 8956
rect 37700 8916 37706 8928
rect 37737 8925 37749 8928
rect 37783 8925 37795 8959
rect 37737 8919 37795 8925
rect 37829 8959 37887 8965
rect 37829 8925 37841 8959
rect 37875 8925 37887 8959
rect 37829 8919 37887 8925
rect 31110 8848 31116 8900
rect 31168 8888 31174 8900
rect 37844 8888 37872 8919
rect 38746 8916 38752 8968
rect 38804 8956 38810 8968
rect 38841 8959 38899 8965
rect 38841 8956 38853 8959
rect 38804 8928 38853 8956
rect 38804 8916 38810 8928
rect 38841 8925 38853 8928
rect 38887 8925 38899 8959
rect 38841 8919 38899 8925
rect 42337 8959 42395 8965
rect 42337 8925 42349 8959
rect 42383 8956 42395 8959
rect 42794 8956 42800 8968
rect 42383 8928 42800 8956
rect 42383 8925 42395 8928
rect 42337 8919 42395 8925
rect 42794 8916 42800 8928
rect 42852 8916 42858 8968
rect 46017 8959 46075 8965
rect 46017 8925 46029 8959
rect 46063 8956 46075 8959
rect 46106 8956 46112 8968
rect 46063 8928 46112 8956
rect 46063 8925 46075 8928
rect 46017 8919 46075 8925
rect 46106 8916 46112 8928
rect 46164 8916 46170 8968
rect 46382 8956 46388 8968
rect 46343 8928 46388 8956
rect 46382 8916 46388 8928
rect 46440 8916 46446 8968
rect 46492 8956 46520 8996
rect 48406 8956 48412 8968
rect 46492 8928 48412 8956
rect 48406 8916 48412 8928
rect 48464 8916 48470 8968
rect 48516 8965 48544 9064
rect 48590 8984 48596 9036
rect 48648 9024 48654 9036
rect 48685 9027 48743 9033
rect 48685 9024 48697 9027
rect 48648 8996 48697 9024
rect 48648 8984 48654 8996
rect 48685 8993 48697 8996
rect 48731 8993 48743 9027
rect 52730 9024 52736 9036
rect 48685 8987 48743 8993
rect 50172 8996 52736 9024
rect 50172 8968 50200 8996
rect 52730 8984 52736 8996
rect 52788 8984 52794 9036
rect 48501 8959 48559 8965
rect 48501 8925 48513 8959
rect 48547 8956 48559 8959
rect 48958 8956 48964 8968
rect 48547 8928 48964 8956
rect 48547 8925 48559 8928
rect 48501 8919 48559 8925
rect 48958 8916 48964 8928
rect 49016 8916 49022 8968
rect 50154 8956 50160 8968
rect 50115 8928 50160 8956
rect 50154 8916 50160 8928
rect 50212 8916 50218 8968
rect 50246 8916 50252 8968
rect 50304 8956 50310 8968
rect 50433 8959 50491 8965
rect 50433 8956 50445 8959
rect 50304 8928 50445 8956
rect 50304 8916 50310 8928
rect 50433 8925 50445 8928
rect 50479 8925 50491 8959
rect 52362 8956 52368 8968
rect 52323 8928 52368 8956
rect 50433 8919 50491 8925
rect 52362 8916 52368 8928
rect 52420 8916 52426 8968
rect 55214 8916 55220 8968
rect 55272 8956 55278 8968
rect 55493 8959 55551 8965
rect 55493 8956 55505 8959
rect 55272 8928 55505 8956
rect 55272 8916 55278 8928
rect 55493 8925 55505 8928
rect 55539 8925 55551 8959
rect 55493 8919 55551 8925
rect 42950 8891 43008 8897
rect 42950 8888 42962 8891
rect 31168 8860 37872 8888
rect 42168 8860 42962 8888
rect 31168 8848 31174 8860
rect 1397 8823 1455 8829
rect 1397 8789 1409 8823
rect 1443 8820 1455 8823
rect 23382 8820 23388 8832
rect 1443 8792 23388 8820
rect 1443 8789 1455 8792
rect 1397 8783 1455 8789
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 36722 8820 36728 8832
rect 36683 8792 36728 8820
rect 36722 8780 36728 8792
rect 36780 8780 36786 8832
rect 42168 8829 42196 8860
rect 42950 8857 42962 8860
rect 42996 8857 43008 8891
rect 42950 8851 43008 8857
rect 46474 8848 46480 8900
rect 46532 8888 46538 8900
rect 46630 8891 46688 8897
rect 46630 8888 46642 8891
rect 46532 8860 46642 8888
rect 46532 8848 46538 8860
rect 46630 8857 46642 8860
rect 46676 8857 46688 8891
rect 46630 8851 46688 8857
rect 46934 8848 46940 8900
rect 46992 8888 46998 8900
rect 48593 8891 48651 8897
rect 48593 8888 48605 8891
rect 46992 8860 48605 8888
rect 46992 8848 46998 8860
rect 48593 8857 48605 8860
rect 48639 8857 48651 8891
rect 52978 8891 53036 8897
rect 52978 8888 52990 8891
rect 48593 8851 48651 8857
rect 52196 8860 52990 8888
rect 42153 8823 42211 8829
rect 42153 8789 42165 8823
rect 42199 8789 42211 8823
rect 42153 8783 42211 8789
rect 50062 8780 50068 8832
rect 50120 8820 50126 8832
rect 50798 8820 50804 8832
rect 50120 8792 50804 8820
rect 50120 8780 50126 8792
rect 50798 8780 50804 8792
rect 50856 8780 50862 8832
rect 52196 8829 52224 8860
rect 52978 8857 52990 8860
rect 53024 8857 53036 8891
rect 60706 8888 60734 9064
rect 60918 9052 60924 9104
rect 60976 9092 60982 9104
rect 60976 9064 84194 9092
rect 60976 9052 60982 9064
rect 67542 8984 67548 9036
rect 67600 9024 67606 9036
rect 68741 9027 68799 9033
rect 68741 9024 68753 9027
rect 67600 8996 68753 9024
rect 67600 8984 67606 8996
rect 68741 8993 68753 8996
rect 68787 8993 68799 9027
rect 84166 9024 84194 9064
rect 87693 9027 87751 9033
rect 87693 9024 87705 9027
rect 84166 8996 87705 9024
rect 68741 8987 68799 8993
rect 87693 8993 87705 8996
rect 87739 8993 87751 9027
rect 87693 8987 87751 8993
rect 68278 8916 68284 8968
rect 68336 8956 68342 8968
rect 68557 8959 68615 8965
rect 68557 8956 68569 8959
rect 68336 8928 68569 8956
rect 68336 8916 68342 8928
rect 68557 8925 68569 8928
rect 68603 8925 68615 8959
rect 87414 8956 87420 8968
rect 87375 8928 87420 8956
rect 68557 8919 68615 8925
rect 87414 8916 87420 8928
rect 87472 8916 87478 8968
rect 86402 8888 86408 8900
rect 60706 8860 86408 8888
rect 52978 8851 53036 8857
rect 86402 8848 86408 8860
rect 86460 8848 86466 8900
rect 52181 8823 52239 8829
rect 52181 8789 52193 8823
rect 52227 8789 52239 8823
rect 52181 8783 52239 8789
rect 53098 8780 53104 8832
rect 53156 8820 53162 8832
rect 54113 8823 54171 8829
rect 54113 8820 54125 8823
rect 53156 8792 54125 8820
rect 53156 8780 53162 8792
rect 54113 8789 54125 8792
rect 54159 8789 54171 8823
rect 54113 8783 54171 8789
rect 68649 8823 68707 8829
rect 68649 8789 68661 8823
rect 68695 8820 68707 8823
rect 70762 8820 70768 8832
rect 68695 8792 70768 8820
rect 68695 8789 68707 8792
rect 68649 8783 68707 8789
rect 70762 8780 70768 8792
rect 70820 8780 70826 8832
rect 1104 8730 88872 8752
rect 1104 8678 22898 8730
rect 22950 8678 22962 8730
rect 23014 8678 23026 8730
rect 23078 8678 23090 8730
rect 23142 8678 23154 8730
rect 23206 8678 44846 8730
rect 44898 8678 44910 8730
rect 44962 8678 44974 8730
rect 45026 8678 45038 8730
rect 45090 8678 45102 8730
rect 45154 8678 66794 8730
rect 66846 8678 66858 8730
rect 66910 8678 66922 8730
rect 66974 8678 66986 8730
rect 67038 8678 67050 8730
rect 67102 8678 88872 8730
rect 1104 8656 88872 8678
rect 38013 8619 38071 8625
rect 38013 8585 38025 8619
rect 38059 8616 38071 8619
rect 40402 8616 40408 8628
rect 38059 8588 40408 8616
rect 38059 8585 38071 8588
rect 38013 8579 38071 8585
rect 40402 8576 40408 8588
rect 40460 8576 40466 8628
rect 42794 8616 42800 8628
rect 42755 8588 42800 8616
rect 42794 8576 42800 8588
rect 42852 8576 42858 8628
rect 43165 8619 43223 8625
rect 43165 8585 43177 8619
rect 43211 8616 43223 8619
rect 44082 8616 44088 8628
rect 43211 8588 44088 8616
rect 43211 8585 43223 8588
rect 43165 8579 43223 8585
rect 44082 8576 44088 8588
rect 44140 8576 44146 8628
rect 46106 8616 46112 8628
rect 46067 8588 46112 8616
rect 46106 8576 46112 8588
rect 46164 8576 46170 8628
rect 46477 8619 46535 8625
rect 46477 8585 46489 8619
rect 46523 8616 46535 8619
rect 47486 8616 47492 8628
rect 46523 8588 47492 8616
rect 46523 8585 46535 8588
rect 46477 8579 46535 8585
rect 47486 8576 47492 8588
rect 47544 8576 47550 8628
rect 48406 8576 48412 8628
rect 48464 8616 48470 8628
rect 49513 8619 49571 8625
rect 49513 8616 49525 8619
rect 48464 8588 49525 8616
rect 48464 8576 48470 8588
rect 49513 8585 49525 8588
rect 49559 8585 49571 8619
rect 50062 8616 50068 8628
rect 49513 8579 49571 8585
rect 49620 8588 50068 8616
rect 39022 8508 39028 8560
rect 39080 8548 39086 8560
rect 43257 8551 43315 8557
rect 43257 8548 43269 8551
rect 39080 8520 43269 8548
rect 39080 8508 39086 8520
rect 43257 8517 43269 8520
rect 43303 8517 43315 8551
rect 49620 8548 49648 8588
rect 50062 8576 50068 8588
rect 50120 8576 50126 8628
rect 50246 8616 50252 8628
rect 50207 8588 50252 8616
rect 50246 8576 50252 8588
rect 50304 8576 50310 8628
rect 52362 8576 52368 8628
rect 52420 8616 52426 8628
rect 52733 8619 52791 8625
rect 52733 8616 52745 8619
rect 52420 8588 52745 8616
rect 52420 8576 52426 8588
rect 52733 8585 52745 8588
rect 52779 8585 52791 8619
rect 53098 8616 53104 8628
rect 53059 8588 53104 8616
rect 52733 8579 52791 8585
rect 53098 8576 53104 8588
rect 53156 8576 53162 8628
rect 67542 8548 67548 8560
rect 43257 8511 43315 8517
rect 43364 8520 49648 8548
rect 49712 8520 67548 8548
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 27430 8480 27436 8492
rect 1719 8452 27436 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 27430 8440 27436 8452
rect 27488 8440 27494 8492
rect 38194 8480 38200 8492
rect 38155 8452 38200 8480
rect 38194 8440 38200 8452
rect 38252 8440 38258 8492
rect 41322 8440 41328 8492
rect 41380 8480 41386 8492
rect 41601 8483 41659 8489
rect 41601 8480 41613 8483
rect 41380 8452 41613 8480
rect 41380 8440 41386 8452
rect 41601 8449 41613 8452
rect 41647 8449 41659 8483
rect 41601 8443 41659 8449
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 33686 8372 33692 8424
rect 33744 8412 33750 8424
rect 41414 8412 41420 8424
rect 33744 8384 41420 8412
rect 33744 8372 33750 8384
rect 41414 8372 41420 8384
rect 41472 8412 41478 8424
rect 41472 8384 41565 8412
rect 41472 8372 41478 8384
rect 42058 8372 42064 8424
rect 42116 8412 42122 8424
rect 43364 8421 43392 8520
rect 43530 8440 43536 8492
rect 43588 8480 43594 8492
rect 48590 8480 48596 8492
rect 43588 8452 48596 8480
rect 43588 8440 43594 8452
rect 43349 8415 43407 8421
rect 43349 8412 43361 8415
rect 42116 8384 43361 8412
rect 42116 8372 42122 8384
rect 43349 8381 43361 8384
rect 43395 8381 43407 8415
rect 43349 8375 43407 8381
rect 45738 8372 45744 8424
rect 45796 8412 45802 8424
rect 46676 8421 46704 8452
rect 48590 8440 48596 8452
rect 48648 8440 48654 8492
rect 49712 8480 49740 8520
rect 67542 8508 67548 8520
rect 67600 8508 67606 8560
rect 49436 8452 49740 8480
rect 46569 8415 46627 8421
rect 46569 8412 46581 8415
rect 45796 8384 46581 8412
rect 45796 8372 45802 8384
rect 46569 8381 46581 8384
rect 46615 8381 46627 8415
rect 46569 8375 46627 8381
rect 46661 8415 46719 8421
rect 46661 8381 46673 8415
rect 46707 8381 46719 8415
rect 49436 8412 49464 8452
rect 49602 8412 49608 8424
rect 46661 8375 46719 8381
rect 47412 8384 49464 8412
rect 49563 8384 49608 8412
rect 39298 8304 39304 8356
rect 39356 8344 39362 8356
rect 47412 8344 47440 8384
rect 49602 8372 49608 8384
rect 49660 8372 49666 8424
rect 49712 8421 49740 8452
rect 50433 8483 50491 8489
rect 50433 8449 50445 8483
rect 50479 8449 50491 8483
rect 50433 8443 50491 8449
rect 53193 8483 53251 8489
rect 53193 8449 53205 8483
rect 53239 8480 53251 8483
rect 55582 8480 55588 8492
rect 53239 8452 55588 8480
rect 53239 8449 53251 8452
rect 53193 8443 53251 8449
rect 49697 8415 49755 8421
rect 49697 8381 49709 8415
rect 49743 8381 49755 8415
rect 49697 8375 49755 8381
rect 39356 8316 47440 8344
rect 49145 8347 49203 8353
rect 39356 8304 39362 8316
rect 49145 8313 49157 8347
rect 49191 8344 49203 8347
rect 50448 8344 50476 8443
rect 55582 8440 55588 8452
rect 55640 8440 55646 8492
rect 88242 8480 88248 8492
rect 88203 8452 88248 8480
rect 88242 8440 88248 8452
rect 88300 8440 88306 8492
rect 53285 8415 53343 8421
rect 53285 8381 53297 8415
rect 53331 8381 53343 8415
rect 53285 8375 53343 8381
rect 49191 8316 50476 8344
rect 49191 8313 49203 8316
rect 49145 8307 49203 8313
rect 50798 8304 50804 8356
rect 50856 8344 50862 8356
rect 53300 8344 53328 8375
rect 50856 8316 53328 8344
rect 50856 8304 50862 8316
rect 82814 8304 82820 8356
rect 82872 8344 82878 8356
rect 88061 8347 88119 8353
rect 88061 8344 88073 8347
rect 82872 8316 88073 8344
rect 82872 8304 82878 8316
rect 88061 8313 88073 8316
rect 88107 8313 88119 8347
rect 88061 8307 88119 8313
rect 41785 8279 41843 8285
rect 41785 8245 41797 8279
rect 41831 8276 41843 8279
rect 41874 8276 41880 8288
rect 41831 8248 41880 8276
rect 41831 8245 41843 8248
rect 41785 8239 41843 8245
rect 41874 8236 41880 8248
rect 41932 8236 41938 8288
rect 1104 8186 88872 8208
rect 1104 8134 11924 8186
rect 11976 8134 11988 8186
rect 12040 8134 12052 8186
rect 12104 8134 12116 8186
rect 12168 8134 12180 8186
rect 12232 8134 33872 8186
rect 33924 8134 33936 8186
rect 33988 8134 34000 8186
rect 34052 8134 34064 8186
rect 34116 8134 34128 8186
rect 34180 8134 55820 8186
rect 55872 8134 55884 8186
rect 55936 8134 55948 8186
rect 56000 8134 56012 8186
rect 56064 8134 56076 8186
rect 56128 8134 77768 8186
rect 77820 8134 77832 8186
rect 77884 8134 77896 8186
rect 77948 8134 77960 8186
rect 78012 8134 78024 8186
rect 78076 8134 88872 8186
rect 1104 8112 88872 8134
rect 46474 8072 46480 8084
rect 46435 8044 46480 8072
rect 46474 8032 46480 8044
rect 46532 8032 46538 8084
rect 41874 7868 41880 7880
rect 41835 7840 41880 7868
rect 41874 7828 41880 7840
rect 41932 7828 41938 7880
rect 46661 7871 46719 7877
rect 46661 7837 46673 7871
rect 46707 7868 46719 7871
rect 48130 7868 48136 7880
rect 46707 7840 48136 7868
rect 46707 7837 46719 7840
rect 46661 7831 46719 7837
rect 48130 7828 48136 7840
rect 48188 7828 48194 7880
rect 64322 7828 64328 7880
rect 64380 7868 64386 7880
rect 87693 7871 87751 7877
rect 87693 7868 87705 7871
rect 64380 7840 87705 7868
rect 64380 7828 64386 7840
rect 87693 7837 87705 7840
rect 87739 7868 87751 7871
rect 88245 7871 88303 7877
rect 88245 7868 88257 7871
rect 87739 7840 88257 7868
rect 87739 7837 87751 7840
rect 87693 7831 87751 7837
rect 88245 7837 88257 7840
rect 88291 7837 88303 7871
rect 88245 7831 88303 7837
rect 20806 7760 20812 7812
rect 20864 7800 20870 7812
rect 58434 7800 58440 7812
rect 20864 7772 58440 7800
rect 20864 7760 20870 7772
rect 58434 7760 58440 7772
rect 58492 7760 58498 7812
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 34422 7732 34428 7744
rect 1728 7704 34428 7732
rect 1728 7692 1734 7704
rect 34422 7692 34428 7704
rect 34480 7692 34486 7744
rect 41693 7735 41751 7741
rect 41693 7701 41705 7735
rect 41739 7732 41751 7735
rect 41966 7732 41972 7744
rect 41739 7704 41972 7732
rect 41739 7701 41751 7704
rect 41693 7695 41751 7701
rect 41966 7692 41972 7704
rect 42024 7692 42030 7744
rect 88058 7732 88064 7744
rect 88019 7704 88064 7732
rect 88058 7692 88064 7704
rect 88116 7692 88122 7744
rect 1104 7642 88872 7664
rect 1104 7590 22898 7642
rect 22950 7590 22962 7642
rect 23014 7590 23026 7642
rect 23078 7590 23090 7642
rect 23142 7590 23154 7642
rect 23206 7590 44846 7642
rect 44898 7590 44910 7642
rect 44962 7590 44974 7642
rect 45026 7590 45038 7642
rect 45090 7590 45102 7642
rect 45154 7590 66794 7642
rect 66846 7590 66858 7642
rect 66910 7590 66922 7642
rect 66974 7590 66986 7642
rect 67038 7590 67050 7642
rect 67102 7590 88872 7642
rect 1104 7568 88872 7590
rect 40310 7528 40316 7540
rect 40271 7500 40316 7528
rect 40310 7488 40316 7500
rect 40368 7488 40374 7540
rect 38654 7420 38660 7472
rect 38712 7460 38718 7472
rect 39025 7463 39083 7469
rect 39025 7460 39037 7463
rect 38712 7432 39037 7460
rect 38712 7420 38718 7432
rect 39025 7429 39037 7432
rect 39071 7429 39083 7463
rect 39025 7423 39083 7429
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 18598 7392 18604 7404
rect 1627 7364 18604 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 88058 7392 88064 7404
rect 88019 7364 88064 7392
rect 88058 7352 88064 7364
rect 88116 7352 88122 7404
rect 36722 7216 36728 7268
rect 36780 7256 36786 7268
rect 88245 7259 88303 7265
rect 88245 7256 88257 7259
rect 36780 7228 88257 7256
rect 36780 7216 36786 7228
rect 88245 7225 88257 7228
rect 88291 7225 88303 7259
rect 88245 7219 88303 7225
rect 1394 7188 1400 7200
rect 1355 7160 1400 7188
rect 1394 7148 1400 7160
rect 1452 7148 1458 7200
rect 1104 7098 88872 7120
rect 1104 7046 11924 7098
rect 11976 7046 11988 7098
rect 12040 7046 12052 7098
rect 12104 7046 12116 7098
rect 12168 7046 12180 7098
rect 12232 7046 33872 7098
rect 33924 7046 33936 7098
rect 33988 7046 34000 7098
rect 34052 7046 34064 7098
rect 34116 7046 34128 7098
rect 34180 7046 55820 7098
rect 55872 7046 55884 7098
rect 55936 7046 55948 7098
rect 56000 7046 56012 7098
rect 56064 7046 56076 7098
rect 56128 7046 77768 7098
rect 77820 7046 77832 7098
rect 77884 7046 77896 7098
rect 77948 7046 77960 7098
rect 78012 7046 78024 7098
rect 78076 7046 88872 7098
rect 1104 7024 88872 7046
rect 49878 6808 49884 6860
rect 49936 6848 49942 6860
rect 53190 6848 53196 6860
rect 49936 6820 53196 6848
rect 49936 6808 49942 6820
rect 53190 6808 53196 6820
rect 53248 6808 53254 6860
rect 26145 6783 26203 6789
rect 26145 6749 26157 6783
rect 26191 6749 26203 6783
rect 26418 6780 26424 6792
rect 26379 6752 26424 6780
rect 26145 6743 26203 6749
rect 26160 6712 26188 6743
rect 26418 6740 26424 6752
rect 26476 6740 26482 6792
rect 39025 6783 39083 6789
rect 39025 6780 39037 6783
rect 31726 6752 39037 6780
rect 31386 6712 31392 6724
rect 26160 6684 31392 6712
rect 31386 6672 31392 6684
rect 31444 6712 31450 6724
rect 31726 6712 31754 6752
rect 39025 6749 39037 6752
rect 39071 6749 39083 6783
rect 39025 6743 39083 6749
rect 39114 6740 39120 6792
rect 39172 6780 39178 6792
rect 39301 6783 39359 6789
rect 39301 6780 39313 6783
rect 39172 6752 39313 6780
rect 39172 6740 39178 6752
rect 39301 6749 39313 6752
rect 39347 6749 39359 6783
rect 39301 6743 39359 6749
rect 56781 6783 56839 6789
rect 56781 6749 56793 6783
rect 56827 6780 56839 6783
rect 56962 6780 56968 6792
rect 56827 6752 56968 6780
rect 56827 6749 56839 6752
rect 56781 6743 56839 6749
rect 56962 6740 56968 6752
rect 57020 6740 57026 6792
rect 31444 6684 31754 6712
rect 38841 6715 38899 6721
rect 31444 6672 31450 6684
rect 38841 6681 38853 6715
rect 38887 6712 38899 6715
rect 39942 6712 39948 6724
rect 38887 6684 39948 6712
rect 38887 6681 38899 6684
rect 38841 6675 38899 6681
rect 39942 6672 39948 6684
rect 40000 6672 40006 6724
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 20772 6616 25973 6644
rect 20772 6604 20778 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 26329 6647 26387 6653
rect 26329 6613 26341 6647
rect 26375 6644 26387 6647
rect 35250 6644 35256 6656
rect 26375 6616 35256 6644
rect 26375 6613 26387 6616
rect 26329 6607 26387 6613
rect 35250 6604 35256 6616
rect 35308 6644 35314 6656
rect 39209 6647 39267 6653
rect 39209 6644 39221 6647
rect 35308 6616 39221 6644
rect 35308 6604 35314 6616
rect 39209 6613 39221 6616
rect 39255 6613 39267 6647
rect 39209 6607 39267 6613
rect 56042 6604 56048 6656
rect 56100 6644 56106 6656
rect 56597 6647 56655 6653
rect 56597 6644 56609 6647
rect 56100 6616 56609 6644
rect 56100 6604 56106 6616
rect 56597 6613 56609 6616
rect 56643 6613 56655 6647
rect 56597 6607 56655 6613
rect 1104 6554 88872 6576
rect 1104 6502 22898 6554
rect 22950 6502 22962 6554
rect 23014 6502 23026 6554
rect 23078 6502 23090 6554
rect 23142 6502 23154 6554
rect 23206 6502 44846 6554
rect 44898 6502 44910 6554
rect 44962 6502 44974 6554
rect 45026 6502 45038 6554
rect 45090 6502 45102 6554
rect 45154 6502 66794 6554
rect 66846 6502 66858 6554
rect 66910 6502 66922 6554
rect 66974 6502 66986 6554
rect 67038 6502 67050 6554
rect 67102 6502 88872 6554
rect 1104 6480 88872 6502
rect 48498 6400 48504 6452
rect 48556 6440 48562 6452
rect 57149 6443 57207 6449
rect 57149 6440 57161 6443
rect 48556 6412 57161 6440
rect 48556 6400 48562 6412
rect 57149 6409 57161 6412
rect 57195 6440 57207 6443
rect 57330 6440 57336 6452
rect 57195 6412 57336 6440
rect 57195 6409 57207 6412
rect 57149 6403 57207 6409
rect 57330 6400 57336 6412
rect 57388 6400 57394 6452
rect 1762 6304 1768 6316
rect 1723 6276 1768 6304
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 55306 6264 55312 6316
rect 55364 6304 55370 6316
rect 55769 6307 55827 6313
rect 55769 6304 55781 6307
rect 55364 6276 55781 6304
rect 55364 6264 55370 6276
rect 55769 6273 55781 6276
rect 55815 6273 55827 6307
rect 56042 6304 56048 6316
rect 56003 6276 56048 6304
rect 55769 6267 55827 6273
rect 56042 6264 56048 6276
rect 56100 6264 56106 6316
rect 87414 6236 87420 6248
rect 87375 6208 87420 6236
rect 87414 6196 87420 6208
rect 87472 6196 87478 6248
rect 87690 6236 87696 6248
rect 87651 6208 87696 6236
rect 87690 6196 87696 6208
rect 87748 6196 87754 6248
rect 31570 6128 31576 6180
rect 31628 6168 31634 6180
rect 34790 6168 34796 6180
rect 31628 6140 34796 6168
rect 31628 6128 31634 6140
rect 34790 6128 34796 6140
rect 34848 6128 34854 6180
rect 63954 6168 63960 6180
rect 56704 6140 63960 6168
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 56704 6100 56732 6140
rect 63954 6128 63960 6140
rect 64012 6128 64018 6180
rect 2087 6072 56732 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 1104 6010 88872 6032
rect 1104 5958 11924 6010
rect 11976 5958 11988 6010
rect 12040 5958 12052 6010
rect 12104 5958 12116 6010
rect 12168 5958 12180 6010
rect 12232 5958 33872 6010
rect 33924 5958 33936 6010
rect 33988 5958 34000 6010
rect 34052 5958 34064 6010
rect 34116 5958 34128 6010
rect 34180 5958 55820 6010
rect 55872 5958 55884 6010
rect 55936 5958 55948 6010
rect 56000 5958 56012 6010
rect 56064 5958 56076 6010
rect 56128 5958 77768 6010
rect 77820 5958 77832 6010
rect 77884 5958 77896 6010
rect 77948 5958 77960 6010
rect 78012 5958 78024 6010
rect 78076 5958 88872 6010
rect 1104 5936 88872 5958
rect 56962 5896 56968 5908
rect 22066 5868 31754 5896
rect 56923 5868 56968 5896
rect 20990 5720 20996 5772
rect 21048 5760 21054 5772
rect 22066 5760 22094 5868
rect 21048 5732 22094 5760
rect 21048 5720 21054 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 1627 5664 2912 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 1394 5556 1400 5568
rect 1355 5528 1400 5556
rect 1394 5516 1400 5528
rect 1452 5516 1458 5568
rect 2884 5565 2912 5664
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 3694 5692 3700 5704
rect 3108 5664 3700 5692
rect 3108 5652 3114 5664
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 25130 5692 25136 5704
rect 25091 5664 25136 5692
rect 25130 5652 25136 5664
rect 25188 5652 25194 5704
rect 25685 5695 25743 5701
rect 25685 5661 25697 5695
rect 25731 5692 25743 5695
rect 25774 5692 25780 5704
rect 25731 5664 25780 5692
rect 25731 5661 25743 5664
rect 25685 5655 25743 5661
rect 25774 5652 25780 5664
rect 25832 5692 25838 5704
rect 25832 5664 26188 5692
rect 25832 5652 25838 5664
rect 26160 5636 26188 5664
rect 25930 5627 25988 5633
rect 25930 5624 25942 5627
rect 24964 5596 25942 5624
rect 24964 5565 24992 5596
rect 25930 5593 25942 5596
rect 25976 5593 25988 5627
rect 25930 5587 25988 5593
rect 26142 5584 26148 5636
rect 26200 5584 26206 5636
rect 2869 5559 2927 5565
rect 2869 5525 2881 5559
rect 2915 5525 2927 5559
rect 2869 5519 2927 5525
rect 24949 5559 25007 5565
rect 24949 5525 24961 5559
rect 24995 5525 25007 5559
rect 24949 5519 25007 5525
rect 26418 5516 26424 5568
rect 26476 5556 26482 5568
rect 27065 5559 27123 5565
rect 27065 5556 27077 5559
rect 26476 5528 27077 5556
rect 26476 5516 26482 5528
rect 27065 5525 27077 5528
rect 27111 5525 27123 5559
rect 31726 5556 31754 5868
rect 56962 5856 56968 5868
rect 57020 5856 57026 5908
rect 56689 5763 56747 5769
rect 56689 5729 56701 5763
rect 56735 5760 56747 5763
rect 57609 5763 57667 5769
rect 57609 5760 57621 5763
rect 56735 5732 57621 5760
rect 56735 5729 56747 5732
rect 56689 5723 56747 5729
rect 57609 5729 57621 5732
rect 57655 5760 57667 5763
rect 57698 5760 57704 5772
rect 57655 5732 57704 5760
rect 57655 5729 57667 5732
rect 57609 5723 57667 5729
rect 57698 5720 57704 5732
rect 57756 5720 57762 5772
rect 57330 5692 57336 5704
rect 57291 5664 57336 5692
rect 57330 5652 57336 5664
rect 57388 5652 57394 5704
rect 57425 5695 57483 5701
rect 57425 5661 57437 5695
rect 57471 5692 57483 5695
rect 87966 5692 87972 5704
rect 57471 5664 70394 5692
rect 87927 5664 87972 5692
rect 57471 5661 57483 5664
rect 57425 5655 57483 5661
rect 70366 5624 70394 5664
rect 87966 5652 87972 5664
rect 88024 5652 88030 5704
rect 87690 5624 87696 5636
rect 41386 5596 60734 5624
rect 70366 5596 87696 5624
rect 41386 5556 41414 5596
rect 31726 5528 41414 5556
rect 60706 5556 60734 5596
rect 87690 5584 87696 5596
rect 87748 5584 87754 5636
rect 88153 5559 88211 5565
rect 88153 5556 88165 5559
rect 60706 5528 88165 5556
rect 27065 5519 27123 5525
rect 88153 5525 88165 5528
rect 88199 5525 88211 5559
rect 88153 5519 88211 5525
rect 1104 5466 88872 5488
rect 1104 5414 22898 5466
rect 22950 5414 22962 5466
rect 23014 5414 23026 5466
rect 23078 5414 23090 5466
rect 23142 5414 23154 5466
rect 23206 5414 44846 5466
rect 44898 5414 44910 5466
rect 44962 5414 44974 5466
rect 45026 5414 45038 5466
rect 45090 5414 45102 5466
rect 45154 5414 66794 5466
rect 66846 5414 66858 5466
rect 66910 5414 66922 5466
rect 66974 5414 66986 5466
rect 67038 5414 67050 5466
rect 67102 5414 88872 5466
rect 1104 5392 88872 5414
rect 24213 5355 24271 5361
rect 24213 5321 24225 5355
rect 24259 5352 24271 5355
rect 25130 5352 25136 5364
rect 24259 5324 25136 5352
rect 24259 5321 24271 5324
rect 24213 5315 24271 5321
rect 25130 5312 25136 5324
rect 25188 5312 25194 5364
rect 27709 5355 27767 5361
rect 27709 5321 27721 5355
rect 27755 5352 27767 5355
rect 29362 5352 29368 5364
rect 27755 5324 29368 5352
rect 27755 5321 27767 5324
rect 27709 5315 27767 5321
rect 24581 5287 24639 5293
rect 24581 5253 24593 5287
rect 24627 5284 24639 5287
rect 26418 5284 26424 5296
rect 24627 5256 26424 5284
rect 24627 5253 24639 5256
rect 24581 5247 24639 5253
rect 26418 5244 26424 5256
rect 26476 5244 26482 5296
rect 23658 5176 23664 5228
rect 23716 5216 23722 5228
rect 26436 5216 26464 5244
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 23716 5188 24808 5216
rect 26436 5188 27169 5216
rect 23716 5176 23722 5188
rect 24780 5160 24808 5188
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 24673 5151 24731 5157
rect 24673 5148 24685 5151
rect 17276 5120 24685 5148
rect 17276 5108 17282 5120
rect 24673 5117 24685 5120
rect 24719 5117 24731 5151
rect 24673 5111 24731 5117
rect 24762 5108 24768 5160
rect 24820 5148 24826 5160
rect 26973 5151 27031 5157
rect 24820 5120 24913 5148
rect 24820 5108 24826 5120
rect 26973 5117 26985 5151
rect 27019 5148 27031 5151
rect 27724 5148 27752 5315
rect 29362 5312 29368 5324
rect 29420 5312 29426 5364
rect 29454 5312 29460 5364
rect 29512 5352 29518 5364
rect 30009 5355 30067 5361
rect 30009 5352 30021 5355
rect 29512 5324 30021 5352
rect 29512 5312 29518 5324
rect 30009 5321 30021 5324
rect 30055 5321 30067 5355
rect 30009 5315 30067 5321
rect 29917 5287 29975 5293
rect 29917 5253 29929 5287
rect 29963 5284 29975 5287
rect 30650 5284 30656 5296
rect 29963 5256 30656 5284
rect 29963 5253 29975 5256
rect 29917 5247 29975 5253
rect 30650 5244 30656 5256
rect 30708 5244 30714 5296
rect 44542 5176 44548 5228
rect 44600 5216 44606 5228
rect 87693 5219 87751 5225
rect 87693 5216 87705 5219
rect 44600 5188 87705 5216
rect 44600 5176 44606 5188
rect 87693 5185 87705 5188
rect 87739 5216 87751 5219
rect 88245 5219 88303 5225
rect 88245 5216 88257 5219
rect 87739 5188 88257 5216
rect 87739 5185 87751 5188
rect 87693 5179 87751 5185
rect 88245 5185 88257 5188
rect 88291 5185 88303 5219
rect 88245 5179 88303 5185
rect 27019 5120 27752 5148
rect 27019 5117 27031 5120
rect 26973 5111 27031 5117
rect 26694 4972 26700 5024
rect 26752 5012 26758 5024
rect 27341 5015 27399 5021
rect 27341 5012 27353 5015
rect 26752 4984 27353 5012
rect 26752 4972 26758 4984
rect 27341 4981 27353 4984
rect 27387 4981 27399 5015
rect 27341 4975 27399 4981
rect 70670 4972 70676 5024
rect 70728 5012 70734 5024
rect 71222 5012 71228 5024
rect 70728 4984 71228 5012
rect 70728 4972 70734 4984
rect 71222 4972 71228 4984
rect 71280 4972 71286 5024
rect 88058 5012 88064 5024
rect 88019 4984 88064 5012
rect 88058 4972 88064 4984
rect 88116 4972 88122 5024
rect 1104 4922 88872 4944
rect 1104 4870 11924 4922
rect 11976 4870 11988 4922
rect 12040 4870 12052 4922
rect 12104 4870 12116 4922
rect 12168 4870 12180 4922
rect 12232 4870 33872 4922
rect 33924 4870 33936 4922
rect 33988 4870 34000 4922
rect 34052 4870 34064 4922
rect 34116 4870 34128 4922
rect 34180 4870 55820 4922
rect 55872 4870 55884 4922
rect 55936 4870 55948 4922
rect 56000 4870 56012 4922
rect 56064 4870 56076 4922
rect 56128 4870 77768 4922
rect 77820 4870 77832 4922
rect 77884 4870 77896 4922
rect 77948 4870 77960 4922
rect 78012 4870 78024 4922
rect 78076 4870 88872 4922
rect 1104 4848 88872 4870
rect 31846 4768 31852 4820
rect 31904 4808 31910 4820
rect 33045 4811 33103 4817
rect 33045 4808 33057 4811
rect 31904 4780 33057 4808
rect 31904 4768 31910 4780
rect 33045 4777 33057 4780
rect 33091 4808 33103 4811
rect 41230 4808 41236 4820
rect 33091 4780 41236 4808
rect 33091 4777 33103 4780
rect 33045 4771 33103 4777
rect 41230 4768 41236 4780
rect 41288 4808 41294 4820
rect 50706 4808 50712 4820
rect 41288 4780 50712 4808
rect 41288 4768 41294 4780
rect 50706 4768 50712 4780
rect 50764 4808 50770 4820
rect 51442 4808 51448 4820
rect 50764 4780 51448 4808
rect 50764 4768 50770 4780
rect 51442 4768 51448 4780
rect 51500 4768 51506 4820
rect 63218 4768 63224 4820
rect 63276 4808 63282 4820
rect 83826 4808 83832 4820
rect 63276 4780 83832 4808
rect 63276 4768 63282 4780
rect 83826 4768 83832 4780
rect 83884 4768 83890 4820
rect 24397 4743 24455 4749
rect 24397 4709 24409 4743
rect 24443 4709 24455 4743
rect 24397 4703 24455 4709
rect 25501 4743 25559 4749
rect 25501 4709 25513 4743
rect 25547 4709 25559 4743
rect 25501 4703 25559 4709
rect 1578 4604 1584 4616
rect 1539 4576 1584 4604
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 24412 4604 24440 4703
rect 24762 4632 24768 4684
rect 24820 4672 24826 4684
rect 24949 4675 25007 4681
rect 24949 4672 24961 4675
rect 24820 4644 24961 4672
rect 24820 4632 24826 4644
rect 24949 4641 24961 4644
rect 24995 4641 25007 4675
rect 25516 4672 25544 4703
rect 37918 4700 37924 4752
rect 37976 4740 37982 4752
rect 87693 4743 87751 4749
rect 87693 4740 87705 4743
rect 37976 4712 87705 4740
rect 37976 4700 37982 4712
rect 87693 4709 87705 4712
rect 87739 4709 87751 4743
rect 87693 4703 87751 4709
rect 26421 4675 26479 4681
rect 26421 4672 26433 4675
rect 25516 4644 26433 4672
rect 24949 4635 25007 4641
rect 26421 4641 26433 4644
rect 26467 4641 26479 4675
rect 26421 4635 26479 4641
rect 29362 4632 29368 4684
rect 29420 4672 29426 4684
rect 55309 4675 55367 4681
rect 55309 4672 55321 4675
rect 29420 4644 55321 4672
rect 29420 4632 29426 4644
rect 55309 4641 55321 4644
rect 55355 4672 55367 4675
rect 56045 4675 56103 4681
rect 56045 4672 56057 4675
rect 55355 4644 56057 4672
rect 55355 4641 55367 4644
rect 55309 4635 55367 4641
rect 56045 4641 56057 4644
rect 56091 4672 56103 4675
rect 56091 4644 60734 4672
rect 56091 4641 56103 4644
rect 56045 4635 56103 4641
rect 25685 4607 25743 4613
rect 25685 4604 25697 4607
rect 24412 4576 25697 4604
rect 25685 4573 25697 4576
rect 25731 4573 25743 4607
rect 26142 4604 26148 4616
rect 26103 4576 26148 4604
rect 25685 4567 25743 4573
rect 26142 4564 26148 4576
rect 26200 4564 26206 4616
rect 55493 4607 55551 4613
rect 55493 4573 55505 4607
rect 55539 4604 55551 4607
rect 57330 4604 57336 4616
rect 55539 4576 57336 4604
rect 55539 4573 55551 4576
rect 55493 4567 55551 4573
rect 57330 4564 57336 4576
rect 57388 4564 57394 4616
rect 60706 4604 60734 4644
rect 71130 4604 71136 4616
rect 60706 4576 71136 4604
rect 71130 4564 71136 4576
rect 71188 4564 71194 4616
rect 87708 4604 87736 4703
rect 88245 4607 88303 4613
rect 88245 4604 88257 4607
rect 87708 4576 88257 4604
rect 88245 4573 88257 4576
rect 88291 4573 88303 4607
rect 88245 4567 88303 4573
rect 17218 4536 17224 4548
rect 6886 4508 17224 4536
rect 1397 4471 1455 4477
rect 1397 4437 1409 4471
rect 1443 4468 1455 4471
rect 6886 4468 6914 4508
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 24857 4539 24915 4545
rect 24857 4536 24869 4539
rect 22066 4508 24869 4536
rect 1443 4440 6914 4468
rect 1443 4437 1455 4440
rect 1397 4431 1455 4437
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 22066 4468 22094 4508
rect 24857 4505 24869 4508
rect 24903 4505 24915 4539
rect 24857 4499 24915 4505
rect 32769 4539 32827 4545
rect 32769 4505 32781 4539
rect 32815 4536 32827 4539
rect 32950 4536 32956 4548
rect 32815 4508 32956 4536
rect 32815 4505 32827 4508
rect 32769 4499 32827 4505
rect 32950 4496 32956 4508
rect 33008 4496 33014 4548
rect 33594 4536 33600 4548
rect 33507 4508 33600 4536
rect 33594 4496 33600 4508
rect 33652 4536 33658 4548
rect 59446 4536 59452 4548
rect 33652 4508 59452 4536
rect 33652 4496 33658 4508
rect 59446 4496 59452 4508
rect 59504 4496 59510 4548
rect 18012 4440 22094 4468
rect 18012 4428 18018 4440
rect 22646 4428 22652 4480
rect 22704 4468 22710 4480
rect 24765 4471 24823 4477
rect 24765 4468 24777 4471
rect 22704 4440 24777 4468
rect 22704 4428 22710 4440
rect 24765 4437 24777 4440
rect 24811 4468 24823 4471
rect 27522 4468 27528 4480
rect 24811 4440 27528 4468
rect 24811 4437 24823 4440
rect 24765 4431 24823 4437
rect 27522 4428 27528 4440
rect 27580 4428 27586 4480
rect 27706 4428 27712 4480
rect 27764 4468 27770 4480
rect 28902 4468 28908 4480
rect 27764 4440 28908 4468
rect 27764 4428 27770 4440
rect 28902 4428 28908 4440
rect 28960 4468 28966 4480
rect 33689 4471 33747 4477
rect 33689 4468 33701 4471
rect 28960 4440 33701 4468
rect 28960 4428 28966 4440
rect 33689 4437 33701 4440
rect 33735 4437 33747 4471
rect 33689 4431 33747 4437
rect 38838 4428 38844 4480
rect 38896 4468 38902 4480
rect 46290 4468 46296 4480
rect 38896 4440 46296 4468
rect 38896 4428 38902 4440
rect 46290 4428 46296 4440
rect 46348 4428 46354 4480
rect 49234 4428 49240 4480
rect 49292 4468 49298 4480
rect 53098 4468 53104 4480
rect 49292 4440 53104 4468
rect 49292 4428 49298 4440
rect 53098 4428 53104 4440
rect 53156 4428 53162 4480
rect 55674 4468 55680 4480
rect 55635 4440 55680 4468
rect 55674 4428 55680 4440
rect 55732 4428 55738 4480
rect 88058 4468 88064 4480
rect 88019 4440 88064 4468
rect 88058 4428 88064 4440
rect 88116 4428 88122 4480
rect 1104 4378 88872 4400
rect 1104 4326 22898 4378
rect 22950 4326 22962 4378
rect 23014 4326 23026 4378
rect 23078 4326 23090 4378
rect 23142 4326 23154 4378
rect 23206 4326 44846 4378
rect 44898 4326 44910 4378
rect 44962 4326 44974 4378
rect 45026 4326 45038 4378
rect 45090 4326 45102 4378
rect 45154 4326 66794 4378
rect 66846 4326 66858 4378
rect 66910 4326 66922 4378
rect 66974 4326 66986 4378
rect 67038 4326 67050 4378
rect 67102 4326 88872 4378
rect 1104 4304 88872 4326
rect 27522 4224 27528 4276
rect 27580 4264 27586 4276
rect 49418 4264 49424 4276
rect 27580 4236 41414 4264
rect 49379 4236 49424 4264
rect 27580 4224 27586 4236
rect 30650 4156 30656 4208
rect 30708 4196 30714 4208
rect 31202 4196 31208 4208
rect 30708 4168 31208 4196
rect 30708 4156 30714 4168
rect 31202 4156 31208 4168
rect 31260 4196 31266 4208
rect 33594 4196 33600 4208
rect 31260 4168 33600 4196
rect 31260 4156 31266 4168
rect 33594 4156 33600 4168
rect 33652 4156 33658 4208
rect 41386 4196 41414 4236
rect 49418 4224 49424 4236
rect 49476 4224 49482 4276
rect 53098 4224 53104 4276
rect 53156 4264 53162 4276
rect 53156 4236 70900 4264
rect 53156 4224 53162 4236
rect 49234 4196 49240 4208
rect 41386 4168 49240 4196
rect 49234 4156 49240 4168
rect 49292 4156 49298 4208
rect 51442 4156 51448 4208
rect 51500 4196 51506 4208
rect 51629 4199 51687 4205
rect 51500 4168 51580 4196
rect 51500 4156 51506 4168
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 2133 4131 2191 4137
rect 2133 4128 2145 4131
rect 1719 4100 2145 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2133 4097 2145 4100
rect 2179 4128 2191 4131
rect 2179 4100 6914 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3992 2007 3995
rect 2774 3992 2780 4004
rect 1995 3964 2780 3992
rect 1995 3961 2007 3964
rect 1949 3955 2007 3961
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 2409 3927 2467 3933
rect 2409 3893 2421 3927
rect 2455 3924 2467 3927
rect 2958 3924 2964 3936
rect 2455 3896 2964 3924
rect 2455 3893 2467 3896
rect 2409 3887 2467 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 6886 3924 6914 4100
rect 25406 4088 25412 4140
rect 25464 4128 25470 4140
rect 44358 4128 44364 4140
rect 25464 4100 44364 4128
rect 25464 4088 25470 4100
rect 44358 4088 44364 4100
rect 44416 4088 44422 4140
rect 49605 4131 49663 4137
rect 49605 4097 49617 4131
rect 49651 4128 49663 4131
rect 49970 4128 49976 4140
rect 49651 4100 49976 4128
rect 49651 4097 49663 4100
rect 49605 4091 49663 4097
rect 49970 4088 49976 4100
rect 50028 4088 50034 4140
rect 19150 4020 19156 4072
rect 19208 4060 19214 4072
rect 45370 4060 45376 4072
rect 19208 4032 45376 4060
rect 19208 4020 19214 4032
rect 45370 4020 45376 4032
rect 45428 4020 45434 4072
rect 51442 4060 51448 4072
rect 46124 4032 51448 4060
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 28994 3992 29000 4004
rect 7156 3964 29000 3992
rect 7156 3952 7162 3964
rect 28994 3952 29000 3964
rect 29052 3952 29058 4004
rect 29178 3952 29184 4004
rect 29236 3992 29242 4004
rect 36538 3992 36544 4004
rect 29236 3964 36544 3992
rect 29236 3952 29242 3964
rect 36538 3952 36544 3964
rect 36596 3952 36602 4004
rect 38102 3952 38108 4004
rect 38160 3992 38166 4004
rect 43438 3992 43444 4004
rect 38160 3964 43444 3992
rect 38160 3952 38166 3964
rect 43438 3952 43444 3964
rect 43496 3952 43502 4004
rect 46124 3924 46152 4032
rect 51442 4020 51448 4032
rect 51500 4020 51506 4072
rect 51552 4060 51580 4168
rect 51629 4165 51641 4199
rect 51675 4196 51687 4199
rect 51810 4196 51816 4208
rect 51675 4168 51816 4196
rect 51675 4165 51687 4168
rect 51629 4159 51687 4165
rect 51810 4156 51816 4168
rect 51868 4156 51874 4208
rect 59446 4156 59452 4208
rect 59504 4196 59510 4208
rect 59541 4199 59599 4205
rect 59541 4196 59553 4199
rect 59504 4168 59553 4196
rect 59504 4156 59510 4168
rect 59541 4165 59553 4168
rect 59587 4196 59599 4199
rect 70670 4196 70676 4208
rect 59587 4168 70676 4196
rect 59587 4165 59599 4168
rect 59541 4159 59599 4165
rect 70670 4156 70676 4168
rect 70728 4156 70734 4208
rect 70872 4205 70900 4236
rect 70857 4199 70915 4205
rect 70857 4165 70869 4199
rect 70903 4196 70915 4199
rect 70903 4168 71360 4196
rect 70903 4165 70915 4168
rect 70857 4159 70915 4165
rect 51721 4131 51779 4137
rect 51721 4097 51733 4131
rect 51767 4128 51779 4131
rect 54018 4128 54024 4140
rect 51767 4100 54024 4128
rect 51767 4097 51779 4100
rect 51721 4091 51779 4097
rect 54018 4088 54024 4100
rect 54076 4088 54082 4140
rect 63586 4128 63592 4140
rect 60706 4100 63592 4128
rect 51813 4063 51871 4069
rect 51813 4060 51825 4063
rect 51552 4032 51825 4060
rect 51813 4029 51825 4032
rect 51859 4029 51871 4063
rect 51813 4023 51871 4029
rect 51902 4020 51908 4072
rect 51960 4060 51966 4072
rect 60706 4060 60734 4100
rect 63586 4088 63592 4100
rect 63644 4128 63650 4140
rect 64046 4128 64052 4140
rect 63644 4100 64052 4128
rect 63644 4088 63650 4100
rect 64046 4088 64052 4100
rect 64104 4088 64110 4140
rect 71332 4137 71360 4168
rect 86788 4168 87828 4196
rect 71317 4131 71375 4137
rect 70366 4100 71268 4128
rect 70366 4060 70394 4100
rect 71130 4060 71136 4072
rect 51960 4032 60734 4060
rect 63696 4032 70394 4060
rect 71091 4032 71136 4060
rect 51960 4020 51966 4032
rect 46474 3952 46480 4004
rect 46532 3992 46538 4004
rect 63696 3992 63724 4032
rect 71130 4020 71136 4032
rect 71188 4020 71194 4072
rect 71240 4060 71268 4100
rect 71317 4097 71329 4131
rect 71363 4128 71375 4131
rect 86788 4128 86816 4168
rect 71363 4100 86816 4128
rect 71363 4097 71375 4100
rect 71317 4091 71375 4097
rect 86862 4088 86868 4140
rect 86920 4128 86926 4140
rect 87141 4131 87199 4137
rect 87141 4128 87153 4131
rect 86920 4100 87153 4128
rect 86920 4088 86926 4100
rect 87141 4097 87153 4100
rect 87187 4097 87199 4131
rect 87690 4128 87696 4140
rect 87651 4100 87696 4128
rect 87141 4091 87199 4097
rect 87690 4088 87696 4100
rect 87748 4088 87754 4140
rect 87800 4128 87828 4168
rect 87874 4128 87880 4140
rect 87800 4100 87880 4128
rect 87874 4088 87880 4100
rect 87932 4088 87938 4140
rect 88245 4131 88303 4137
rect 88245 4097 88257 4131
rect 88291 4097 88303 4131
rect 88245 4091 88303 4097
rect 71240 4032 72556 4060
rect 46532 3964 63724 3992
rect 46532 3952 46538 3964
rect 63862 3952 63868 4004
rect 63920 3992 63926 4004
rect 72528 3992 72556 4032
rect 72602 4020 72608 4072
rect 72660 4060 72666 4072
rect 88260 4060 88288 4091
rect 72660 4032 88288 4060
rect 72660 4020 72666 4032
rect 81526 3992 81532 4004
rect 63920 3964 72188 3992
rect 72528 3964 81532 3992
rect 63920 3952 63926 3964
rect 6886 3896 46152 3924
rect 46290 3884 46296 3936
rect 46348 3924 46354 3936
rect 49694 3924 49700 3936
rect 46348 3896 49700 3924
rect 46348 3884 46354 3896
rect 49694 3884 49700 3896
rect 49752 3884 49758 3936
rect 51261 3927 51319 3933
rect 51261 3893 51273 3927
rect 51307 3924 51319 3927
rect 51626 3924 51632 3936
rect 51307 3896 51632 3924
rect 51307 3893 51319 3896
rect 51261 3887 51319 3893
rect 51626 3884 51632 3896
rect 51684 3884 51690 3936
rect 59630 3924 59636 3936
rect 59591 3896 59636 3924
rect 59630 3884 59636 3896
rect 59688 3884 59694 3936
rect 71501 3927 71559 3933
rect 71501 3893 71513 3927
rect 71547 3924 71559 3927
rect 71590 3924 71596 3936
rect 71547 3896 71596 3924
rect 71547 3893 71559 3896
rect 71501 3887 71559 3893
rect 71590 3884 71596 3896
rect 71648 3884 71654 3936
rect 72160 3924 72188 3964
rect 81526 3952 81532 3964
rect 81584 3952 81590 4004
rect 87509 3995 87567 4001
rect 87509 3961 87521 3995
rect 87555 3992 87567 3995
rect 88242 3992 88248 4004
rect 87555 3964 88248 3992
rect 87555 3961 87567 3964
rect 87509 3955 87567 3961
rect 88242 3952 88248 3964
rect 88300 3952 88306 4004
rect 86589 3927 86647 3933
rect 86589 3924 86601 3927
rect 72160 3896 86601 3924
rect 86589 3893 86601 3896
rect 86635 3924 86647 3927
rect 86862 3924 86868 3936
rect 86635 3896 86868 3924
rect 86635 3893 86647 3896
rect 86589 3887 86647 3893
rect 86862 3884 86868 3896
rect 86920 3884 86926 3936
rect 86957 3927 87015 3933
rect 86957 3893 86969 3927
rect 87003 3924 87015 3927
rect 87874 3924 87880 3936
rect 87003 3896 87880 3924
rect 87003 3893 87015 3896
rect 86957 3887 87015 3893
rect 87874 3884 87880 3896
rect 87932 3884 87938 3936
rect 88058 3924 88064 3936
rect 88019 3896 88064 3924
rect 88058 3884 88064 3896
rect 88116 3884 88122 3936
rect 1104 3834 88872 3856
rect 1104 3782 11924 3834
rect 11976 3782 11988 3834
rect 12040 3782 12052 3834
rect 12104 3782 12116 3834
rect 12168 3782 12180 3834
rect 12232 3782 33872 3834
rect 33924 3782 33936 3834
rect 33988 3782 34000 3834
rect 34052 3782 34064 3834
rect 34116 3782 34128 3834
rect 34180 3782 55820 3834
rect 55872 3782 55884 3834
rect 55936 3782 55948 3834
rect 56000 3782 56012 3834
rect 56064 3782 56076 3834
rect 56128 3782 77768 3834
rect 77820 3782 77832 3834
rect 77884 3782 77896 3834
rect 77948 3782 77960 3834
rect 78012 3782 78024 3834
rect 78076 3782 88872 3834
rect 1104 3760 88872 3782
rect 17218 3680 17224 3732
rect 17276 3720 17282 3732
rect 27433 3723 27491 3729
rect 27433 3720 27445 3723
rect 17276 3692 27445 3720
rect 17276 3680 17282 3692
rect 27433 3689 27445 3692
rect 27479 3689 27491 3723
rect 27433 3683 27491 3689
rect 27890 3680 27896 3732
rect 27948 3720 27954 3732
rect 29178 3720 29184 3732
rect 27948 3692 29184 3720
rect 27948 3680 27954 3692
rect 29178 3680 29184 3692
rect 29236 3680 29242 3732
rect 30834 3720 30840 3732
rect 30795 3692 30840 3720
rect 30834 3680 30840 3692
rect 30892 3720 30898 3732
rect 31386 3720 31392 3732
rect 30892 3692 31392 3720
rect 30892 3680 30898 3692
rect 31386 3680 31392 3692
rect 31444 3680 31450 3732
rect 31478 3680 31484 3732
rect 31536 3720 31542 3732
rect 34698 3720 34704 3732
rect 31536 3692 34704 3720
rect 31536 3680 31542 3692
rect 34698 3680 34704 3692
rect 34756 3680 34762 3732
rect 34882 3680 34888 3732
rect 34940 3720 34946 3732
rect 42610 3720 42616 3732
rect 34940 3692 42616 3720
rect 34940 3680 34946 3692
rect 42610 3680 42616 3692
rect 42668 3680 42674 3732
rect 42702 3680 42708 3732
rect 42760 3720 42766 3732
rect 46290 3720 46296 3732
rect 42760 3692 46296 3720
rect 42760 3680 42766 3692
rect 46290 3680 46296 3692
rect 46348 3680 46354 3732
rect 47854 3680 47860 3732
rect 47912 3720 47918 3732
rect 49053 3723 49111 3729
rect 47912 3692 47992 3720
rect 47912 3680 47918 3692
rect 658 3612 664 3664
rect 716 3652 722 3664
rect 2501 3655 2559 3661
rect 2501 3652 2513 3655
rect 716 3624 2513 3652
rect 716 3612 722 3624
rect 2501 3621 2513 3624
rect 2547 3621 2559 3655
rect 2501 3615 2559 3621
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10008 3624 19334 3652
rect 10008 3612 10014 3624
rect 11698 3584 11704 3596
rect 1596 3556 11704 3584
rect 1596 3525 1624 3556
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 19306 3584 19334 3624
rect 22738 3612 22744 3664
rect 22796 3652 22802 3664
rect 41874 3652 41880 3664
rect 22796 3624 41880 3652
rect 22796 3612 22802 3624
rect 41874 3612 41880 3624
rect 41932 3612 41938 3664
rect 19306 3556 27384 3584
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 3510 3516 3516 3528
rect 2731 3488 3516 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 2148 3448 2176 3479
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 18230 3516 18236 3528
rect 9364 3488 18236 3516
rect 9364 3476 9370 3488
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 24394 3516 24400 3528
rect 24355 3488 24400 3516
rect 24394 3476 24400 3488
rect 24452 3476 24458 3528
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 24946 3476 24952 3528
rect 25004 3516 25010 3528
rect 26053 3519 26111 3525
rect 26053 3516 26065 3519
rect 25004 3488 26065 3516
rect 25004 3476 25010 3488
rect 26053 3485 26065 3488
rect 26099 3485 26111 3519
rect 26694 3516 26700 3528
rect 26655 3488 26700 3516
rect 26053 3479 26111 3485
rect 26694 3476 26700 3488
rect 26752 3476 26758 3528
rect 27157 3519 27215 3525
rect 27157 3485 27169 3519
rect 27203 3485 27215 3519
rect 27157 3479 27215 3485
rect 27249 3519 27307 3525
rect 27249 3485 27261 3519
rect 27295 3485 27307 3519
rect 27356 3516 27384 3556
rect 28368 3556 33456 3584
rect 28368 3516 28396 3556
rect 28445 3519 28503 3525
rect 28445 3516 28457 3519
rect 27356 3488 28457 3516
rect 27249 3479 27307 3485
rect 28445 3485 28457 3488
rect 28491 3485 28503 3519
rect 28445 3479 28503 3485
rect 4982 3448 4988 3460
rect 2148 3420 4988 3448
rect 4982 3408 4988 3420
rect 5040 3448 5046 3460
rect 5040 3420 6914 3448
rect 5040 3408 5046 3420
rect 1394 3380 1400 3392
rect 1355 3352 1400 3380
rect 1394 3340 1400 3352
rect 1452 3340 1458 3392
rect 1486 3340 1492 3392
rect 1544 3380 1550 3392
rect 1949 3383 2007 3389
rect 1949 3380 1961 3383
rect 1544 3352 1961 3380
rect 1544 3340 1550 3352
rect 1949 3349 1961 3352
rect 1995 3349 2007 3383
rect 6886 3380 6914 3420
rect 13814 3408 13820 3460
rect 13872 3448 13878 3460
rect 20714 3448 20720 3460
rect 13872 3420 20720 3448
rect 13872 3408 13878 3420
rect 20714 3408 20720 3420
rect 20772 3408 20778 3460
rect 21174 3380 21180 3392
rect 6886 3352 21180 3380
rect 1949 3343 2007 3349
rect 21174 3340 21180 3352
rect 21232 3340 21238 3392
rect 24762 3380 24768 3392
rect 24723 3352 24768 3380
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 25774 3340 25780 3392
rect 25832 3380 25838 3392
rect 25869 3383 25927 3389
rect 25869 3380 25881 3383
rect 25832 3352 25881 3380
rect 25832 3340 25838 3352
rect 25869 3349 25881 3352
rect 25915 3349 25927 3383
rect 25869 3343 25927 3349
rect 26513 3383 26571 3389
rect 26513 3349 26525 3383
rect 26559 3380 26571 3383
rect 26602 3380 26608 3392
rect 26559 3352 26608 3380
rect 26559 3349 26571 3352
rect 26513 3343 26571 3349
rect 26602 3340 26608 3352
rect 26660 3340 26666 3392
rect 27172 3380 27200 3479
rect 27264 3448 27292 3479
rect 28534 3476 28540 3528
rect 28592 3516 28598 3528
rect 30742 3516 30748 3528
rect 28592 3488 30748 3516
rect 28592 3476 28598 3488
rect 30742 3476 30748 3488
rect 30800 3476 30806 3528
rect 31202 3516 31208 3528
rect 31163 3488 31208 3516
rect 31202 3476 31208 3488
rect 31260 3476 31266 3528
rect 31386 3516 31392 3528
rect 31347 3488 31392 3516
rect 31386 3476 31392 3488
rect 31444 3476 31450 3528
rect 33042 3516 33048 3528
rect 33003 3488 33048 3516
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33428 3516 33456 3556
rect 33502 3544 33508 3596
rect 33560 3584 33566 3596
rect 33965 3587 34023 3593
rect 33965 3584 33977 3587
rect 33560 3556 33977 3584
rect 33560 3544 33566 3556
rect 33965 3553 33977 3556
rect 34011 3553 34023 3587
rect 33965 3547 34023 3553
rect 35526 3544 35532 3596
rect 35584 3584 35590 3596
rect 38102 3584 38108 3596
rect 35584 3556 38108 3584
rect 35584 3544 35590 3556
rect 38102 3544 38108 3556
rect 38160 3544 38166 3596
rect 39298 3544 39304 3596
rect 39356 3584 39362 3596
rect 41414 3584 41420 3596
rect 39356 3556 41420 3584
rect 39356 3544 39362 3556
rect 41414 3544 41420 3556
rect 41472 3584 41478 3596
rect 42702 3584 42708 3596
rect 41472 3556 42708 3584
rect 41472 3544 41478 3556
rect 42702 3544 42708 3556
rect 42760 3544 42766 3596
rect 45370 3544 45376 3596
rect 45428 3584 45434 3596
rect 47486 3584 47492 3596
rect 45428 3556 47492 3584
rect 45428 3544 45434 3556
rect 47486 3544 47492 3556
rect 47544 3544 47550 3596
rect 47765 3587 47823 3593
rect 47765 3553 47777 3587
rect 47811 3584 47823 3587
rect 47964 3584 47992 3692
rect 49053 3689 49065 3723
rect 49099 3720 49111 3723
rect 49602 3720 49608 3732
rect 49099 3692 49608 3720
rect 49099 3689 49111 3692
rect 49053 3683 49111 3689
rect 49602 3680 49608 3692
rect 49660 3680 49666 3732
rect 49694 3680 49700 3732
rect 49752 3720 49758 3732
rect 49752 3692 60734 3720
rect 49752 3680 49758 3692
rect 48222 3612 48228 3664
rect 48280 3652 48286 3664
rect 51350 3652 51356 3664
rect 48280 3624 51356 3652
rect 48280 3612 48286 3624
rect 51350 3612 51356 3624
rect 51408 3612 51414 3664
rect 60706 3652 60734 3692
rect 64138 3680 64144 3732
rect 64196 3720 64202 3732
rect 87782 3720 87788 3732
rect 64196 3692 87788 3720
rect 64196 3680 64202 3692
rect 87782 3680 87788 3692
rect 87840 3680 87846 3732
rect 87874 3680 87880 3732
rect 87932 3720 87938 3732
rect 89530 3720 89536 3732
rect 87932 3692 89536 3720
rect 87932 3680 87938 3692
rect 89530 3680 89536 3692
rect 89588 3680 89594 3732
rect 76742 3652 76748 3664
rect 60706 3624 76748 3652
rect 76742 3612 76748 3624
rect 76800 3612 76806 3664
rect 86405 3655 86463 3661
rect 86405 3621 86417 3655
rect 86451 3652 86463 3655
rect 86678 3652 86684 3664
rect 86451 3624 86684 3652
rect 86451 3621 86463 3624
rect 86405 3615 86463 3621
rect 86678 3612 86684 3624
rect 86736 3612 86742 3664
rect 87598 3612 87604 3664
rect 87656 3652 87662 3664
rect 88337 3655 88395 3661
rect 88337 3652 88349 3655
rect 87656 3624 88349 3652
rect 87656 3612 87662 3624
rect 88337 3621 88349 3624
rect 88383 3621 88395 3655
rect 88337 3615 88395 3621
rect 47811 3556 47992 3584
rect 47811 3553 47823 3556
rect 47765 3547 47823 3553
rect 48130 3544 48136 3596
rect 48188 3584 48194 3596
rect 48188 3556 49464 3584
rect 48188 3544 48194 3556
rect 33152 3488 33364 3516
rect 33428 3488 36492 3516
rect 30006 3448 30012 3460
rect 27264 3420 28396 3448
rect 27706 3380 27712 3392
rect 27172 3352 27712 3380
rect 27706 3340 27712 3352
rect 27764 3340 27770 3392
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28261 3383 28319 3389
rect 28261 3380 28273 3383
rect 27948 3352 28273 3380
rect 27948 3340 27954 3352
rect 28261 3349 28273 3352
rect 28307 3349 28319 3383
rect 28368 3380 28396 3420
rect 28644 3420 30012 3448
rect 28644 3380 28672 3420
rect 30006 3408 30012 3420
rect 30064 3448 30070 3460
rect 30282 3448 30288 3460
rect 30064 3420 30288 3448
rect 30064 3408 30070 3420
rect 30282 3408 30288 3420
rect 30340 3408 30346 3460
rect 31294 3408 31300 3460
rect 31352 3448 31358 3460
rect 33152 3448 33180 3488
rect 31352 3420 33180 3448
rect 33336 3448 33364 3488
rect 33781 3451 33839 3457
rect 33781 3448 33793 3451
rect 33336 3420 33793 3448
rect 31352 3408 31358 3420
rect 33781 3417 33793 3420
rect 33827 3448 33839 3451
rect 33962 3448 33968 3460
rect 33827 3420 33968 3448
rect 33827 3417 33839 3420
rect 33781 3411 33839 3417
rect 33962 3408 33968 3420
rect 34020 3408 34026 3460
rect 36464 3448 36492 3488
rect 36538 3476 36544 3528
rect 36596 3516 36602 3528
rect 43438 3516 43444 3528
rect 36596 3488 43444 3516
rect 36596 3476 36602 3488
rect 43438 3476 43444 3488
rect 43496 3476 43502 3528
rect 46014 3476 46020 3528
rect 46072 3516 46078 3528
rect 48866 3516 48872 3528
rect 46072 3488 48872 3516
rect 46072 3476 46078 3488
rect 48866 3476 48872 3488
rect 48924 3476 48930 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49237 3519 49295 3525
rect 49237 3516 49249 3519
rect 49016 3488 49249 3516
rect 49016 3476 49022 3488
rect 49237 3485 49249 3488
rect 49283 3485 49295 3519
rect 49237 3479 49295 3485
rect 37274 3448 37280 3460
rect 36464 3420 37280 3448
rect 37274 3408 37280 3420
rect 37332 3408 37338 3460
rect 41230 3408 41236 3460
rect 41288 3448 41294 3460
rect 48682 3448 48688 3460
rect 41288 3420 48688 3448
rect 41288 3408 41294 3420
rect 48682 3408 48688 3420
rect 48740 3408 48746 3460
rect 28368 3352 28672 3380
rect 28261 3343 28319 3349
rect 28718 3340 28724 3392
rect 28776 3380 28782 3392
rect 31478 3380 31484 3392
rect 28776 3352 31484 3380
rect 28776 3340 28782 3352
rect 31478 3340 31484 3352
rect 31536 3340 31542 3392
rect 31573 3383 31631 3389
rect 31573 3349 31585 3383
rect 31619 3380 31631 3383
rect 31662 3380 31668 3392
rect 31619 3352 31668 3380
rect 31619 3349 31631 3352
rect 31573 3343 31631 3349
rect 31662 3340 31668 3352
rect 31720 3340 31726 3392
rect 32582 3340 32588 3392
rect 32640 3380 32646 3392
rect 32861 3383 32919 3389
rect 32861 3380 32873 3383
rect 32640 3352 32873 3380
rect 32640 3340 32646 3352
rect 32861 3349 32873 3352
rect 32907 3349 32919 3383
rect 32861 3343 32919 3349
rect 33042 3340 33048 3392
rect 33100 3380 33106 3392
rect 33413 3383 33471 3389
rect 33413 3380 33425 3383
rect 33100 3352 33425 3380
rect 33100 3340 33106 3352
rect 33413 3349 33425 3352
rect 33459 3349 33471 3383
rect 33413 3343 33471 3349
rect 33873 3383 33931 3389
rect 33873 3349 33885 3383
rect 33919 3380 33931 3383
rect 39390 3380 39396 3392
rect 33919 3352 39396 3380
rect 33919 3349 33931 3352
rect 33873 3343 33931 3349
rect 39390 3340 39396 3352
rect 39448 3340 39454 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 45186 3380 45192 3392
rect 41932 3352 45192 3380
rect 41932 3340 41938 3352
rect 45186 3340 45192 3352
rect 45244 3340 45250 3392
rect 47118 3380 47124 3392
rect 47079 3352 47124 3380
rect 47118 3340 47124 3352
rect 47176 3340 47182 3392
rect 47486 3380 47492 3392
rect 47447 3352 47492 3380
rect 47486 3340 47492 3352
rect 47544 3340 47550 3392
rect 47581 3383 47639 3389
rect 47581 3349 47593 3383
rect 47627 3380 47639 3383
rect 49234 3380 49240 3392
rect 47627 3352 49240 3380
rect 47627 3349 47639 3352
rect 47581 3343 47639 3349
rect 49234 3340 49240 3352
rect 49292 3340 49298 3392
rect 49436 3380 49464 3556
rect 49694 3544 49700 3596
rect 49752 3584 49758 3596
rect 50154 3584 50160 3596
rect 49752 3556 50160 3584
rect 49752 3544 49758 3556
rect 50154 3544 50160 3556
rect 50212 3584 50218 3596
rect 51537 3587 51595 3593
rect 51537 3584 51549 3587
rect 50212 3556 51549 3584
rect 50212 3544 50218 3556
rect 51537 3553 51549 3556
rect 51583 3553 51595 3587
rect 51537 3547 51595 3553
rect 52546 3544 52552 3596
rect 52604 3584 52610 3596
rect 58342 3584 58348 3596
rect 52604 3556 58348 3584
rect 52604 3544 52610 3556
rect 58342 3544 58348 3556
rect 58400 3544 58406 3596
rect 58618 3544 58624 3596
rect 58676 3584 58682 3596
rect 73522 3584 73528 3596
rect 58676 3556 73528 3584
rect 58676 3544 58682 3556
rect 73522 3544 73528 3556
rect 73580 3544 73586 3596
rect 50246 3476 50252 3528
rect 50304 3516 50310 3528
rect 50341 3519 50399 3525
rect 50341 3516 50353 3519
rect 50304 3488 50353 3516
rect 50304 3476 50310 3488
rect 50341 3485 50353 3488
rect 50387 3485 50399 3519
rect 50522 3516 50528 3528
rect 50483 3488 50528 3516
rect 50341 3479 50399 3485
rect 50522 3476 50528 3488
rect 50580 3476 50586 3528
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 62390 3516 62396 3528
rect 51408 3488 62396 3516
rect 51408 3476 51414 3488
rect 62390 3476 62396 3488
rect 62448 3476 62454 3528
rect 70210 3476 70216 3528
rect 70268 3516 70274 3528
rect 75178 3516 75184 3528
rect 70268 3488 75184 3516
rect 70268 3476 70274 3488
rect 75178 3476 75184 3488
rect 75236 3476 75242 3528
rect 86586 3516 86592 3528
rect 86547 3488 86592 3516
rect 86586 3476 86592 3488
rect 86644 3516 86650 3528
rect 86865 3519 86923 3525
rect 86865 3516 86877 3519
rect 86644 3488 86877 3516
rect 86644 3476 86650 3488
rect 86865 3485 86877 3488
rect 86911 3485 86923 3519
rect 86865 3479 86923 3485
rect 88061 3519 88119 3525
rect 88061 3485 88073 3519
rect 88107 3516 88119 3519
rect 88150 3516 88156 3528
rect 88107 3488 88156 3516
rect 88107 3485 88119 3488
rect 88061 3479 88119 3485
rect 88150 3476 88156 3488
rect 88208 3476 88214 3528
rect 88521 3519 88579 3525
rect 88521 3485 88533 3519
rect 88567 3485 88579 3519
rect 88521 3479 88579 3485
rect 49510 3408 49516 3460
rect 49568 3448 49574 3460
rect 50709 3451 50767 3457
rect 50709 3448 50721 3451
rect 49568 3420 50721 3448
rect 49568 3408 49574 3420
rect 50709 3417 50721 3420
rect 50755 3417 50767 3451
rect 50709 3411 50767 3417
rect 51442 3408 51448 3460
rect 51500 3448 51506 3460
rect 51782 3451 51840 3457
rect 51782 3448 51794 3451
rect 51500 3420 51794 3448
rect 51500 3408 51506 3420
rect 51782 3417 51794 3420
rect 51828 3417 51840 3451
rect 51782 3411 51840 3417
rect 51920 3420 53144 3448
rect 51920 3380 51948 3420
rect 49436 3352 51948 3380
rect 52914 3340 52920 3392
rect 52972 3380 52978 3392
rect 53116 3380 53144 3420
rect 53190 3408 53196 3460
rect 53248 3448 53254 3460
rect 87325 3451 87383 3457
rect 87325 3448 87337 3451
rect 53248 3420 87337 3448
rect 53248 3408 53254 3420
rect 87325 3417 87337 3420
rect 87371 3448 87383 3451
rect 88536 3448 88564 3479
rect 87371 3420 88564 3448
rect 87371 3417 87383 3420
rect 87325 3411 87383 3417
rect 87693 3383 87751 3389
rect 87693 3380 87705 3383
rect 52972 3352 53017 3380
rect 53116 3352 87705 3380
rect 52972 3340 52978 3352
rect 87693 3349 87705 3352
rect 87739 3380 87751 3383
rect 87739 3352 88932 3380
rect 87739 3349 87751 3352
rect 87693 3343 87751 3349
rect 1104 3290 88872 3312
rect 1104 3238 22898 3290
rect 22950 3238 22962 3290
rect 23014 3238 23026 3290
rect 23078 3238 23090 3290
rect 23142 3238 23154 3290
rect 23206 3238 44846 3290
rect 44898 3238 44910 3290
rect 44962 3238 44974 3290
rect 45026 3238 45038 3290
rect 45090 3238 45102 3290
rect 45154 3238 66794 3290
rect 66846 3238 66858 3290
rect 66910 3238 66922 3290
rect 66974 3238 66986 3290
rect 67038 3238 67050 3290
rect 67102 3238 88872 3290
rect 1104 3216 88872 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 1670 3176 1676 3188
rect 1627 3148 1676 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 3510 3176 3516 3188
rect 3471 3148 3516 3176
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 16574 3176 16580 3188
rect 3620 3148 16580 3176
rect 14 3000 20 3052
rect 72 3040 78 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 72 3012 1409 3040
rect 72 3000 78 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3620 3040 3648 3148
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 24210 3176 24216 3188
rect 17144 3148 24216 3176
rect 4522 3068 4528 3120
rect 4580 3108 4586 3120
rect 9306 3108 9312 3120
rect 4580 3080 9312 3108
rect 4580 3068 4586 3080
rect 9306 3068 9312 3080
rect 9364 3068 9370 3120
rect 9416 3080 12296 3108
rect 3191 3012 3648 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 2240 2904 2268 3003
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 4798 3040 4804 3052
rect 3752 3012 3845 3040
rect 4759 3012 4804 3040
rect 3752 3000 3758 3012
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 4982 3040 4988 3052
rect 4943 3012 4988 3040
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 5215 3012 5733 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 5721 3009 5733 3012
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3040 6791 3043
rect 7098 3040 7104 3052
rect 6779 3012 7104 3040
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 9416 3049 9444 3080
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9950 3040 9956 3052
rect 9911 3012 9956 3040
rect 9401 3003 9459 3009
rect 3712 2972 3740 3000
rect 9416 2972 9444 3003
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 3712 2944 9444 2972
rect 4522 2904 4528 2916
rect 2240 2876 4528 2904
rect 4522 2864 4528 2876
rect 4580 2864 4586 2916
rect 9217 2907 9275 2913
rect 9217 2873 9229 2907
rect 9263 2904 9275 2907
rect 9950 2904 9956 2916
rect 9263 2876 9956 2904
rect 9263 2873 9275 2876
rect 9217 2867 9275 2873
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 12176 2904 12204 3003
rect 12268 2972 12296 3080
rect 13814 3040 13820 3052
rect 13775 3012 13820 3040
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16816 3012 17049 3040
rect 16816 3000 16822 3012
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 17144 2972 17172 3148
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 46014 3176 46020 3188
rect 26068 3148 46020 3176
rect 26068 3108 26096 3148
rect 46014 3136 46020 3148
rect 46072 3136 46078 3188
rect 46937 3179 46995 3185
rect 46937 3145 46949 3179
rect 46983 3176 46995 3179
rect 46983 3148 47716 3176
rect 46983 3145 46995 3148
rect 46937 3139 46995 3145
rect 19444 3080 26096 3108
rect 19444 3049 19472 3080
rect 26142 3068 26148 3120
rect 26200 3108 26206 3120
rect 31754 3108 31760 3120
rect 26200 3080 31760 3108
rect 26200 3068 26206 3080
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3040 17739 3043
rect 19429 3043 19487 3049
rect 17727 3012 19288 3040
rect 17727 3009 17739 3012
rect 17681 3003 17739 3009
rect 12268 2944 17172 2972
rect 17218 2904 17224 2916
rect 12176 2876 17224 2904
rect 17218 2864 17224 2876
rect 17276 2864 17282 2916
rect 17954 2904 17960 2916
rect 17328 2876 17960 2904
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 2041 2839 2099 2845
rect 2041 2836 2053 2839
rect 2004 2808 2053 2836
rect 2004 2796 2010 2808
rect 2041 2805 2053 2808
rect 2087 2805 2099 2839
rect 2041 2799 2099 2805
rect 2961 2839 3019 2845
rect 2961 2805 2973 2839
rect 3007 2836 3019 2839
rect 4890 2836 4896 2848
rect 3007 2808 4896 2836
rect 3007 2805 3019 2808
rect 2961 2799 3019 2805
rect 4890 2796 4896 2808
rect 4948 2796 4954 2848
rect 5534 2836 5540 2848
rect 5495 2808 5540 2836
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 6512 2808 6561 2836
rect 6512 2796 6518 2808
rect 6549 2805 6561 2808
rect 6595 2805 6607 2839
rect 9766 2836 9772 2848
rect 9727 2808 9772 2836
rect 6549 2799 6607 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 10226 2796 10232 2848
rect 10284 2836 10290 2848
rect 11977 2839 12035 2845
rect 11977 2836 11989 2839
rect 10284 2808 11989 2836
rect 10284 2796 10290 2808
rect 11977 2805 11989 2808
rect 12023 2805 12035 2839
rect 11977 2799 12035 2805
rect 13538 2796 13544 2848
rect 13596 2836 13602 2848
rect 13633 2839 13691 2845
rect 13633 2836 13645 2839
rect 13596 2808 13645 2836
rect 13596 2796 13602 2808
rect 13633 2805 13645 2808
rect 13679 2805 13691 2839
rect 13633 2799 13691 2805
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 17328 2836 17356 2876
rect 17954 2864 17960 2876
rect 18012 2864 18018 2916
rect 19260 2913 19288 3012
rect 19429 3009 19441 3043
rect 19475 3009 19487 3043
rect 19429 3003 19487 3009
rect 19797 3043 19855 3049
rect 19797 3009 19809 3043
rect 19843 3040 19855 3043
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 19843 3012 20269 3040
rect 19843 3009 19855 3012
rect 19797 3003 19855 3009
rect 20257 3009 20269 3012
rect 20303 3040 20315 3043
rect 22738 3040 22744 3052
rect 20303 3012 22744 3040
rect 20303 3009 20315 3012
rect 20257 3003 20315 3009
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 23017 3043 23075 3049
rect 23017 3009 23029 3043
rect 23063 3040 23075 3043
rect 24762 3040 24768 3052
rect 23063 3012 24768 3040
rect 23063 3009 23075 3012
rect 23017 3003 23075 3009
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 25406 3040 25412 3052
rect 25367 3012 25412 3040
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 25958 3040 25964 3052
rect 25871 3012 25964 3040
rect 25958 3000 25964 3012
rect 26016 3000 26022 3052
rect 26326 3040 26332 3052
rect 26287 3012 26332 3040
rect 26326 3000 26332 3012
rect 26384 3000 26390 3052
rect 27433 3043 27491 3049
rect 27433 3009 27445 3043
rect 27479 3040 27491 3043
rect 27706 3040 27712 3052
rect 27479 3012 27712 3040
rect 27479 3009 27491 3012
rect 27433 3003 27491 3009
rect 27706 3000 27712 3012
rect 27764 3000 27770 3052
rect 27816 3049 27844 3080
rect 31754 3068 31760 3080
rect 31812 3108 31818 3120
rect 33962 3108 33968 3120
rect 31812 3080 32352 3108
rect 33923 3080 33968 3108
rect 31812 3068 31818 3080
rect 27801 3043 27859 3049
rect 27801 3009 27813 3043
rect 27847 3009 27859 3043
rect 28057 3043 28115 3049
rect 28057 3040 28069 3043
rect 27801 3003 27859 3009
rect 27908 3012 28069 3040
rect 24210 2932 24216 2984
rect 24268 2972 24274 2984
rect 25976 2972 26004 3000
rect 24268 2944 26004 2972
rect 24268 2932 24274 2944
rect 26234 2932 26240 2984
rect 26292 2972 26298 2984
rect 26421 2975 26479 2981
rect 26421 2972 26433 2975
rect 26292 2944 26433 2972
rect 26292 2932 26298 2944
rect 26421 2941 26433 2944
rect 26467 2941 26479 2975
rect 27908 2972 27936 3012
rect 28057 3009 28069 3012
rect 28103 3009 28115 3043
rect 29825 3043 29883 3049
rect 29825 3040 29837 3043
rect 28057 3003 28115 3009
rect 29380 3012 29837 3040
rect 26421 2935 26479 2941
rect 27264 2944 27936 2972
rect 19245 2907 19303 2913
rect 19245 2873 19257 2907
rect 19291 2873 19303 2907
rect 19245 2867 19303 2873
rect 24394 2864 24400 2916
rect 24452 2904 24458 2916
rect 27264 2913 27292 2944
rect 27249 2907 27307 2913
rect 24452 2876 25912 2904
rect 24452 2864 24458 2876
rect 16899 2808 17356 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 17497 2839 17555 2845
rect 17497 2836 17509 2839
rect 17460 2808 17509 2836
rect 17460 2796 17466 2808
rect 17497 2805 17509 2808
rect 17543 2805 17555 2839
rect 17497 2799 17555 2805
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 20073 2839 20131 2845
rect 20073 2836 20085 2839
rect 20036 2808 20085 2836
rect 20036 2796 20042 2808
rect 20073 2805 20085 2808
rect 20119 2805 20131 2839
rect 22830 2836 22836 2848
rect 22791 2808 22836 2836
rect 20073 2799 20131 2805
rect 22830 2796 22836 2808
rect 22888 2796 22894 2848
rect 25130 2796 25136 2848
rect 25188 2836 25194 2848
rect 25225 2839 25283 2845
rect 25225 2836 25237 2839
rect 25188 2808 25237 2836
rect 25188 2796 25194 2808
rect 25225 2805 25237 2808
rect 25271 2805 25283 2839
rect 25225 2799 25283 2805
rect 25406 2796 25412 2848
rect 25464 2836 25470 2848
rect 25777 2839 25835 2845
rect 25777 2836 25789 2839
rect 25464 2808 25789 2836
rect 25464 2796 25470 2808
rect 25777 2805 25789 2808
rect 25823 2805 25835 2839
rect 25884 2836 25912 2876
rect 27249 2873 27261 2907
rect 27295 2873 27307 2907
rect 29178 2904 29184 2916
rect 29091 2876 29184 2904
rect 27249 2867 27307 2873
rect 29178 2864 29184 2876
rect 29236 2904 29242 2916
rect 29380 2904 29408 3012
rect 29825 3009 29837 3012
rect 29871 3009 29883 3043
rect 29825 3003 29883 3009
rect 30009 3043 30067 3049
rect 30009 3009 30021 3043
rect 30055 3040 30067 3043
rect 30561 3043 30619 3049
rect 30561 3040 30573 3043
rect 30055 3012 30573 3040
rect 30055 3009 30067 3012
rect 30009 3003 30067 3009
rect 30561 3009 30573 3012
rect 30607 3009 30619 3043
rect 31662 3040 31668 3052
rect 31623 3012 31668 3040
rect 30561 3003 30619 3009
rect 31662 3000 31668 3012
rect 31720 3000 31726 3052
rect 32324 3049 32352 3080
rect 33962 3068 33968 3080
rect 34020 3068 34026 3120
rect 34698 3068 34704 3120
rect 34756 3108 34762 3120
rect 39114 3108 39120 3120
rect 34756 3080 39120 3108
rect 34756 3068 34762 3080
rect 39114 3068 39120 3080
rect 39172 3108 39178 3120
rect 39669 3111 39727 3117
rect 39172 3080 39528 3108
rect 39172 3068 39178 3080
rect 32309 3043 32367 3049
rect 32309 3009 32321 3043
rect 32355 3009 32367 3043
rect 32582 3040 32588 3052
rect 32543 3012 32588 3040
rect 32309 3003 32367 3009
rect 32582 3000 32588 3012
rect 32640 3000 32646 3052
rect 34333 3043 34391 3049
rect 34333 3009 34345 3043
rect 34379 3040 34391 3043
rect 34793 3043 34851 3049
rect 34793 3040 34805 3043
rect 34379 3012 34805 3040
rect 34379 3009 34391 3012
rect 34333 3003 34391 3009
rect 34793 3009 34805 3012
rect 34839 3040 34851 3043
rect 34882 3040 34888 3052
rect 34839 3012 34888 3040
rect 34839 3009 34851 3012
rect 34793 3003 34851 3009
rect 34882 3000 34888 3012
rect 34940 3000 34946 3052
rect 38657 3043 38715 3049
rect 38657 3009 38669 3043
rect 38703 3040 38715 3043
rect 38930 3040 38936 3052
rect 38703 3012 38936 3040
rect 38703 3009 38715 3012
rect 38657 3003 38715 3009
rect 38930 3000 38936 3012
rect 38988 3000 38994 3052
rect 39025 3043 39083 3049
rect 39025 3009 39037 3043
rect 39071 3040 39083 3043
rect 39298 3040 39304 3052
rect 39071 3012 39304 3040
rect 39071 3009 39083 3012
rect 39025 3003 39083 3009
rect 39298 3000 39304 3012
rect 39356 3000 39362 3052
rect 39500 3049 39528 3080
rect 39669 3077 39681 3111
rect 39715 3108 39727 3111
rect 39715 3080 41414 3108
rect 39715 3077 39727 3080
rect 39669 3071 39727 3077
rect 39485 3043 39543 3049
rect 39485 3009 39497 3043
rect 39531 3009 39543 3043
rect 40218 3040 40224 3052
rect 40179 3012 40224 3040
rect 39485 3003 39543 3009
rect 40218 3000 40224 3012
rect 40276 3000 40282 3052
rect 41386 3040 41414 3080
rect 41598 3068 41604 3120
rect 41656 3108 41662 3120
rect 43254 3108 43260 3120
rect 41656 3080 43260 3108
rect 41656 3068 41662 3080
rect 43254 3068 43260 3080
rect 43312 3068 43318 3120
rect 41969 3043 42027 3049
rect 41969 3040 41981 3043
rect 41386 3012 41981 3040
rect 41969 3009 41981 3012
rect 42015 3009 42027 3043
rect 41969 3003 42027 3009
rect 42613 3043 42671 3049
rect 42613 3009 42625 3043
rect 42659 3040 42671 3043
rect 43898 3040 43904 3052
rect 42659 3012 43904 3040
rect 42659 3009 42671 3012
rect 42613 3003 42671 3009
rect 43898 3000 43904 3012
rect 43956 3000 43962 3052
rect 47118 3040 47124 3052
rect 47079 3012 47124 3040
rect 47118 3000 47124 3012
rect 47176 3000 47182 3052
rect 47581 3043 47639 3049
rect 47581 3040 47593 3043
rect 47228 3012 47593 3040
rect 29641 2975 29699 2981
rect 29641 2941 29653 2975
rect 29687 2972 29699 2975
rect 29687 2944 34744 2972
rect 29687 2941 29699 2944
rect 29641 2935 29699 2941
rect 29236 2876 29408 2904
rect 29236 2864 29242 2876
rect 33502 2864 33508 2916
rect 33560 2904 33566 2916
rect 34609 2907 34667 2913
rect 34609 2904 34621 2907
rect 33560 2876 34621 2904
rect 33560 2864 33566 2876
rect 34609 2873 34621 2876
rect 34655 2873 34667 2907
rect 34716 2904 34744 2944
rect 39390 2932 39396 2984
rect 39448 2972 39454 2984
rect 46290 2972 46296 2984
rect 39448 2944 46296 2972
rect 39448 2932 39454 2944
rect 46290 2932 46296 2944
rect 46348 2932 46354 2984
rect 46382 2932 46388 2984
rect 46440 2972 46446 2984
rect 47228 2972 47256 3012
rect 47581 3009 47593 3012
rect 47627 3009 47639 3043
rect 47688 3040 47716 3148
rect 50338 3136 50344 3188
rect 50396 3176 50402 3188
rect 50985 3179 51043 3185
rect 50985 3176 50997 3179
rect 50396 3148 50997 3176
rect 50396 3136 50402 3148
rect 50985 3145 50997 3148
rect 51031 3176 51043 3179
rect 51994 3176 52000 3188
rect 51031 3148 51856 3176
rect 51955 3148 52000 3176
rect 51031 3145 51043 3148
rect 50985 3139 51043 3145
rect 49418 3068 49424 3120
rect 49476 3108 49482 3120
rect 49850 3111 49908 3117
rect 49850 3108 49862 3111
rect 49476 3080 49862 3108
rect 49476 3068 49482 3080
rect 49850 3077 49862 3080
rect 49896 3077 49908 3111
rect 51828 3108 51856 3148
rect 51994 3136 52000 3148
rect 52052 3136 52058 3188
rect 52178 3136 52184 3188
rect 52236 3176 52242 3188
rect 59630 3176 59636 3188
rect 52236 3148 59636 3176
rect 52236 3136 52242 3148
rect 59630 3136 59636 3148
rect 59688 3176 59694 3188
rect 59688 3148 61608 3176
rect 59688 3136 59694 3148
rect 51828 3080 60734 3108
rect 49850 3071 49908 3077
rect 47857 3043 47915 3049
rect 47857 3040 47869 3043
rect 47688 3012 47869 3040
rect 47581 3003 47639 3009
rect 47857 3009 47869 3012
rect 47903 3009 47915 3043
rect 49602 3040 49608 3052
rect 49563 3012 49608 3040
rect 47857 3003 47915 3009
rect 49602 3000 49608 3012
rect 49660 3000 49666 3052
rect 50246 3040 50252 3052
rect 49712 3012 50252 3040
rect 49712 2972 49740 3012
rect 50246 3000 50252 3012
rect 50304 3000 50310 3052
rect 51626 3000 51632 3052
rect 51684 3040 51690 3052
rect 52181 3043 52239 3049
rect 51684 3012 51729 3040
rect 51684 3000 51690 3012
rect 52181 3009 52193 3043
rect 52227 3009 52239 3043
rect 52181 3003 52239 3009
rect 53009 3043 53067 3049
rect 53009 3009 53021 3043
rect 53055 3040 53067 3043
rect 53469 3043 53527 3049
rect 53469 3040 53481 3043
rect 53055 3012 53481 3040
rect 53055 3009 53067 3012
rect 53009 3003 53067 3009
rect 53469 3009 53481 3012
rect 53515 3040 53527 3043
rect 53650 3040 53656 3052
rect 53515 3012 53656 3040
rect 53515 3009 53527 3012
rect 53469 3003 53527 3009
rect 46440 2944 47256 2972
rect 47596 2944 49740 2972
rect 51276 2944 51680 2972
rect 46440 2932 46446 2944
rect 41598 2904 41604 2916
rect 34716 2876 41604 2904
rect 34609 2867 34667 2873
rect 41598 2864 41604 2876
rect 41656 2864 41662 2916
rect 41785 2907 41843 2913
rect 41785 2873 41797 2907
rect 41831 2904 41843 2907
rect 43438 2904 43444 2916
rect 41831 2876 43444 2904
rect 41831 2873 41843 2876
rect 41785 2867 41843 2873
rect 43438 2864 43444 2876
rect 43496 2864 43502 2916
rect 47596 2904 47624 2944
rect 47412 2876 47624 2904
rect 29454 2836 29460 2848
rect 25884 2808 29460 2836
rect 25777 2799 25835 2805
rect 29454 2796 29460 2808
rect 29512 2796 29518 2848
rect 30374 2836 30380 2848
rect 30335 2808 30380 2836
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 31478 2836 31484 2848
rect 31439 2808 31484 2836
rect 31478 2796 31484 2808
rect 31536 2796 31542 2848
rect 35710 2796 35716 2848
rect 35768 2836 35774 2848
rect 37458 2836 37464 2848
rect 35768 2808 37464 2836
rect 35768 2796 35774 2808
rect 37458 2796 37464 2808
rect 37516 2796 37522 2848
rect 38473 2839 38531 2845
rect 38473 2805 38485 2839
rect 38519 2836 38531 2839
rect 39758 2836 39764 2848
rect 38519 2808 39764 2836
rect 38519 2805 38531 2808
rect 38473 2799 38531 2805
rect 39758 2796 39764 2808
rect 39816 2796 39822 2848
rect 39942 2796 39948 2848
rect 40000 2836 40006 2848
rect 40037 2839 40095 2845
rect 40037 2836 40049 2839
rect 40000 2808 40049 2836
rect 40000 2796 40006 2808
rect 40037 2805 40049 2808
rect 40083 2805 40095 2839
rect 40037 2799 40095 2805
rect 42429 2839 42487 2845
rect 42429 2805 42441 2839
rect 42475 2836 42487 2839
rect 42794 2836 42800 2848
rect 42475 2808 42800 2836
rect 42475 2805 42487 2808
rect 42429 2799 42487 2805
rect 42794 2796 42800 2808
rect 42852 2796 42858 2848
rect 43254 2796 43260 2848
rect 43312 2836 43318 2848
rect 47412 2836 47440 2876
rect 43312 2808 47440 2836
rect 43312 2796 43318 2808
rect 47486 2796 47492 2848
rect 47544 2836 47550 2848
rect 49145 2839 49203 2845
rect 49145 2836 49157 2839
rect 47544 2808 49157 2836
rect 47544 2796 47550 2808
rect 49145 2805 49157 2808
rect 49191 2836 49203 2839
rect 51276 2836 51304 2944
rect 51442 2904 51448 2916
rect 51403 2876 51448 2904
rect 51442 2864 51448 2876
rect 51500 2864 51506 2916
rect 51652 2904 51680 2944
rect 51718 2932 51724 2984
rect 51776 2972 51782 2984
rect 52196 2972 52224 3003
rect 53650 3000 53656 3012
rect 53708 3000 53714 3052
rect 53745 3043 53803 3049
rect 53745 3009 53757 3043
rect 53791 3009 53803 3043
rect 53745 3003 53803 3009
rect 54113 3043 54171 3049
rect 54113 3009 54125 3043
rect 54159 3009 54171 3043
rect 54113 3003 54171 3009
rect 53760 2972 53788 3003
rect 51776 2944 52224 2972
rect 53300 2944 53788 2972
rect 54128 2972 54156 3003
rect 55674 3000 55680 3052
rect 55732 3040 55738 3052
rect 55861 3043 55919 3049
rect 55861 3040 55873 3043
rect 55732 3012 55873 3040
rect 55732 3000 55738 3012
rect 55861 3009 55873 3012
rect 55907 3009 55919 3043
rect 55861 3003 55919 3009
rect 58069 3043 58127 3049
rect 58069 3009 58081 3043
rect 58115 3009 58127 3043
rect 58618 3040 58624 3052
rect 58579 3012 58624 3040
rect 58069 3003 58127 3009
rect 54938 2972 54944 2984
rect 54128 2944 54944 2972
rect 51776 2932 51782 2944
rect 51902 2904 51908 2916
rect 51652 2876 51908 2904
rect 51902 2864 51908 2876
rect 51960 2864 51966 2916
rect 52178 2864 52184 2916
rect 52236 2904 52242 2916
rect 53300 2913 53328 2944
rect 54938 2932 54944 2944
rect 54996 2972 55002 2984
rect 58084 2972 58112 3003
rect 58618 3000 58624 3012
rect 58676 3000 58682 3052
rect 54996 2944 58112 2972
rect 60706 2972 60734 3080
rect 61580 3049 61608 3148
rect 63494 3136 63500 3188
rect 63552 3176 63558 3188
rect 71409 3179 71467 3185
rect 63552 3148 64828 3176
rect 63552 3136 63558 3148
rect 61933 3111 61991 3117
rect 61933 3077 61945 3111
rect 61979 3108 61991 3111
rect 61979 3080 63908 3108
rect 61979 3077 61991 3080
rect 61933 3071 61991 3077
rect 61565 3043 61623 3049
rect 61565 3009 61577 3043
rect 61611 3009 61623 3043
rect 61565 3003 61623 3009
rect 61749 3043 61807 3049
rect 61749 3009 61761 3043
rect 61795 3009 61807 3043
rect 61749 3003 61807 3009
rect 61764 2972 61792 3003
rect 63126 3000 63132 3052
rect 63184 3040 63190 3052
rect 63880 3049 63908 3080
rect 64800 3049 64828 3148
rect 71409 3145 71421 3179
rect 71455 3145 71467 3179
rect 71409 3139 71467 3145
rect 71424 3108 71452 3139
rect 75178 3136 75184 3188
rect 75236 3176 75242 3188
rect 85945 3179 86003 3185
rect 75236 3148 84194 3176
rect 75236 3136 75242 3148
rect 76742 3108 76748 3120
rect 71424 3080 72188 3108
rect 76703 3080 76748 3108
rect 63221 3043 63279 3049
rect 63221 3040 63233 3043
rect 63184 3012 63233 3040
rect 63184 3000 63190 3012
rect 63221 3009 63233 3012
rect 63267 3040 63279 3043
rect 63497 3043 63555 3049
rect 63497 3040 63509 3043
rect 63267 3012 63509 3040
rect 63267 3009 63279 3012
rect 63221 3003 63279 3009
rect 63497 3009 63509 3012
rect 63543 3009 63555 3043
rect 63497 3003 63555 3009
rect 63865 3043 63923 3049
rect 63865 3009 63877 3043
rect 63911 3009 63923 3043
rect 63865 3003 63923 3009
rect 64785 3043 64843 3049
rect 64785 3009 64797 3043
rect 64831 3009 64843 3043
rect 64785 3003 64843 3009
rect 68741 3043 68799 3049
rect 68741 3009 68753 3043
rect 68787 3040 68799 3043
rect 71590 3040 71596 3052
rect 68787 3012 70394 3040
rect 71551 3012 71596 3040
rect 68787 3009 68799 3012
rect 68741 3003 68799 3009
rect 60706 2944 63172 2972
rect 54996 2932 55002 2944
rect 53285 2907 53343 2913
rect 52236 2876 53052 2904
rect 52236 2864 52242 2876
rect 49191 2808 51304 2836
rect 53024 2836 53052 2876
rect 53285 2873 53297 2907
rect 53331 2873 53343 2907
rect 53285 2867 53343 2873
rect 53561 2839 53619 2845
rect 53561 2836 53573 2839
rect 53024 2808 53573 2836
rect 49191 2805 49203 2808
rect 49145 2799 49203 2805
rect 53561 2805 53573 2808
rect 53607 2805 53619 2839
rect 53561 2799 53619 2805
rect 53929 2839 53987 2845
rect 53929 2805 53941 2839
rect 53975 2836 53987 2839
rect 54386 2836 54392 2848
rect 53975 2808 54392 2836
rect 53975 2805 53987 2808
rect 53929 2799 53987 2805
rect 54386 2796 54392 2808
rect 54444 2796 54450 2848
rect 55677 2839 55735 2845
rect 55677 2805 55689 2839
rect 55723 2836 55735 2839
rect 56594 2836 56600 2848
rect 55723 2808 56600 2836
rect 55723 2805 55735 2808
rect 55677 2799 55735 2805
rect 56594 2796 56600 2808
rect 56652 2796 56658 2848
rect 57885 2839 57943 2845
rect 57885 2805 57897 2839
rect 57931 2836 57943 2839
rect 58342 2836 58348 2848
rect 57931 2808 58348 2836
rect 57931 2805 57943 2808
rect 57885 2799 57943 2805
rect 58342 2796 58348 2808
rect 58400 2796 58406 2848
rect 58437 2839 58495 2845
rect 58437 2805 58449 2839
rect 58483 2836 58495 2839
rect 59170 2836 59176 2848
rect 58483 2808 59176 2836
rect 58483 2805 58495 2808
rect 58437 2799 58495 2805
rect 59170 2796 59176 2808
rect 59228 2796 59234 2848
rect 62482 2796 62488 2848
rect 62540 2836 62546 2848
rect 63037 2839 63095 2845
rect 63037 2836 63049 2839
rect 62540 2808 63049 2836
rect 62540 2796 62546 2808
rect 63037 2805 63049 2808
rect 63083 2805 63095 2839
rect 63144 2836 63172 2944
rect 64414 2932 64420 2984
rect 64472 2972 64478 2984
rect 64509 2975 64567 2981
rect 64509 2972 64521 2975
rect 64472 2944 64521 2972
rect 64472 2932 64478 2944
rect 64509 2941 64521 2944
rect 64555 2941 64567 2975
rect 70366 2972 70394 3012
rect 71590 3000 71596 3012
rect 71648 3000 71654 3052
rect 72160 3049 72188 3080
rect 76742 3068 76748 3080
rect 76800 3068 76806 3120
rect 77110 3108 77116 3120
rect 77071 3080 77116 3108
rect 77110 3068 77116 3080
rect 77168 3108 77174 3120
rect 79686 3108 79692 3120
rect 77168 3080 79692 3108
rect 77168 3068 77174 3080
rect 77680 3049 77708 3080
rect 79686 3068 79692 3080
rect 79744 3068 79750 3120
rect 72145 3043 72203 3049
rect 72145 3009 72157 3043
rect 72191 3009 72203 3043
rect 77665 3043 77723 3049
rect 72145 3003 72203 3009
rect 75196 3012 77616 3040
rect 75196 2972 75224 3012
rect 70366 2944 75224 2972
rect 64509 2935 64567 2941
rect 76742 2932 76748 2984
rect 76800 2972 76806 2984
rect 77481 2975 77539 2981
rect 77481 2972 77493 2975
rect 76800 2944 77493 2972
rect 76800 2932 76806 2944
rect 77481 2941 77493 2944
rect 77527 2941 77539 2975
rect 77588 2972 77616 3012
rect 77665 3009 77677 3043
rect 77711 3009 77723 3043
rect 77665 3003 77723 3009
rect 77849 3043 77907 3049
rect 77849 3009 77861 3043
rect 77895 3040 77907 3043
rect 78677 3043 78735 3049
rect 78677 3040 78689 3043
rect 77895 3012 78689 3040
rect 77895 3009 77907 3012
rect 77849 3003 77907 3009
rect 78677 3009 78689 3012
rect 78723 3009 78735 3043
rect 81526 3040 81532 3052
rect 81487 3012 81532 3040
rect 78677 3003 78735 3009
rect 81526 3000 81532 3012
rect 81584 3040 81590 3052
rect 82081 3043 82139 3049
rect 82081 3040 82093 3043
rect 81584 3012 82093 3040
rect 81584 3000 81590 3012
rect 82081 3009 82093 3012
rect 82127 3009 82139 3043
rect 84166 3040 84194 3148
rect 85945 3145 85957 3179
rect 85991 3145 86003 3179
rect 85945 3139 86003 3145
rect 86773 3179 86831 3185
rect 86773 3145 86785 3179
rect 86819 3176 86831 3179
rect 87690 3176 87696 3188
rect 86819 3148 87696 3176
rect 86819 3145 86831 3148
rect 86773 3139 86831 3145
rect 85960 3108 85988 3139
rect 87690 3136 87696 3148
rect 87748 3136 87754 3188
rect 87782 3136 87788 3188
rect 87840 3176 87846 3188
rect 88153 3179 88211 3185
rect 88153 3176 88165 3179
rect 87840 3148 88165 3176
rect 87840 3136 87846 3148
rect 88153 3145 88165 3148
rect 88199 3145 88211 3179
rect 88334 3176 88340 3188
rect 88295 3148 88340 3176
rect 88153 3139 88211 3145
rect 88334 3136 88340 3148
rect 88392 3136 88398 3188
rect 85960 3080 87552 3108
rect 87524 3049 87552 3080
rect 86129 3043 86187 3049
rect 86129 3040 86141 3043
rect 84166 3012 86141 3040
rect 82081 3003 82139 3009
rect 86129 3009 86141 3012
rect 86175 3009 86187 3043
rect 86957 3043 87015 3049
rect 86957 3040 86969 3043
rect 86129 3003 86187 3009
rect 86236 3012 86969 3040
rect 85022 2972 85028 2984
rect 77588 2944 85028 2972
rect 77481 2935 77539 2941
rect 85022 2932 85028 2944
rect 85080 2932 85086 2984
rect 85114 2932 85120 2984
rect 85172 2972 85178 2984
rect 86236 2972 86264 3012
rect 86957 3009 86969 3012
rect 87003 3009 87015 3043
rect 86957 3003 87015 3009
rect 87509 3043 87567 3049
rect 87509 3009 87521 3043
rect 87555 3009 87567 3043
rect 87509 3003 87567 3009
rect 88061 3043 88119 3049
rect 88061 3009 88073 3043
rect 88107 3009 88119 3043
rect 88061 3003 88119 3009
rect 88521 3043 88579 3049
rect 88521 3009 88533 3043
rect 88567 3040 88579 3043
rect 88904 3040 88932 3352
rect 88567 3012 88932 3040
rect 88567 3009 88579 3012
rect 88521 3003 88579 3009
rect 85172 2944 86264 2972
rect 85172 2932 85178 2944
rect 86862 2932 86868 2984
rect 86920 2972 86926 2984
rect 88076 2972 88104 3003
rect 86920 2944 88104 2972
rect 86920 2932 86926 2944
rect 63681 2907 63739 2913
rect 63681 2873 63693 2907
rect 63727 2904 63739 2907
rect 85482 2904 85488 2916
rect 63727 2876 85488 2904
rect 63727 2873 63739 2876
rect 63681 2867 63739 2873
rect 85482 2864 85488 2876
rect 85540 2864 85546 2916
rect 67450 2836 67456 2848
rect 63144 2808 67456 2836
rect 63037 2799 63095 2805
rect 67450 2796 67456 2808
rect 67508 2796 67514 2848
rect 68370 2796 68376 2848
rect 68428 2836 68434 2848
rect 68557 2839 68615 2845
rect 68557 2836 68569 2839
rect 68428 2808 68569 2836
rect 68428 2796 68434 2808
rect 68557 2805 68569 2808
rect 68603 2805 68615 2839
rect 68557 2799 68615 2805
rect 71498 2796 71504 2848
rect 71556 2836 71562 2848
rect 71961 2839 72019 2845
rect 71961 2836 71973 2839
rect 71556 2808 71973 2836
rect 71556 2796 71562 2808
rect 71961 2805 71973 2808
rect 72007 2805 72019 2839
rect 71961 2799 72019 2805
rect 78493 2839 78551 2845
rect 78493 2805 78505 2839
rect 78539 2836 78551 2839
rect 79962 2836 79968 2848
rect 78539 2808 79968 2836
rect 78539 2805 78551 2808
rect 78493 2799 78551 2805
rect 79962 2796 79968 2808
rect 80020 2796 80026 2848
rect 81802 2796 81808 2848
rect 81860 2836 81866 2848
rect 81897 2839 81955 2845
rect 81897 2836 81909 2839
rect 81860 2808 81909 2836
rect 81860 2796 81866 2808
rect 81897 2805 81909 2808
rect 81943 2805 81955 2839
rect 81897 2799 81955 2805
rect 86954 2796 86960 2848
rect 87012 2836 87018 2848
rect 87325 2839 87383 2845
rect 87325 2836 87337 2839
rect 87012 2808 87337 2836
rect 87012 2796 87018 2808
rect 87325 2805 87337 2808
rect 87371 2805 87383 2839
rect 87325 2799 87383 2805
rect 1104 2746 88872 2768
rect 1104 2694 11924 2746
rect 11976 2694 11988 2746
rect 12040 2694 12052 2746
rect 12104 2694 12116 2746
rect 12168 2694 12180 2746
rect 12232 2694 33872 2746
rect 33924 2694 33936 2746
rect 33988 2694 34000 2746
rect 34052 2694 34064 2746
rect 34116 2694 34128 2746
rect 34180 2694 55820 2746
rect 55872 2694 55884 2746
rect 55936 2694 55948 2746
rect 56000 2694 56012 2746
rect 56064 2694 56076 2746
rect 56128 2694 77768 2746
rect 77820 2694 77832 2746
rect 77884 2694 77896 2746
rect 77948 2694 77960 2746
rect 78012 2694 78024 2746
rect 78076 2694 88872 2746
rect 1104 2672 88872 2694
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 11747 2604 27752 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 4154 2524 4160 2576
rect 4212 2564 4218 2576
rect 4709 2567 4767 2573
rect 4709 2564 4721 2567
rect 4212 2536 4721 2564
rect 4212 2524 4218 2536
rect 4709 2533 4721 2536
rect 4755 2533 4767 2567
rect 21174 2564 21180 2576
rect 4709 2527 4767 2533
rect 6886 2536 21180 2564
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2496 6699 2499
rect 6886 2496 6914 2536
rect 21174 2524 21180 2536
rect 21232 2524 21238 2576
rect 23290 2524 23296 2576
rect 23348 2564 23354 2576
rect 24029 2567 24087 2573
rect 24029 2564 24041 2567
rect 23348 2536 24041 2564
rect 23348 2524 23354 2536
rect 24029 2533 24041 2536
rect 24075 2533 24087 2567
rect 24029 2527 24087 2533
rect 25225 2567 25283 2573
rect 25225 2533 25237 2567
rect 25271 2564 25283 2567
rect 26418 2564 26424 2576
rect 25271 2536 26424 2564
rect 25271 2533 25283 2536
rect 25225 2527 25283 2533
rect 26418 2524 26424 2536
rect 26476 2524 26482 2576
rect 26510 2524 26516 2576
rect 26568 2564 26574 2576
rect 27246 2564 27252 2576
rect 26568 2536 27252 2564
rect 26568 2524 26574 2536
rect 27246 2524 27252 2536
rect 27304 2524 27310 2576
rect 27341 2567 27399 2573
rect 27341 2533 27353 2567
rect 27387 2564 27399 2567
rect 27522 2564 27528 2576
rect 27387 2536 27528 2564
rect 27387 2533 27399 2536
rect 27341 2527 27399 2533
rect 27522 2524 27528 2536
rect 27580 2524 27586 2576
rect 10226 2496 10232 2508
rect 6687 2468 6914 2496
rect 8496 2468 10232 2496
rect 6687 2465 6699 2468
rect 6641 2459 6699 2465
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 2777 2431 2835 2437
rect 2777 2428 2789 2431
rect 2363 2400 2789 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2777 2397 2789 2400
rect 2823 2428 2835 2431
rect 2866 2428 2872 2440
rect 2823 2400 2872 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3326 2428 3332 2440
rect 3287 2400 3332 2428
rect 3326 2388 3332 2400
rect 3384 2388 3390 2440
rect 4890 2428 4896 2440
rect 4851 2400 4896 2428
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5534 2428 5540 2440
rect 5491 2400 5540 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5868 2400 6377 2428
rect 5868 2388 5874 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8496 2437 8524 2468
rect 10226 2456 10232 2468
rect 10284 2456 10290 2508
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 15838 2496 15844 2508
rect 13127 2468 15844 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 15838 2456 15844 2468
rect 15896 2456 15902 2508
rect 18690 2456 18696 2508
rect 18748 2496 18754 2508
rect 19245 2499 19303 2505
rect 19245 2496 19257 2499
rect 18748 2468 19257 2496
rect 18748 2456 18754 2468
rect 19245 2465 19257 2468
rect 19291 2465 19303 2499
rect 20162 2496 20168 2508
rect 19245 2459 19303 2465
rect 19444 2468 20168 2496
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7800 2400 7941 2428
rect 7800 2388 7806 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9766 2428 9772 2440
rect 9355 2400 9772 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 9950 2428 9956 2440
rect 9911 2400 9956 2428
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10502 2428 10508 2440
rect 10463 2400 10508 2428
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2428 11115 2431
rect 12161 2431 12219 2437
rect 11103 2400 12112 2428
rect 11103 2397 11115 2400
rect 11057 2391 11115 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1581 2363 1639 2369
rect 1581 2360 1593 2363
rect 1360 2332 1593 2360
rect 1360 2320 1366 2332
rect 1581 2329 1593 2332
rect 1627 2329 1639 2363
rect 1581 2323 1639 2329
rect 1949 2363 2007 2369
rect 1949 2329 1961 2363
rect 1995 2360 2007 2363
rect 2682 2360 2688 2372
rect 1995 2332 2688 2360
rect 1995 2329 2007 2332
rect 1949 2323 2007 2329
rect 2682 2320 2688 2332
rect 2740 2320 2746 2372
rect 3878 2320 3884 2372
rect 3936 2360 3942 2372
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 3936 2332 4169 2360
rect 3936 2320 3942 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 11606 2360 11612 2372
rect 11567 2332 11612 2360
rect 4157 2323 4215 2329
rect 11606 2320 11612 2332
rect 11664 2320 11670 2372
rect 12084 2360 12112 2400
rect 12161 2397 12173 2431
rect 12207 2428 12219 2431
rect 12250 2428 12256 2440
rect 12207 2400 12256 2428
rect 12207 2397 12219 2400
rect 12161 2391 12219 2397
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2428 12863 2431
rect 12894 2428 12900 2440
rect 12851 2400 12900 2428
rect 12851 2397 12863 2400
rect 12805 2391 12863 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2428 14151 2431
rect 14182 2428 14188 2440
rect 14139 2400 14188 2428
rect 14139 2397 14151 2400
rect 14093 2391 14151 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 14366 2428 14372 2440
rect 14327 2400 14372 2428
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15746 2428 15752 2440
rect 15335 2400 15752 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16172 2400 16681 2428
rect 16172 2388 16178 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16942 2428 16948 2440
rect 16903 2400 16948 2428
rect 16669 2391 16727 2397
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18233 2431 18291 2437
rect 18233 2428 18245 2431
rect 18104 2400 18245 2428
rect 18104 2388 18110 2400
rect 18233 2397 18245 2400
rect 18279 2397 18291 2431
rect 18233 2391 18291 2397
rect 18785 2431 18843 2437
rect 18785 2397 18797 2431
rect 18831 2428 18843 2431
rect 19444 2428 19472 2468
rect 20162 2456 20168 2468
rect 20220 2456 20226 2508
rect 22830 2496 22836 2508
rect 21376 2468 22836 2496
rect 18831 2400 19472 2428
rect 19521 2431 19579 2437
rect 18831 2397 18843 2400
rect 18785 2391 18843 2397
rect 19521 2397 19533 2431
rect 19567 2397 19579 2431
rect 20806 2428 20812 2440
rect 20767 2400 20812 2428
rect 19521 2391 19579 2397
rect 15378 2360 15384 2372
rect 12084 2332 15384 2360
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 19536 2360 19564 2391
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 21376 2437 21404 2468
rect 22830 2456 22836 2468
rect 22888 2456 22894 2508
rect 27614 2496 27620 2508
rect 26896 2468 27620 2496
rect 21361 2431 21419 2437
rect 21361 2397 21373 2431
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21968 2400 22017 2428
rect 21968 2388 21974 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2428 23535 2431
rect 23934 2428 23940 2440
rect 23523 2400 23940 2428
rect 23523 2397 23535 2400
rect 23477 2391 23535 2397
rect 23934 2388 23940 2400
rect 23992 2388 23998 2440
rect 24210 2428 24216 2440
rect 24171 2400 24216 2428
rect 24210 2388 24216 2400
rect 24268 2388 24274 2440
rect 24762 2428 24768 2440
rect 24723 2400 24768 2428
rect 24762 2388 24768 2400
rect 24820 2388 24826 2440
rect 25406 2428 25412 2440
rect 25367 2400 25412 2428
rect 25406 2388 25412 2400
rect 25464 2388 25470 2440
rect 26053 2431 26111 2437
rect 26053 2397 26065 2431
rect 26099 2428 26111 2431
rect 26510 2428 26516 2440
rect 26099 2400 26516 2428
rect 26099 2397 26111 2400
rect 26053 2391 26111 2397
rect 26510 2388 26516 2400
rect 26568 2388 26574 2440
rect 26789 2431 26847 2437
rect 26789 2397 26801 2431
rect 26835 2428 26847 2431
rect 26896 2428 26924 2468
rect 27614 2456 27620 2468
rect 27672 2456 27678 2508
rect 27724 2496 27752 2604
rect 27798 2592 27804 2644
rect 27856 2632 27862 2644
rect 27893 2635 27951 2641
rect 27893 2632 27905 2635
rect 27856 2604 27905 2632
rect 27856 2592 27862 2604
rect 27893 2601 27905 2604
rect 27939 2601 27951 2635
rect 27893 2595 27951 2601
rect 29914 2592 29920 2644
rect 29972 2632 29978 2644
rect 30374 2632 30380 2644
rect 29972 2604 30380 2632
rect 29972 2592 29978 2604
rect 30374 2592 30380 2604
rect 30432 2592 30438 2644
rect 31110 2592 31116 2644
rect 31168 2632 31174 2644
rect 45462 2632 45468 2644
rect 31168 2604 45468 2632
rect 31168 2592 31174 2604
rect 45462 2592 45468 2604
rect 45520 2592 45526 2644
rect 46290 2592 46296 2644
rect 46348 2632 46354 2644
rect 48685 2635 48743 2641
rect 48685 2632 48697 2635
rect 46348 2604 48697 2632
rect 46348 2592 46354 2604
rect 48685 2601 48697 2604
rect 48731 2601 48743 2635
rect 48685 2595 48743 2601
rect 49970 2592 49976 2644
rect 50028 2632 50034 2644
rect 50157 2635 50215 2641
rect 50157 2632 50169 2635
rect 50028 2604 50169 2632
rect 50028 2592 50034 2604
rect 50157 2601 50169 2604
rect 50203 2601 50215 2635
rect 50157 2595 50215 2601
rect 50246 2592 50252 2644
rect 50304 2632 50310 2644
rect 51905 2635 51963 2641
rect 51905 2632 51917 2635
rect 50304 2604 51917 2632
rect 50304 2592 50310 2604
rect 51905 2601 51917 2604
rect 51951 2601 51963 2635
rect 51905 2595 51963 2601
rect 53282 2592 53288 2644
rect 53340 2632 53346 2644
rect 55309 2635 55367 2641
rect 55309 2632 55321 2635
rect 53340 2604 55321 2632
rect 53340 2592 53346 2604
rect 55309 2601 55321 2604
rect 55355 2601 55367 2635
rect 55309 2595 55367 2601
rect 55582 2592 55588 2644
rect 55640 2632 55646 2644
rect 55861 2635 55919 2641
rect 55861 2632 55873 2635
rect 55640 2604 55873 2632
rect 55640 2592 55646 2604
rect 55861 2601 55873 2604
rect 55907 2601 55919 2635
rect 55861 2595 55919 2601
rect 59262 2592 59268 2644
rect 59320 2632 59326 2644
rect 60461 2635 60519 2641
rect 60461 2632 60473 2635
rect 59320 2604 60473 2632
rect 59320 2592 59326 2604
rect 60461 2601 60473 2604
rect 60507 2601 60519 2635
rect 61286 2632 61292 2644
rect 61247 2604 61292 2632
rect 60461 2595 60519 2601
rect 61286 2592 61292 2604
rect 61344 2592 61350 2644
rect 63678 2592 63684 2644
rect 63736 2632 63742 2644
rect 69014 2632 69020 2644
rect 63736 2604 68876 2632
rect 68975 2604 69020 2632
rect 63736 2592 63742 2604
rect 31662 2564 31668 2576
rect 28552 2536 31668 2564
rect 28552 2505 28580 2536
rect 31662 2524 31668 2536
rect 31720 2524 31726 2576
rect 31846 2524 31852 2576
rect 31904 2564 31910 2576
rect 31904 2536 34836 2564
rect 31904 2524 31910 2536
rect 28537 2499 28595 2505
rect 27724 2468 28028 2496
rect 26835 2400 26924 2428
rect 27525 2431 27583 2437
rect 26835 2397 26847 2400
rect 26789 2391 26847 2397
rect 27525 2397 27537 2431
rect 27571 2428 27583 2431
rect 27890 2428 27896 2440
rect 27571 2400 27896 2428
rect 27571 2397 27583 2400
rect 27525 2391 27583 2397
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 28000 2428 28028 2468
rect 28537 2465 28549 2499
rect 28583 2465 28595 2499
rect 31570 2496 31576 2508
rect 28537 2459 28595 2465
rect 28644 2468 31576 2496
rect 28644 2428 28672 2468
rect 31570 2456 31576 2468
rect 31628 2456 31634 2508
rect 34808 2496 34836 2536
rect 34882 2524 34888 2576
rect 34940 2564 34946 2576
rect 38746 2564 38752 2576
rect 34940 2536 38752 2564
rect 34940 2524 34946 2536
rect 38746 2524 38752 2536
rect 38804 2524 38810 2576
rect 38930 2524 38936 2576
rect 38988 2564 38994 2576
rect 38988 2536 40632 2564
rect 38988 2524 38994 2536
rect 34808 2468 36308 2496
rect 29914 2428 29920 2440
rect 28000 2400 28672 2428
rect 29875 2400 29920 2428
rect 29914 2388 29920 2400
rect 29972 2388 29978 2440
rect 30469 2431 30527 2437
rect 30469 2397 30481 2431
rect 30515 2397 30527 2431
rect 30469 2391 30527 2397
rect 26142 2360 26148 2372
rect 19536 2332 26148 2360
rect 26142 2320 26148 2332
rect 26200 2320 26206 2372
rect 26970 2360 26976 2372
rect 26344 2332 26976 2360
rect 2590 2292 2596 2304
rect 2551 2264 2596 2292
rect 2590 2252 2596 2264
rect 2648 2252 2654 2304
rect 3145 2295 3203 2301
rect 3145 2261 3157 2295
rect 3191 2292 3203 2295
rect 3234 2292 3240 2304
rect 3191 2264 3240 2292
rect 3191 2261 3203 2264
rect 3145 2255 3203 2261
rect 3234 2252 3240 2264
rect 3292 2252 3298 2304
rect 4246 2292 4252 2304
rect 4207 2264 4252 2292
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5261 2295 5319 2301
rect 5261 2292 5273 2295
rect 5224 2264 5273 2292
rect 5224 2252 5230 2264
rect 5261 2261 5273 2264
rect 5307 2261 5319 2295
rect 5261 2255 5319 2261
rect 7745 2295 7803 2301
rect 7745 2261 7757 2295
rect 7791 2292 7803 2295
rect 8202 2292 8208 2304
rect 7791 2264 8208 2292
rect 7791 2261 7803 2264
rect 7745 2255 7803 2261
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 8297 2295 8355 2301
rect 8297 2261 8309 2295
rect 8343 2292 8355 2295
rect 8386 2292 8392 2304
rect 8343 2264 8392 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 9088 2264 9137 2292
rect 9088 2252 9094 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9732 2264 9781 2292
rect 9732 2252 9738 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 10318 2292 10324 2304
rect 10279 2264 10324 2292
rect 9769 2255 9827 2261
rect 10318 2252 10324 2264
rect 10376 2252 10382 2304
rect 10873 2295 10931 2301
rect 10873 2261 10885 2295
rect 10919 2292 10931 2295
rect 10962 2292 10968 2304
rect 10919 2264 10968 2292
rect 10919 2261 10931 2264
rect 10873 2255 10931 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 12342 2292 12348 2304
rect 12303 2264 12348 2292
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15565 2295 15623 2301
rect 15565 2292 15577 2295
rect 15528 2264 15577 2292
rect 15528 2252 15534 2264
rect 15565 2261 15577 2264
rect 15611 2261 15623 2295
rect 15565 2255 15623 2261
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 19334 2292 19340 2304
rect 18647 2264 19340 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 19334 2252 19340 2264
rect 19392 2252 19398 2304
rect 20622 2292 20628 2304
rect 20583 2264 20628 2292
rect 20622 2252 20628 2264
rect 20680 2252 20686 2304
rect 21177 2295 21235 2301
rect 21177 2261 21189 2295
rect 21223 2292 21235 2295
rect 21266 2292 21272 2304
rect 21223 2264 21272 2292
rect 21223 2261 21235 2264
rect 21177 2255 21235 2261
rect 21266 2252 21272 2264
rect 21324 2252 21330 2304
rect 22186 2292 22192 2304
rect 22147 2264 22192 2292
rect 22186 2252 22192 2264
rect 22244 2252 22250 2304
rect 23753 2295 23811 2301
rect 23753 2261 23765 2295
rect 23799 2292 23811 2295
rect 23842 2292 23848 2304
rect 23799 2264 23848 2292
rect 23799 2261 23811 2264
rect 23753 2255 23811 2261
rect 23842 2252 23848 2264
rect 23900 2252 23906 2304
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24394 2292 24400 2304
rect 24084 2264 24400 2292
rect 24084 2252 24090 2264
rect 24394 2252 24400 2264
rect 24452 2252 24458 2304
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 26344 2301 26372 2332
rect 26970 2320 26976 2332
rect 27028 2320 27034 2372
rect 27798 2320 27804 2372
rect 27856 2360 27862 2372
rect 28353 2363 28411 2369
rect 28353 2360 28365 2363
rect 27856 2332 28365 2360
rect 27856 2320 27862 2332
rect 28353 2329 28365 2332
rect 28399 2329 28411 2363
rect 28353 2323 28411 2329
rect 28994 2320 29000 2372
rect 29052 2360 29058 2372
rect 30484 2360 30512 2391
rect 31478 2388 31484 2440
rect 31536 2428 31542 2440
rect 31657 2431 31715 2437
rect 31657 2428 31669 2431
rect 31536 2400 31669 2428
rect 31536 2388 31542 2400
rect 31657 2397 31669 2400
rect 31703 2397 31715 2431
rect 31657 2391 31715 2397
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32916 2400 32965 2428
rect 32916 2388 32922 2400
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 33229 2431 33287 2437
rect 33229 2397 33241 2431
rect 33275 2428 33287 2431
rect 34790 2428 34796 2440
rect 33275 2400 34796 2428
rect 33275 2397 33287 2400
rect 33229 2391 33287 2397
rect 34790 2388 34796 2400
rect 34848 2388 34854 2440
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2428 34943 2431
rect 35342 2428 35348 2440
rect 34931 2400 35348 2428
rect 34931 2397 34943 2400
rect 34885 2391 34943 2397
rect 35342 2388 35348 2400
rect 35400 2388 35406 2440
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 36280 2437 36308 2468
rect 36354 2456 36360 2508
rect 36412 2496 36418 2508
rect 36412 2468 38654 2496
rect 36412 2456 36418 2468
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 36265 2431 36323 2437
rect 36265 2397 36277 2431
rect 36311 2397 36323 2431
rect 36814 2428 36820 2440
rect 36775 2400 36820 2428
rect 36265 2391 36323 2397
rect 36814 2388 36820 2400
rect 36872 2388 36878 2440
rect 37642 2428 37648 2440
rect 37603 2400 37648 2428
rect 37642 2388 37648 2400
rect 37700 2388 37706 2440
rect 38626 2424 38654 2468
rect 39758 2456 39764 2508
rect 39816 2496 39822 2508
rect 40129 2499 40187 2505
rect 39816 2468 39988 2496
rect 39816 2456 39822 2468
rect 38746 2424 38752 2440
rect 38626 2396 38752 2424
rect 38746 2388 38752 2396
rect 38804 2388 38810 2440
rect 38933 2407 38991 2413
rect 38933 2373 38945 2407
rect 38979 2404 38991 2407
rect 38979 2376 39068 2404
rect 39298 2388 39304 2440
rect 39356 2428 39362 2440
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 39356 2400 39865 2428
rect 39356 2388 39362 2400
rect 39853 2397 39865 2400
rect 39899 2397 39911 2431
rect 39960 2428 39988 2468
rect 40129 2465 40141 2499
rect 40175 2496 40187 2499
rect 40494 2496 40500 2508
rect 40175 2468 40500 2496
rect 40175 2465 40187 2468
rect 40129 2459 40187 2465
rect 40494 2456 40500 2468
rect 40552 2456 40558 2508
rect 40604 2496 40632 2536
rect 43714 2524 43720 2576
rect 43772 2564 43778 2576
rect 44361 2567 44419 2573
rect 44361 2564 44373 2567
rect 43772 2536 44373 2564
rect 43772 2524 43778 2536
rect 44361 2533 44373 2536
rect 44407 2533 44419 2567
rect 44361 2527 44419 2533
rect 45189 2567 45247 2573
rect 45189 2533 45201 2567
rect 45235 2533 45247 2567
rect 45189 2527 45247 2533
rect 45204 2496 45232 2527
rect 45278 2524 45284 2576
rect 45336 2564 45342 2576
rect 45336 2536 68692 2564
rect 45336 2524 45342 2536
rect 46842 2496 46848 2508
rect 40604 2468 44128 2496
rect 45204 2468 46848 2496
rect 41233 2431 41291 2437
rect 41233 2428 41245 2431
rect 39960 2400 41245 2428
rect 39853 2391 39911 2397
rect 41233 2397 41245 2400
rect 41279 2397 41291 2431
rect 41966 2428 41972 2440
rect 41927 2400 41972 2428
rect 41233 2391 41291 2397
rect 41966 2388 41972 2400
rect 42024 2388 42030 2440
rect 42794 2428 42800 2440
rect 42755 2400 42800 2428
rect 42794 2388 42800 2400
rect 42852 2388 42858 2440
rect 43438 2428 43444 2440
rect 43399 2400 43444 2428
rect 43438 2388 43444 2400
rect 43496 2388 43502 2440
rect 43993 2431 44051 2437
rect 43993 2397 44005 2431
rect 44039 2397 44051 2431
rect 43993 2391 44051 2397
rect 38979 2373 38991 2376
rect 31110 2360 31116 2372
rect 29052 2332 30328 2360
rect 30484 2332 31116 2360
rect 29052 2320 29058 2332
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24544 2264 24593 2292
rect 24544 2252 24550 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 26329 2295 26387 2301
rect 26329 2261 26341 2295
rect 26375 2261 26387 2295
rect 26329 2255 26387 2261
rect 26605 2295 26663 2301
rect 26605 2261 26617 2295
rect 26651 2292 26663 2295
rect 27062 2292 27068 2304
rect 26651 2264 27068 2292
rect 26651 2261 26663 2264
rect 26605 2255 26663 2261
rect 27062 2252 27068 2264
rect 27120 2252 27126 2304
rect 28258 2292 28264 2304
rect 28219 2264 28264 2292
rect 28258 2252 28264 2264
rect 28316 2292 28322 2304
rect 29178 2292 29184 2304
rect 28316 2264 29184 2292
rect 28316 2252 28322 2264
rect 29178 2252 29184 2264
rect 29236 2252 29242 2304
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 30300 2301 30328 2332
rect 31110 2320 31116 2332
rect 31168 2320 31174 2372
rect 31294 2320 31300 2372
rect 31352 2360 31358 2372
rect 32401 2363 32459 2369
rect 32401 2360 32413 2363
rect 31352 2332 32413 2360
rect 31352 2320 31358 2332
rect 32401 2329 32413 2332
rect 32447 2329 32459 2363
rect 32401 2323 32459 2329
rect 32674 2320 32680 2372
rect 32732 2360 32738 2372
rect 38933 2367 38991 2373
rect 39040 2360 39068 2376
rect 39114 2360 39120 2372
rect 32732 2332 37596 2360
rect 39040 2332 39120 2360
rect 32732 2320 32738 2332
rect 29733 2295 29791 2301
rect 29733 2292 29745 2295
rect 29696 2264 29745 2292
rect 29696 2252 29702 2264
rect 29733 2261 29745 2264
rect 29779 2261 29791 2295
rect 29733 2255 29791 2261
rect 30285 2295 30343 2301
rect 30285 2261 30297 2295
rect 30331 2261 30343 2295
rect 30285 2255 30343 2261
rect 31481 2295 31539 2301
rect 31481 2261 31493 2295
rect 31527 2292 31539 2295
rect 32214 2292 32220 2304
rect 31527 2264 32220 2292
rect 31527 2261 31539 2264
rect 31481 2255 31539 2261
rect 32214 2252 32220 2264
rect 32272 2252 32278 2304
rect 32493 2295 32551 2301
rect 32493 2261 32505 2295
rect 32539 2292 32551 2295
rect 34054 2292 34060 2304
rect 32539 2264 34060 2292
rect 32539 2261 32551 2264
rect 32493 2255 32551 2261
rect 34054 2252 34060 2264
rect 34112 2252 34118 2304
rect 34146 2252 34152 2304
rect 34204 2292 34210 2304
rect 34701 2295 34759 2301
rect 34701 2292 34713 2295
rect 34204 2264 34713 2292
rect 34204 2252 34210 2264
rect 34701 2261 34713 2264
rect 34747 2261 34759 2295
rect 36078 2292 36084 2304
rect 36039 2264 36084 2292
rect 34701 2255 34759 2261
rect 36078 2252 36084 2264
rect 36136 2252 36142 2304
rect 36633 2295 36691 2301
rect 36633 2261 36645 2295
rect 36679 2292 36691 2295
rect 36722 2292 36728 2304
rect 36679 2264 36728 2292
rect 36679 2261 36691 2264
rect 36633 2255 36691 2261
rect 36722 2252 36728 2264
rect 36780 2252 36786 2304
rect 37366 2252 37372 2304
rect 37424 2292 37430 2304
rect 37461 2295 37519 2301
rect 37461 2292 37473 2295
rect 37424 2264 37473 2292
rect 37424 2252 37430 2264
rect 37461 2261 37473 2264
rect 37507 2261 37519 2295
rect 37568 2292 37596 2332
rect 39114 2320 39120 2332
rect 39172 2320 39178 2372
rect 41690 2320 41696 2372
rect 41748 2360 41754 2372
rect 44008 2360 44036 2391
rect 41748 2332 44036 2360
rect 44100 2360 44128 2468
rect 46842 2456 46848 2468
rect 46900 2456 46906 2508
rect 50706 2496 50712 2508
rect 46952 2468 49740 2496
rect 50667 2468 50712 2496
rect 44450 2388 44456 2440
rect 44508 2428 44514 2440
rect 44545 2431 44603 2437
rect 44545 2428 44557 2431
rect 44508 2400 44557 2428
rect 44508 2388 44514 2400
rect 44545 2397 44557 2400
rect 44591 2397 44603 2431
rect 44545 2391 44603 2397
rect 45186 2388 45192 2440
rect 45244 2428 45250 2440
rect 45373 2431 45431 2437
rect 45373 2428 45385 2431
rect 45244 2400 45385 2428
rect 45244 2388 45250 2400
rect 45373 2397 45385 2400
rect 45419 2397 45431 2431
rect 45373 2391 45431 2397
rect 46293 2431 46351 2437
rect 46293 2397 46305 2431
rect 46339 2428 46351 2431
rect 46382 2428 46388 2440
rect 46339 2400 46388 2428
rect 46339 2397 46351 2400
rect 46293 2391 46351 2397
rect 46382 2388 46388 2400
rect 46440 2388 46446 2440
rect 46569 2431 46627 2437
rect 46569 2397 46581 2431
rect 46615 2428 46627 2431
rect 46750 2428 46756 2440
rect 46615 2400 46756 2428
rect 46615 2397 46627 2400
rect 46569 2391 46627 2397
rect 46750 2388 46756 2400
rect 46808 2388 46814 2440
rect 46952 2360 46980 2468
rect 47026 2388 47032 2440
rect 47084 2428 47090 2440
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 47084 2400 47777 2428
rect 47084 2388 47090 2400
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 48222 2388 48228 2440
rect 48280 2424 48286 2440
rect 48317 2431 48375 2437
rect 48317 2424 48329 2431
rect 48280 2397 48329 2424
rect 48363 2397 48375 2431
rect 48280 2396 48375 2397
rect 48280 2388 48286 2396
rect 48317 2391 48375 2396
rect 48406 2388 48412 2440
rect 48464 2428 48470 2440
rect 48869 2431 48927 2437
rect 48869 2428 48881 2431
rect 48464 2400 48881 2428
rect 48464 2388 48470 2400
rect 48869 2397 48881 2400
rect 48915 2397 48927 2431
rect 48869 2391 48927 2397
rect 49513 2431 49571 2437
rect 49513 2397 49525 2431
rect 49559 2428 49571 2431
rect 49602 2428 49608 2440
rect 49559 2400 49608 2428
rect 49559 2397 49571 2400
rect 49513 2391 49571 2397
rect 49602 2388 49608 2400
rect 49660 2388 49666 2440
rect 49712 2428 49740 2468
rect 50706 2456 50712 2468
rect 50764 2456 50770 2508
rect 50982 2456 50988 2508
rect 51040 2496 51046 2508
rect 51040 2468 62160 2496
rect 51040 2456 51046 2468
rect 52089 2431 52147 2437
rect 52089 2428 52101 2431
rect 49712 2400 52101 2428
rect 52089 2397 52101 2400
rect 52135 2397 52147 2431
rect 54386 2428 54392 2440
rect 54347 2400 54392 2428
rect 52089 2391 52147 2397
rect 54386 2388 54392 2400
rect 54444 2388 54450 2440
rect 54754 2388 54760 2440
rect 54812 2428 54818 2440
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 54812 2400 55505 2428
rect 54812 2388 54818 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 55493 2391 55551 2397
rect 56045 2431 56103 2437
rect 56045 2397 56057 2431
rect 56091 2397 56103 2431
rect 56594 2428 56600 2440
rect 56555 2400 56600 2428
rect 56045 2391 56103 2397
rect 44100 2332 46980 2360
rect 41748 2320 41754 2332
rect 47854 2320 47860 2372
rect 47912 2360 47918 2372
rect 47912 2332 48176 2360
rect 47912 2320 47918 2332
rect 38654 2292 38660 2304
rect 37568 2264 38660 2292
rect 37461 2255 37519 2261
rect 38654 2252 38660 2264
rect 38712 2252 38718 2304
rect 38746 2252 38752 2304
rect 38804 2292 38810 2304
rect 38804 2264 38849 2292
rect 38804 2252 38810 2264
rect 40586 2252 40592 2304
rect 40644 2292 40650 2304
rect 41049 2295 41107 2301
rect 41049 2292 41061 2295
rect 40644 2264 41061 2292
rect 40644 2252 40650 2264
rect 41049 2261 41061 2264
rect 41095 2261 41107 2295
rect 41049 2255 41107 2261
rect 41785 2295 41843 2301
rect 41785 2261 41797 2295
rect 41831 2292 41843 2295
rect 41874 2292 41880 2304
rect 41831 2264 41880 2292
rect 41831 2261 41843 2264
rect 41785 2255 41843 2261
rect 41874 2252 41880 2264
rect 41932 2252 41938 2304
rect 42518 2252 42524 2304
rect 42576 2292 42582 2304
rect 42613 2295 42671 2301
rect 42613 2292 42625 2295
rect 42576 2264 42625 2292
rect 42576 2252 42582 2264
rect 42613 2261 42625 2264
rect 42659 2261 42671 2295
rect 42613 2255 42671 2261
rect 43162 2252 43168 2304
rect 43220 2292 43226 2304
rect 43257 2295 43315 2301
rect 43257 2292 43269 2295
rect 43220 2264 43269 2292
rect 43220 2252 43226 2264
rect 43257 2261 43269 2264
rect 43303 2261 43315 2295
rect 43806 2292 43812 2304
rect 43767 2264 43812 2292
rect 43257 2255 43315 2261
rect 43806 2252 43812 2264
rect 43864 2252 43870 2304
rect 45554 2252 45560 2304
rect 45612 2292 45618 2304
rect 48038 2292 48044 2304
rect 45612 2264 48044 2292
rect 45612 2252 45618 2264
rect 48038 2252 48044 2264
rect 48096 2252 48102 2304
rect 48148 2301 48176 2332
rect 48424 2332 50844 2360
rect 48133 2295 48191 2301
rect 48133 2261 48145 2295
rect 48179 2261 48191 2295
rect 48133 2255 48191 2261
rect 48222 2252 48228 2304
rect 48280 2292 48286 2304
rect 48424 2292 48452 2332
rect 48280 2264 48452 2292
rect 48280 2252 48286 2264
rect 48774 2252 48780 2304
rect 48832 2292 48838 2304
rect 49605 2295 49663 2301
rect 49605 2292 49617 2295
rect 48832 2264 49617 2292
rect 48832 2252 48838 2264
rect 49605 2261 49617 2264
rect 49651 2261 49663 2295
rect 49605 2255 49663 2261
rect 50338 2252 50344 2304
rect 50396 2292 50402 2304
rect 50525 2295 50583 2301
rect 50525 2292 50537 2295
rect 50396 2264 50537 2292
rect 50396 2252 50402 2264
rect 50525 2261 50537 2264
rect 50571 2261 50583 2295
rect 50525 2255 50583 2261
rect 50614 2252 50620 2304
rect 50672 2292 50678 2304
rect 50816 2292 50844 2332
rect 50890 2320 50896 2372
rect 50948 2360 50954 2372
rect 51353 2363 51411 2369
rect 51353 2360 51365 2363
rect 50948 2332 51365 2360
rect 50948 2320 50954 2332
rect 51353 2329 51365 2332
rect 51399 2329 51411 2363
rect 51353 2323 51411 2329
rect 52822 2320 52828 2372
rect 52880 2360 52886 2372
rect 53101 2363 53159 2369
rect 53101 2360 53113 2363
rect 52880 2332 53113 2360
rect 52880 2320 52886 2332
rect 53101 2329 53113 2332
rect 53147 2329 53159 2363
rect 53101 2323 53159 2329
rect 55398 2320 55404 2372
rect 55456 2360 55462 2372
rect 56060 2360 56088 2391
rect 56594 2388 56600 2400
rect 56652 2388 56658 2440
rect 57146 2428 57152 2440
rect 57107 2400 57152 2428
rect 57146 2388 57152 2400
rect 57204 2388 57210 2440
rect 57974 2388 57980 2440
rect 58032 2428 58038 2440
rect 58069 2431 58127 2437
rect 58069 2428 58081 2431
rect 58032 2400 58081 2428
rect 58032 2388 58038 2400
rect 58069 2397 58081 2400
rect 58115 2397 58127 2431
rect 58069 2391 58127 2397
rect 58342 2388 58348 2440
rect 58400 2428 58406 2440
rect 58621 2431 58679 2437
rect 58621 2428 58633 2431
rect 58400 2400 58633 2428
rect 58400 2388 58406 2400
rect 58621 2397 58633 2400
rect 58667 2397 58679 2431
rect 59170 2428 59176 2440
rect 59131 2400 59176 2428
rect 58621 2391 58679 2397
rect 59170 2388 59176 2400
rect 59228 2388 59234 2440
rect 59262 2388 59268 2440
rect 59320 2428 59326 2440
rect 59725 2431 59783 2437
rect 59725 2428 59737 2431
rect 59320 2400 59737 2428
rect 59320 2388 59326 2400
rect 59725 2397 59737 2400
rect 59771 2397 59783 2431
rect 59725 2391 59783 2397
rect 59906 2388 59912 2440
rect 59964 2428 59970 2440
rect 60645 2431 60703 2437
rect 60645 2428 60657 2431
rect 59964 2400 60657 2428
rect 59964 2388 59970 2400
rect 60645 2397 60657 2400
rect 60691 2397 60703 2431
rect 60645 2391 60703 2397
rect 61194 2388 61200 2440
rect 61252 2428 61258 2440
rect 62132 2437 62160 2468
rect 62206 2456 62212 2508
rect 62264 2496 62270 2508
rect 62264 2468 64874 2496
rect 62264 2456 62270 2468
rect 61473 2431 61531 2437
rect 61473 2428 61485 2431
rect 61252 2400 61485 2428
rect 61252 2388 61258 2400
rect 61473 2397 61485 2400
rect 61519 2397 61531 2431
rect 61473 2391 61531 2397
rect 62117 2431 62175 2437
rect 62117 2397 62129 2431
rect 62163 2397 62175 2431
rect 62117 2391 62175 2397
rect 63126 2388 63132 2440
rect 63184 2428 63190 2440
rect 63221 2431 63279 2437
rect 63221 2428 63233 2431
rect 63184 2400 63233 2428
rect 63184 2388 63190 2400
rect 63221 2397 63233 2400
rect 63267 2397 63279 2431
rect 63494 2428 63500 2440
rect 63455 2400 63500 2428
rect 63221 2391 63279 2397
rect 63494 2388 63500 2400
rect 63552 2388 63558 2440
rect 55456 2332 56088 2360
rect 64846 2360 64874 2468
rect 64966 2456 64972 2508
rect 65024 2496 65030 2508
rect 65024 2468 66392 2496
rect 65024 2456 65030 2468
rect 65797 2431 65855 2437
rect 65797 2397 65809 2431
rect 65843 2428 65855 2431
rect 66254 2428 66260 2440
rect 65843 2400 66260 2428
rect 65843 2397 65855 2400
rect 65797 2391 65855 2397
rect 66254 2388 66260 2400
rect 66312 2388 66318 2440
rect 66364 2437 66392 2468
rect 66349 2431 66407 2437
rect 66349 2397 66361 2431
rect 66395 2397 66407 2431
rect 66349 2391 66407 2397
rect 66438 2388 66444 2440
rect 66496 2428 66502 2440
rect 66901 2431 66959 2437
rect 66901 2428 66913 2431
rect 66496 2400 66913 2428
rect 66496 2388 66502 2400
rect 66901 2397 66913 2400
rect 66947 2397 66959 2431
rect 67450 2428 67456 2440
rect 67411 2400 67456 2428
rect 66901 2391 66959 2397
rect 67450 2388 67456 2400
rect 67508 2388 67514 2440
rect 68370 2428 68376 2440
rect 68331 2400 68376 2428
rect 68370 2388 68376 2400
rect 68428 2388 68434 2440
rect 68664 2428 68692 2536
rect 68848 2496 68876 2604
rect 69014 2592 69020 2604
rect 69072 2592 69078 2644
rect 70762 2632 70768 2644
rect 70723 2604 70768 2632
rect 70762 2592 70768 2604
rect 70820 2592 70826 2644
rect 71317 2635 71375 2641
rect 71317 2601 71329 2635
rect 71363 2632 71375 2635
rect 71406 2632 71412 2644
rect 71363 2604 71412 2632
rect 71363 2601 71375 2604
rect 71317 2595 71375 2601
rect 71406 2592 71412 2604
rect 71464 2592 71470 2644
rect 71590 2592 71596 2644
rect 71648 2632 71654 2644
rect 71648 2604 84194 2632
rect 71648 2592 71654 2604
rect 68922 2524 68928 2576
rect 68980 2564 68986 2576
rect 68980 2536 76052 2564
rect 68980 2524 68986 2536
rect 75089 2499 75147 2505
rect 75089 2496 75101 2499
rect 68848 2468 75101 2496
rect 75089 2465 75101 2468
rect 75135 2465 75147 2499
rect 75089 2459 75147 2465
rect 68830 2428 68836 2440
rect 68664 2400 68836 2428
rect 68830 2388 68836 2400
rect 68888 2388 68894 2440
rect 68922 2388 68928 2440
rect 68980 2428 68986 2440
rect 69201 2431 69259 2437
rect 69201 2428 69213 2431
rect 68980 2400 69213 2428
rect 68980 2388 68986 2400
rect 69201 2397 69213 2400
rect 69247 2397 69259 2431
rect 69201 2391 69259 2397
rect 69845 2431 69903 2437
rect 69845 2397 69857 2431
rect 69891 2397 69903 2431
rect 69845 2391 69903 2397
rect 69860 2360 69888 2391
rect 70210 2388 70216 2440
rect 70268 2428 70274 2440
rect 70949 2431 71007 2437
rect 70949 2428 70961 2431
rect 70268 2400 70961 2428
rect 70268 2388 70274 2400
rect 70949 2397 70961 2400
rect 70995 2397 71007 2431
rect 70949 2391 71007 2397
rect 71501 2431 71559 2437
rect 71501 2397 71513 2431
rect 71547 2397 71559 2431
rect 71501 2391 71559 2397
rect 64846 2332 69888 2360
rect 55456 2320 55462 2332
rect 70854 2320 70860 2372
rect 70912 2360 70918 2372
rect 71516 2360 71544 2391
rect 72142 2388 72148 2440
rect 72200 2428 72206 2440
rect 72237 2431 72295 2437
rect 72237 2428 72249 2431
rect 72200 2400 72249 2428
rect 72200 2388 72206 2400
rect 72237 2397 72249 2400
rect 72283 2397 72295 2431
rect 73522 2428 73528 2440
rect 73483 2400 73528 2428
rect 72237 2391 72295 2397
rect 73522 2388 73528 2400
rect 73580 2388 73586 2440
rect 74074 2388 74080 2440
rect 74132 2428 74138 2440
rect 74353 2431 74411 2437
rect 74353 2428 74365 2431
rect 74132 2400 74365 2428
rect 74132 2388 74138 2400
rect 74353 2397 74365 2400
rect 74399 2397 74411 2431
rect 74353 2391 74411 2397
rect 70912 2332 71544 2360
rect 70912 2320 70918 2332
rect 74718 2320 74724 2372
rect 74776 2360 74782 2372
rect 74905 2363 74963 2369
rect 74905 2360 74917 2363
rect 74776 2332 74917 2360
rect 74776 2320 74782 2332
rect 74905 2329 74917 2332
rect 74951 2329 74963 2363
rect 76024 2360 76052 2536
rect 78582 2524 78588 2576
rect 78640 2564 78646 2576
rect 79045 2567 79103 2573
rect 79045 2564 79057 2567
rect 78640 2536 79057 2564
rect 78640 2524 78646 2536
rect 79045 2533 79057 2536
rect 79091 2533 79103 2567
rect 79045 2527 79103 2533
rect 79226 2524 79232 2576
rect 79284 2564 79290 2576
rect 79965 2567 80023 2573
rect 79965 2564 79977 2567
rect 79284 2536 79977 2564
rect 79284 2524 79290 2536
rect 79965 2533 79977 2536
rect 80011 2533 80023 2567
rect 80790 2564 80796 2576
rect 80751 2536 80796 2564
rect 79965 2527 80023 2533
rect 80790 2524 80796 2536
rect 80848 2524 80854 2576
rect 81158 2524 81164 2576
rect 81216 2564 81222 2576
rect 81713 2567 81771 2573
rect 81713 2564 81725 2567
rect 81216 2536 81725 2564
rect 81216 2524 81222 2536
rect 81713 2533 81725 2536
rect 81759 2533 81771 2567
rect 84166 2564 84194 2604
rect 84166 2536 85436 2564
rect 81713 2527 81771 2533
rect 76116 2468 85344 2496
rect 76116 2437 76144 2468
rect 76101 2431 76159 2437
rect 76101 2397 76113 2431
rect 76147 2397 76159 2431
rect 76742 2428 76748 2440
rect 76703 2400 76748 2428
rect 76101 2391 76159 2397
rect 76742 2388 76748 2400
rect 76800 2388 76806 2440
rect 77018 2388 77024 2440
rect 77076 2428 77082 2440
rect 77573 2431 77631 2437
rect 77573 2428 77585 2431
rect 77076 2400 77585 2428
rect 77076 2388 77082 2400
rect 77573 2397 77585 2400
rect 77619 2397 77631 2431
rect 78677 2431 78735 2437
rect 78677 2428 78689 2431
rect 77573 2391 77631 2397
rect 77680 2400 78689 2428
rect 77680 2360 77708 2400
rect 78677 2397 78689 2400
rect 78723 2428 78735 2431
rect 79229 2431 79287 2437
rect 79229 2428 79241 2431
rect 78723 2400 79241 2428
rect 78723 2397 78735 2400
rect 78677 2391 78735 2397
rect 79229 2397 79241 2400
rect 79275 2397 79287 2431
rect 79502 2428 79508 2440
rect 79463 2400 79508 2428
rect 79229 2391 79287 2397
rect 79502 2388 79508 2400
rect 79560 2428 79566 2440
rect 79781 2431 79839 2437
rect 79781 2428 79793 2431
rect 79560 2400 79793 2428
rect 79560 2388 79566 2400
rect 79781 2397 79793 2400
rect 79827 2397 79839 2431
rect 79781 2391 79839 2397
rect 79962 2388 79968 2440
rect 80020 2428 80026 2440
rect 80149 2431 80207 2437
rect 80149 2428 80161 2431
rect 80020 2400 80161 2428
rect 80020 2388 80026 2400
rect 80149 2397 80161 2400
rect 80195 2397 80207 2431
rect 80149 2391 80207 2397
rect 80425 2431 80483 2437
rect 80425 2397 80437 2431
rect 80471 2397 80483 2431
rect 80425 2391 80483 2397
rect 76024 2332 77708 2360
rect 74905 2323 74963 2329
rect 77938 2320 77944 2372
rect 77996 2360 78002 2372
rect 77996 2332 79364 2360
rect 77996 2320 78002 2332
rect 50982 2292 50988 2304
rect 50672 2264 50717 2292
rect 50816 2264 50988 2292
rect 50672 2252 50678 2264
rect 50982 2252 50988 2264
rect 51040 2252 51046 2304
rect 51442 2292 51448 2304
rect 51403 2264 51448 2292
rect 51442 2252 51448 2264
rect 51500 2252 51506 2304
rect 53190 2292 53196 2304
rect 53151 2264 53196 2292
rect 53190 2252 53196 2264
rect 53248 2252 53254 2304
rect 54110 2252 54116 2304
rect 54168 2292 54174 2304
rect 54205 2295 54263 2301
rect 54205 2292 54217 2295
rect 54168 2264 54217 2292
rect 54168 2252 54174 2264
rect 54205 2261 54217 2264
rect 54251 2261 54263 2295
rect 54205 2255 54263 2261
rect 56042 2252 56048 2304
rect 56100 2292 56106 2304
rect 56413 2295 56471 2301
rect 56413 2292 56425 2295
rect 56100 2264 56425 2292
rect 56100 2252 56106 2264
rect 56413 2261 56425 2264
rect 56459 2261 56471 2295
rect 56413 2255 56471 2261
rect 56686 2252 56692 2304
rect 56744 2292 56750 2304
rect 56965 2295 57023 2301
rect 56965 2292 56977 2295
rect 56744 2264 56977 2292
rect 56744 2252 56750 2264
rect 56965 2261 56977 2264
rect 57011 2261 57023 2295
rect 56965 2255 57023 2261
rect 57330 2252 57336 2304
rect 57388 2292 57394 2304
rect 57885 2295 57943 2301
rect 57885 2292 57897 2295
rect 57388 2264 57897 2292
rect 57388 2252 57394 2264
rect 57885 2261 57897 2264
rect 57931 2261 57943 2295
rect 57885 2255 57943 2261
rect 57974 2252 57980 2304
rect 58032 2292 58038 2304
rect 58437 2295 58495 2301
rect 58437 2292 58449 2295
rect 58032 2264 58449 2292
rect 58032 2252 58038 2264
rect 58437 2261 58449 2264
rect 58483 2261 58495 2295
rect 58437 2255 58495 2261
rect 58618 2252 58624 2304
rect 58676 2292 58682 2304
rect 58989 2295 59047 2301
rect 58989 2292 59001 2295
rect 58676 2264 59001 2292
rect 58676 2252 58682 2264
rect 58989 2261 59001 2264
rect 59035 2261 59047 2295
rect 58989 2255 59047 2261
rect 61838 2252 61844 2304
rect 61896 2292 61902 2304
rect 61933 2295 61991 2301
rect 61933 2292 61945 2295
rect 61896 2264 61945 2292
rect 61896 2252 61902 2264
rect 61933 2261 61945 2264
rect 61979 2261 61991 2295
rect 61933 2255 61991 2261
rect 65058 2252 65064 2304
rect 65116 2292 65122 2304
rect 65613 2295 65671 2301
rect 65613 2292 65625 2295
rect 65116 2264 65625 2292
rect 65116 2252 65122 2264
rect 65613 2261 65625 2264
rect 65659 2261 65671 2295
rect 65613 2255 65671 2261
rect 65702 2252 65708 2304
rect 65760 2292 65766 2304
rect 66165 2295 66223 2301
rect 66165 2292 66177 2295
rect 65760 2264 66177 2292
rect 65760 2252 65766 2264
rect 66165 2261 66177 2264
rect 66211 2261 66223 2295
rect 66714 2292 66720 2304
rect 66675 2264 66720 2292
rect 66165 2255 66223 2261
rect 66714 2252 66720 2264
rect 66772 2252 66778 2304
rect 67174 2252 67180 2304
rect 67232 2292 67238 2304
rect 67269 2295 67327 2301
rect 67269 2292 67281 2295
rect 67232 2264 67281 2292
rect 67232 2252 67238 2264
rect 67269 2261 67281 2264
rect 67315 2261 67327 2295
rect 67269 2255 67327 2261
rect 67634 2252 67640 2304
rect 67692 2292 67698 2304
rect 68189 2295 68247 2301
rect 68189 2292 68201 2295
rect 67692 2264 68201 2292
rect 67692 2252 67698 2264
rect 68189 2261 68201 2264
rect 68235 2261 68247 2295
rect 68189 2255 68247 2261
rect 69566 2252 69572 2304
rect 69624 2292 69630 2304
rect 69661 2295 69719 2301
rect 69661 2292 69673 2295
rect 69624 2264 69673 2292
rect 69624 2252 69630 2264
rect 69661 2261 69673 2264
rect 69707 2261 69719 2295
rect 72418 2292 72424 2304
rect 72379 2264 72424 2292
rect 69661 2255 69719 2261
rect 72418 2252 72424 2264
rect 72476 2252 72482 2304
rect 72786 2252 72792 2304
rect 72844 2292 72850 2304
rect 73341 2295 73399 2301
rect 73341 2292 73353 2295
rect 72844 2264 73353 2292
rect 72844 2252 72850 2264
rect 73341 2261 73353 2264
rect 73387 2261 73399 2295
rect 73341 2255 73399 2261
rect 75362 2252 75368 2304
rect 75420 2292 75426 2304
rect 75917 2295 75975 2301
rect 75917 2292 75929 2295
rect 75420 2264 75929 2292
rect 75420 2252 75426 2264
rect 75917 2261 75929 2264
rect 75963 2261 75975 2295
rect 75917 2255 75975 2261
rect 76561 2295 76619 2301
rect 76561 2261 76573 2295
rect 76607 2292 76619 2295
rect 76650 2292 76656 2304
rect 76607 2264 76656 2292
rect 76607 2261 76619 2264
rect 76561 2255 76619 2261
rect 76650 2252 76656 2264
rect 76708 2252 76714 2304
rect 77018 2292 77024 2304
rect 76979 2264 77024 2292
rect 77018 2252 77024 2264
rect 77076 2252 77082 2304
rect 77294 2252 77300 2304
rect 77352 2292 77358 2304
rect 79336 2301 79364 2332
rect 79686 2320 79692 2372
rect 79744 2360 79750 2372
rect 80440 2360 80468 2391
rect 80514 2388 80520 2440
rect 80572 2428 80578 2440
rect 80609 2431 80667 2437
rect 80609 2428 80621 2431
rect 80572 2400 80621 2428
rect 80572 2388 80578 2400
rect 80609 2397 80621 2400
rect 80655 2397 80667 2431
rect 81897 2431 81955 2437
rect 81897 2428 81909 2431
rect 80609 2391 80667 2397
rect 81452 2400 81909 2428
rect 79744 2332 80468 2360
rect 79744 2320 79750 2332
rect 81452 2304 81480 2400
rect 81897 2397 81909 2400
rect 81943 2397 81955 2431
rect 83826 2428 83832 2440
rect 83787 2400 83832 2428
rect 81897 2391 81955 2397
rect 83826 2388 83832 2400
rect 83884 2388 83890 2440
rect 84657 2431 84715 2437
rect 84657 2428 84669 2431
rect 84212 2400 84669 2428
rect 82446 2320 82452 2372
rect 82504 2360 82510 2372
rect 82633 2363 82691 2369
rect 82633 2360 82645 2363
rect 82504 2332 82645 2360
rect 82504 2320 82510 2332
rect 82633 2329 82645 2332
rect 82679 2329 82691 2363
rect 82633 2323 82691 2329
rect 84212 2304 84240 2400
rect 84657 2397 84669 2400
rect 84703 2397 84715 2431
rect 84657 2391 84715 2397
rect 85022 2388 85028 2440
rect 85080 2428 85086 2440
rect 85117 2431 85175 2437
rect 85117 2428 85129 2431
rect 85080 2400 85129 2428
rect 85080 2388 85086 2400
rect 85117 2397 85129 2400
rect 85163 2397 85175 2431
rect 85117 2391 85175 2397
rect 85316 2360 85344 2468
rect 85408 2428 85436 2536
rect 86310 2524 86316 2576
rect 86368 2564 86374 2576
rect 86865 2567 86923 2573
rect 86865 2564 86877 2567
rect 86368 2536 86877 2564
rect 86368 2524 86374 2536
rect 86865 2533 86877 2536
rect 86911 2533 86923 2567
rect 86865 2527 86923 2533
rect 85482 2456 85488 2508
rect 85540 2496 85546 2508
rect 85540 2468 87092 2496
rect 85540 2456 85546 2468
rect 87064 2437 87092 2468
rect 86405 2431 86463 2437
rect 86405 2428 86417 2431
rect 85408 2400 86417 2428
rect 86405 2397 86417 2400
rect 86451 2428 86463 2431
rect 86681 2431 86739 2437
rect 86681 2428 86693 2431
rect 86451 2400 86693 2428
rect 86451 2397 86463 2400
rect 86405 2391 86463 2397
rect 86681 2397 86693 2400
rect 86727 2397 86739 2431
rect 86681 2391 86739 2397
rect 87049 2431 87107 2437
rect 87049 2397 87061 2431
rect 87095 2397 87107 2431
rect 87049 2391 87107 2397
rect 87877 2363 87935 2369
rect 85316 2332 87092 2360
rect 87064 2304 87092 2332
rect 87877 2329 87889 2363
rect 87923 2360 87935 2363
rect 88886 2360 88892 2372
rect 87923 2332 88892 2360
rect 87923 2329 87935 2332
rect 87877 2323 87935 2329
rect 88886 2320 88892 2332
rect 88944 2320 88950 2372
rect 77389 2295 77447 2301
rect 77389 2292 77401 2295
rect 77352 2264 77401 2292
rect 77352 2252 77358 2264
rect 77389 2261 77401 2264
rect 77435 2261 77447 2295
rect 77389 2255 77447 2261
rect 79321 2295 79379 2301
rect 79321 2261 79333 2295
rect 79367 2261 79379 2295
rect 79321 2255 79379 2261
rect 80054 2252 80060 2304
rect 80112 2292 80118 2304
rect 80241 2295 80299 2301
rect 80241 2292 80253 2295
rect 80112 2264 80253 2292
rect 80112 2252 80118 2264
rect 80241 2261 80253 2264
rect 80287 2261 80299 2295
rect 81434 2292 81440 2304
rect 81395 2264 81440 2292
rect 80241 2255 80299 2261
rect 81434 2252 81440 2264
rect 81492 2252 81498 2304
rect 82722 2292 82728 2304
rect 82683 2264 82728 2292
rect 82722 2252 82728 2264
rect 82780 2252 82786 2304
rect 83090 2252 83096 2304
rect 83148 2292 83154 2304
rect 83645 2295 83703 2301
rect 83645 2292 83657 2295
rect 83148 2264 83657 2292
rect 83148 2252 83154 2264
rect 83645 2261 83657 2264
rect 83691 2261 83703 2295
rect 83645 2255 83703 2261
rect 84194 2252 84200 2304
rect 84252 2292 84258 2304
rect 84252 2264 84297 2292
rect 84252 2252 84258 2264
rect 84378 2252 84384 2304
rect 84436 2292 84442 2304
rect 84473 2295 84531 2301
rect 84473 2292 84485 2295
rect 84436 2264 84485 2292
rect 84436 2252 84442 2264
rect 84473 2261 84485 2264
rect 84519 2261 84531 2295
rect 85298 2292 85304 2304
rect 85259 2264 85304 2292
rect 84473 2255 84531 2261
rect 85298 2252 85304 2264
rect 85356 2252 85362 2304
rect 85666 2252 85672 2304
rect 85724 2292 85730 2304
rect 86221 2295 86279 2301
rect 86221 2292 86233 2295
rect 85724 2264 86233 2292
rect 85724 2252 85730 2264
rect 86221 2261 86233 2264
rect 86267 2261 86279 2295
rect 86221 2255 86279 2261
rect 87046 2252 87052 2304
rect 87104 2252 87110 2304
rect 87966 2292 87972 2304
rect 87927 2264 87972 2292
rect 87966 2252 87972 2264
rect 88024 2252 88030 2304
rect 1104 2202 88872 2224
rect 1104 2150 22898 2202
rect 22950 2150 22962 2202
rect 23014 2150 23026 2202
rect 23078 2150 23090 2202
rect 23142 2150 23154 2202
rect 23206 2150 44846 2202
rect 44898 2150 44910 2202
rect 44962 2150 44974 2202
rect 45026 2150 45038 2202
rect 45090 2150 45102 2202
rect 45154 2150 66794 2202
rect 66846 2150 66858 2202
rect 66910 2150 66922 2202
rect 66974 2150 66986 2202
rect 67038 2150 67050 2202
rect 67102 2150 88872 2202
rect 1104 2128 88872 2150
rect 24762 2048 24768 2100
rect 24820 2088 24826 2100
rect 28810 2088 28816 2100
rect 24820 2060 28816 2088
rect 24820 2048 24826 2060
rect 28810 2048 28816 2060
rect 28868 2048 28874 2100
rect 28902 2048 28908 2100
rect 28960 2088 28966 2100
rect 62022 2088 62028 2100
rect 28960 2060 62028 2088
rect 28960 2048 28966 2060
rect 62022 2048 62028 2060
rect 62080 2048 62086 2100
rect 64690 2048 64696 2100
rect 64748 2088 64754 2100
rect 82722 2088 82728 2100
rect 64748 2060 82728 2088
rect 64748 2048 64754 2060
rect 82722 2048 82728 2060
rect 82780 2048 82786 2100
rect 15746 1980 15752 2032
rect 15804 2020 15810 2032
rect 45554 2020 45560 2032
rect 15804 1992 45560 2020
rect 15804 1980 15810 1992
rect 45554 1980 45560 1992
rect 45612 1980 45618 2032
rect 45646 1980 45652 2032
rect 45704 2020 45710 2032
rect 48774 2020 48780 2032
rect 45704 1992 48780 2020
rect 45704 1980 45710 1992
rect 48774 1980 48780 1992
rect 48832 1980 48838 2032
rect 48866 1980 48872 2032
rect 48924 2020 48930 2032
rect 50430 2020 50436 2032
rect 48924 1992 50436 2020
rect 48924 1980 48930 1992
rect 50430 1980 50436 1992
rect 50488 1980 50494 2032
rect 50614 1980 50620 2032
rect 50672 2020 50678 2032
rect 51626 2020 51632 2032
rect 50672 1992 51632 2020
rect 50672 1980 50678 1992
rect 51626 1980 51632 1992
rect 51684 1980 51690 2032
rect 52914 1980 52920 2032
rect 52972 2020 52978 2032
rect 81434 2020 81440 2032
rect 52972 1992 81440 2020
rect 52972 1980 52978 1992
rect 81434 1980 81440 1992
rect 81492 1980 81498 2032
rect 8202 1912 8208 1964
rect 8260 1952 8266 1964
rect 8260 1924 12572 1952
rect 8260 1912 8266 1924
rect 12544 1884 12572 1924
rect 22186 1912 22192 1964
rect 22244 1952 22250 1964
rect 28902 1952 28908 1964
rect 22244 1924 28908 1952
rect 22244 1912 22250 1924
rect 28902 1912 28908 1924
rect 28960 1912 28966 1964
rect 59354 1952 59360 1964
rect 29104 1924 59360 1952
rect 27798 1884 27804 1896
rect 6886 1856 12434 1884
rect 12544 1856 27804 1884
rect 2866 1776 2872 1828
rect 2924 1816 2930 1828
rect 6886 1816 6914 1856
rect 2924 1788 6914 1816
rect 12406 1816 12434 1856
rect 27798 1844 27804 1856
rect 27856 1844 27862 1896
rect 12406 1788 24348 1816
rect 2924 1776 2930 1788
rect 10502 1708 10508 1760
rect 10560 1748 10566 1760
rect 24210 1748 24216 1760
rect 10560 1720 24216 1748
rect 10560 1708 10566 1720
rect 24210 1708 24216 1720
rect 24268 1708 24274 1760
rect 24320 1748 24348 1788
rect 24394 1776 24400 1828
rect 24452 1816 24458 1828
rect 26326 1816 26332 1828
rect 24452 1788 26332 1816
rect 24452 1776 24458 1788
rect 26326 1776 26332 1788
rect 26384 1776 26390 1828
rect 26510 1776 26516 1828
rect 26568 1816 26574 1828
rect 26568 1788 26740 1816
rect 26568 1776 26574 1788
rect 26602 1748 26608 1760
rect 24320 1720 26608 1748
rect 26602 1708 26608 1720
rect 26660 1708 26666 1760
rect 26712 1748 26740 1788
rect 26970 1776 26976 1828
rect 27028 1816 27034 1828
rect 27706 1816 27712 1828
rect 27028 1788 27712 1816
rect 27028 1776 27034 1788
rect 27706 1776 27712 1788
rect 27764 1776 27770 1828
rect 29104 1816 29132 1924
rect 59354 1912 59360 1924
rect 59412 1912 59418 1964
rect 63402 1912 63408 1964
rect 63460 1952 63466 1964
rect 66714 1952 66720 1964
rect 63460 1924 66720 1952
rect 63460 1912 63466 1924
rect 66714 1912 66720 1924
rect 66772 1912 66778 1964
rect 31662 1844 31668 1896
rect 31720 1884 31726 1896
rect 53190 1884 53196 1896
rect 31720 1856 53196 1884
rect 31720 1844 31726 1856
rect 53190 1844 53196 1856
rect 53248 1844 53254 1896
rect 58986 1844 58992 1896
rect 59044 1884 59050 1896
rect 62298 1884 62304 1896
rect 59044 1856 62304 1884
rect 59044 1844 59050 1856
rect 62298 1844 62304 1856
rect 62356 1844 62362 1896
rect 64138 1844 64144 1896
rect 64196 1884 64202 1896
rect 76742 1884 76748 1896
rect 64196 1856 76748 1884
rect 64196 1844 64202 1856
rect 76742 1844 76748 1856
rect 76800 1844 76806 1896
rect 28000 1788 29132 1816
rect 28000 1748 28028 1788
rect 31386 1776 31392 1828
rect 31444 1816 31450 1828
rect 84194 1816 84200 1828
rect 31444 1788 84200 1816
rect 31444 1776 31450 1788
rect 84194 1776 84200 1788
rect 84252 1776 84258 1828
rect 26712 1720 28028 1748
rect 28626 1708 28632 1760
rect 28684 1748 28690 1760
rect 87966 1748 87972 1760
rect 28684 1720 87972 1748
rect 28684 1708 28690 1720
rect 87966 1708 87972 1720
rect 88024 1708 88030 1760
rect 12342 1640 12348 1692
rect 12400 1680 12406 1692
rect 45554 1680 45560 1692
rect 12400 1652 45560 1680
rect 12400 1640 12406 1652
rect 45554 1640 45560 1652
rect 45612 1640 45618 1692
rect 45830 1640 45836 1692
rect 45888 1680 45894 1692
rect 79502 1680 79508 1692
rect 45888 1652 79508 1680
rect 45888 1640 45894 1652
rect 79502 1640 79508 1652
rect 79560 1640 79566 1692
rect 16942 1572 16948 1624
rect 17000 1612 17006 1624
rect 45370 1612 45376 1624
rect 17000 1584 45376 1612
rect 17000 1572 17006 1584
rect 45370 1572 45376 1584
rect 45428 1572 45434 1624
rect 47118 1572 47124 1624
rect 47176 1612 47182 1624
rect 85298 1612 85304 1624
rect 47176 1584 85304 1612
rect 47176 1572 47182 1584
rect 85298 1572 85304 1584
rect 85356 1572 85362 1624
rect 4246 1504 4252 1556
rect 4304 1544 4310 1556
rect 26050 1544 26056 1556
rect 4304 1516 26056 1544
rect 4304 1504 4310 1516
rect 26050 1504 26056 1516
rect 26108 1504 26114 1556
rect 26142 1504 26148 1556
rect 26200 1544 26206 1556
rect 30190 1544 30196 1556
rect 26200 1516 30196 1544
rect 26200 1504 26206 1516
rect 30190 1504 30196 1516
rect 30248 1504 30254 1556
rect 30282 1504 30288 1556
rect 30340 1544 30346 1556
rect 31754 1544 31760 1556
rect 30340 1516 31760 1544
rect 30340 1504 30346 1516
rect 31754 1504 31760 1516
rect 31812 1504 31818 1556
rect 31846 1504 31852 1556
rect 31904 1544 31910 1556
rect 72418 1544 72424 1556
rect 31904 1516 72424 1544
rect 31904 1504 31910 1516
rect 72418 1504 72424 1516
rect 72476 1504 72482 1556
rect 22002 1436 22008 1488
rect 22060 1476 22066 1488
rect 51442 1476 51448 1488
rect 22060 1448 51448 1476
rect 22060 1436 22066 1448
rect 51442 1436 51448 1448
rect 51500 1436 51506 1488
rect 62206 1476 62212 1488
rect 51552 1448 62212 1476
rect 14366 1368 14372 1420
rect 14424 1408 14430 1420
rect 23566 1408 23572 1420
rect 14424 1380 23572 1408
rect 14424 1368 14430 1380
rect 23566 1368 23572 1380
rect 23624 1368 23630 1420
rect 23934 1368 23940 1420
rect 23992 1408 23998 1420
rect 30282 1408 30288 1420
rect 23992 1380 30288 1408
rect 23992 1368 23998 1380
rect 30282 1368 30288 1380
rect 30340 1368 30346 1420
rect 45554 1408 45560 1420
rect 30392 1380 45560 1408
rect 26050 1300 26056 1352
rect 26108 1340 26114 1352
rect 29086 1340 29092 1352
rect 26108 1312 29092 1340
rect 26108 1300 26114 1312
rect 29086 1300 29092 1312
rect 29144 1300 29150 1352
rect 25866 1232 25872 1284
rect 25924 1272 25930 1284
rect 30392 1272 30420 1380
rect 45554 1368 45560 1380
rect 45612 1368 45618 1420
rect 45738 1368 45744 1420
rect 45796 1368 45802 1420
rect 47118 1408 47124 1420
rect 45848 1380 47124 1408
rect 45370 1300 45376 1352
rect 45428 1340 45434 1352
rect 45756 1340 45784 1368
rect 45428 1312 45784 1340
rect 45428 1300 45434 1312
rect 25924 1244 30420 1272
rect 25924 1232 25930 1244
rect 38654 1232 38660 1284
rect 38712 1272 38718 1284
rect 39114 1272 39120 1284
rect 38712 1244 39120 1272
rect 38712 1232 38718 1244
rect 39114 1232 39120 1244
rect 39172 1232 39178 1284
rect 39206 1232 39212 1284
rect 39264 1272 39270 1284
rect 45848 1272 45876 1380
rect 47118 1368 47124 1380
rect 47176 1368 47182 1420
rect 50798 1408 50804 1420
rect 47228 1380 50804 1408
rect 46750 1300 46756 1352
rect 46808 1340 46814 1352
rect 47228 1340 47256 1380
rect 50798 1368 50804 1380
rect 50856 1368 50862 1420
rect 51552 1408 51580 1448
rect 62206 1436 62212 1448
rect 62264 1436 62270 1488
rect 62298 1436 62304 1488
rect 62356 1476 62362 1488
rect 71590 1476 71596 1488
rect 62356 1448 71596 1476
rect 62356 1436 62362 1448
rect 71590 1436 71596 1448
rect 71648 1436 71654 1488
rect 77018 1476 77024 1488
rect 74506 1448 77024 1476
rect 50908 1380 51580 1408
rect 46808 1312 47256 1340
rect 46808 1300 46814 1312
rect 49418 1300 49424 1352
rect 49476 1340 49482 1352
rect 50908 1340 50936 1380
rect 51626 1368 51632 1420
rect 51684 1408 51690 1420
rect 63494 1408 63500 1420
rect 51684 1380 63500 1408
rect 51684 1368 51690 1380
rect 63494 1368 63500 1380
rect 63552 1368 63558 1420
rect 64046 1368 64052 1420
rect 64104 1408 64110 1420
rect 74506 1408 74534 1448
rect 77018 1436 77024 1448
rect 77076 1436 77082 1488
rect 64104 1380 74534 1408
rect 64104 1368 64110 1380
rect 49476 1312 50936 1340
rect 49476 1300 49482 1312
rect 39264 1244 45876 1272
rect 39264 1232 39270 1244
rect 27614 1164 27620 1216
rect 27672 1204 27678 1216
rect 28350 1204 28356 1216
rect 27672 1176 28356 1204
rect 27672 1164 27678 1176
rect 28350 1164 28356 1176
rect 28408 1164 28414 1216
<< via1 >>
rect 11924 27718 11976 27770
rect 11988 27718 12040 27770
rect 12052 27718 12104 27770
rect 12116 27718 12168 27770
rect 12180 27718 12232 27770
rect 33872 27718 33924 27770
rect 33936 27718 33988 27770
rect 34000 27718 34052 27770
rect 34064 27718 34116 27770
rect 34128 27718 34180 27770
rect 55820 27718 55872 27770
rect 55884 27718 55936 27770
rect 55948 27718 56000 27770
rect 56012 27718 56064 27770
rect 56076 27718 56128 27770
rect 77768 27718 77820 27770
rect 77832 27718 77884 27770
rect 77896 27718 77948 27770
rect 77960 27718 78012 27770
rect 78024 27718 78076 27770
rect 25872 27616 25924 27668
rect 2688 27591 2740 27600
rect 2688 27557 2697 27591
rect 2697 27557 2731 27591
rect 2731 27557 2740 27591
rect 2688 27548 2740 27557
rect 5264 27591 5316 27600
rect 5264 27557 5273 27591
rect 5273 27557 5307 27591
rect 5307 27557 5316 27591
rect 5264 27548 5316 27557
rect 7748 27591 7800 27600
rect 7748 27557 7757 27591
rect 7757 27557 7791 27591
rect 7791 27557 7800 27591
rect 7748 27548 7800 27557
rect 8484 27591 8536 27600
rect 8484 27557 8493 27591
rect 8493 27557 8527 27591
rect 8527 27557 8536 27591
rect 8484 27548 8536 27557
rect 9128 27591 9180 27600
rect 9128 27557 9137 27591
rect 9137 27557 9171 27591
rect 9171 27557 9180 27591
rect 9128 27548 9180 27557
rect 9220 27548 9272 27600
rect 12164 27548 12216 27600
rect 14280 27591 14332 27600
rect 14280 27557 14289 27591
rect 14289 27557 14323 27591
rect 14323 27557 14332 27591
rect 14280 27548 14332 27557
rect 14924 27591 14976 27600
rect 14924 27557 14933 27591
rect 14933 27557 14967 27591
rect 14967 27557 14976 27591
rect 14924 27548 14976 27557
rect 15568 27591 15620 27600
rect 15568 27557 15577 27591
rect 15577 27557 15611 27591
rect 15611 27557 15620 27591
rect 15568 27548 15620 27557
rect 18052 27591 18104 27600
rect 18052 27557 18061 27591
rect 18061 27557 18095 27591
rect 18095 27557 18104 27591
rect 18052 27548 18104 27557
rect 18604 27591 18656 27600
rect 18604 27557 18613 27591
rect 18613 27557 18647 27591
rect 18647 27557 18656 27591
rect 18604 27548 18656 27557
rect 19984 27548 20036 27600
rect 20628 27591 20680 27600
rect 20628 27557 20637 27591
rect 20637 27557 20671 27591
rect 20671 27557 20680 27591
rect 20628 27548 20680 27557
rect 22008 27591 22060 27600
rect 22008 27557 22017 27591
rect 22017 27557 22051 27591
rect 22051 27557 22060 27591
rect 22008 27548 22060 27557
rect 22560 27591 22612 27600
rect 22560 27557 22569 27591
rect 22569 27557 22603 27591
rect 22603 27557 22612 27591
rect 22560 27548 22612 27557
rect 24584 27591 24636 27600
rect 5816 27480 5868 27532
rect 11612 27523 11664 27532
rect 1308 27412 1360 27464
rect 2228 27455 2280 27464
rect 2228 27421 2237 27455
rect 2237 27421 2271 27455
rect 2271 27421 2280 27455
rect 2228 27412 2280 27421
rect 3148 27412 3200 27464
rect 3240 27412 3292 27464
rect 4712 27455 4764 27464
rect 4712 27421 4721 27455
rect 4721 27421 4755 27455
rect 4755 27421 4764 27455
rect 4712 27412 4764 27421
rect 6644 27455 6696 27464
rect 6644 27421 6653 27455
rect 6653 27421 6687 27455
rect 6687 27421 6696 27455
rect 6644 27412 6696 27421
rect 9220 27412 9272 27464
rect 9680 27412 9732 27464
rect 10508 27455 10560 27464
rect 10508 27421 10517 27455
rect 10517 27421 10551 27455
rect 10551 27421 10560 27455
rect 10508 27412 10560 27421
rect 11612 27489 11621 27523
rect 11621 27489 11655 27523
rect 11655 27489 11664 27523
rect 11612 27480 11664 27489
rect 23112 27523 23164 27532
rect 23112 27489 23121 27523
rect 23121 27489 23155 27523
rect 23155 27489 23164 27523
rect 23112 27480 23164 27489
rect 24584 27557 24593 27591
rect 24593 27557 24627 27591
rect 24627 27557 24636 27591
rect 24584 27548 24636 27557
rect 26424 27548 26476 27600
rect 27160 27591 27212 27600
rect 27160 27557 27169 27591
rect 27169 27557 27203 27591
rect 27203 27557 27212 27591
rect 27160 27548 27212 27557
rect 27804 27591 27856 27600
rect 27804 27557 27813 27591
rect 27813 27557 27847 27591
rect 27847 27557 27856 27591
rect 27804 27548 27856 27557
rect 31300 27616 31352 27668
rect 36544 27616 36596 27668
rect 29736 27591 29788 27600
rect 29736 27557 29745 27591
rect 29745 27557 29779 27591
rect 29779 27557 29788 27591
rect 29736 27548 29788 27557
rect 33508 27591 33560 27600
rect 33508 27557 33517 27591
rect 33517 27557 33551 27591
rect 33551 27557 33560 27591
rect 33508 27548 33560 27557
rect 34244 27548 34296 27600
rect 34888 27591 34940 27600
rect 34888 27557 34897 27591
rect 34897 27557 34931 27591
rect 34931 27557 34940 27591
rect 34888 27548 34940 27557
rect 35532 27591 35584 27600
rect 35532 27557 35541 27591
rect 35541 27557 35575 27591
rect 35575 27557 35584 27591
rect 35532 27548 35584 27557
rect 36084 27591 36136 27600
rect 36084 27557 36093 27591
rect 36093 27557 36127 27591
rect 36127 27557 36136 27591
rect 36084 27548 36136 27557
rect 36176 27548 36228 27600
rect 37280 27548 37332 27600
rect 37464 27591 37516 27600
rect 37464 27557 37473 27591
rect 37473 27557 37507 27591
rect 37507 27557 37516 27591
rect 37464 27548 37516 27557
rect 37556 27548 37608 27600
rect 38108 27591 38160 27600
rect 38108 27557 38117 27591
rect 38117 27557 38151 27591
rect 38151 27557 38160 27591
rect 38108 27548 38160 27557
rect 38752 27591 38804 27600
rect 38752 27557 38761 27591
rect 38761 27557 38795 27591
rect 38795 27557 38804 27591
rect 38752 27548 38804 27557
rect 39304 27548 39356 27600
rect 40684 27591 40736 27600
rect 40684 27557 40693 27591
rect 40693 27557 40727 27591
rect 40727 27557 40736 27591
rect 40684 27548 40736 27557
rect 42616 27591 42668 27600
rect 29368 27480 29420 27532
rect 30840 27523 30892 27532
rect 30840 27489 30849 27523
rect 30849 27489 30883 27523
rect 30883 27489 30892 27523
rect 30840 27480 30892 27489
rect 31576 27480 31628 27532
rect 32680 27480 32732 27532
rect 42616 27557 42625 27591
rect 42625 27557 42659 27591
rect 42659 27557 42668 27591
rect 42616 27548 42668 27557
rect 43260 27591 43312 27600
rect 43260 27557 43269 27591
rect 43269 27557 43303 27591
rect 43303 27557 43312 27591
rect 43260 27548 43312 27557
rect 43812 27591 43864 27600
rect 43812 27557 43821 27591
rect 43821 27557 43855 27591
rect 43855 27557 43864 27591
rect 43812 27548 43864 27557
rect 45192 27591 45244 27600
rect 45192 27557 45201 27591
rect 45201 27557 45235 27591
rect 45235 27557 45244 27591
rect 45192 27548 45244 27557
rect 45836 27591 45888 27600
rect 45836 27557 45845 27591
rect 45845 27557 45879 27591
rect 45879 27557 45888 27591
rect 45836 27548 45888 27557
rect 46480 27591 46532 27600
rect 46480 27557 46489 27591
rect 46489 27557 46523 27591
rect 46523 27557 46532 27591
rect 46480 27548 46532 27557
rect 52276 27616 52328 27668
rect 49056 27591 49108 27600
rect 49056 27557 49065 27591
rect 49065 27557 49099 27591
rect 49099 27557 49108 27591
rect 49056 27548 49108 27557
rect 51080 27591 51132 27600
rect 51080 27557 51089 27591
rect 51089 27557 51123 27591
rect 51123 27557 51132 27591
rect 51080 27548 51132 27557
rect 51264 27548 51316 27600
rect 52460 27548 52512 27600
rect 55680 27548 55732 27600
rect 56232 27548 56284 27600
rect 56784 27591 56836 27600
rect 56784 27557 56793 27591
rect 56793 27557 56827 27591
rect 56827 27557 56836 27591
rect 56784 27548 56836 27557
rect 57336 27548 57388 27600
rect 59360 27591 59412 27600
rect 59360 27557 59369 27591
rect 59369 27557 59403 27591
rect 59403 27557 59412 27591
rect 59360 27548 59412 27557
rect 59912 27548 59964 27600
rect 60556 27548 60608 27600
rect 61936 27591 61988 27600
rect 61936 27557 61945 27591
rect 61945 27557 61979 27591
rect 61979 27557 61988 27591
rect 61936 27548 61988 27557
rect 62488 27548 62540 27600
rect 65064 27548 65116 27600
rect 65708 27548 65760 27600
rect 66352 27548 66404 27600
rect 69020 27548 69072 27600
rect 70400 27548 70452 27600
rect 71504 27548 71556 27600
rect 72424 27591 72476 27600
rect 72424 27557 72433 27591
rect 72433 27557 72467 27591
rect 72467 27557 72476 27591
rect 72424 27548 72476 27557
rect 74264 27591 74316 27600
rect 74264 27557 74273 27591
rect 74273 27557 74307 27591
rect 74307 27557 74316 27591
rect 74264 27548 74316 27557
rect 74816 27591 74868 27600
rect 74816 27557 74825 27591
rect 74825 27557 74859 27591
rect 74859 27557 74868 27591
rect 74816 27548 74868 27557
rect 76840 27591 76892 27600
rect 76840 27557 76849 27591
rect 76849 27557 76883 27591
rect 76883 27557 76892 27591
rect 76840 27548 76892 27557
rect 77392 27591 77444 27600
rect 77392 27557 77401 27591
rect 77401 27557 77435 27591
rect 77435 27557 77444 27591
rect 77392 27548 77444 27557
rect 81992 27591 82044 27600
rect 81992 27557 82001 27591
rect 82001 27557 82035 27591
rect 82035 27557 82044 27591
rect 81992 27548 82044 27557
rect 83096 27548 83148 27600
rect 83740 27548 83792 27600
rect 85672 27548 85724 27600
rect 12256 27412 12308 27464
rect 12808 27455 12860 27464
rect 12808 27421 12817 27455
rect 12817 27421 12851 27455
rect 12851 27421 12860 27455
rect 12808 27412 12860 27421
rect 13084 27455 13136 27464
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 14464 27455 14516 27464
rect 14464 27421 14473 27455
rect 14473 27421 14507 27455
rect 14507 27421 14516 27455
rect 14464 27412 14516 27421
rect 15108 27455 15160 27464
rect 15108 27421 15117 27455
rect 15117 27421 15151 27455
rect 15151 27421 15160 27455
rect 15108 27412 15160 27421
rect 15752 27455 15804 27464
rect 15752 27421 15761 27455
rect 15761 27421 15795 27455
rect 15795 27421 15804 27455
rect 15752 27412 15804 27421
rect 16580 27412 16632 27464
rect 18052 27412 18104 27464
rect 18236 27455 18288 27464
rect 18236 27421 18245 27455
rect 18245 27421 18279 27455
rect 18279 27421 18288 27455
rect 18236 27412 18288 27421
rect 18788 27455 18840 27464
rect 18788 27421 18797 27455
rect 18797 27421 18831 27455
rect 18831 27421 18840 27455
rect 18788 27412 18840 27421
rect 19616 27455 19668 27464
rect 19616 27421 19625 27455
rect 19625 27421 19659 27455
rect 19659 27421 19668 27455
rect 19616 27412 19668 27421
rect 20260 27455 20312 27464
rect 20260 27421 20269 27455
rect 20269 27421 20303 27455
rect 20303 27421 20312 27455
rect 20260 27412 20312 27421
rect 20352 27412 20404 27464
rect 21364 27455 21416 27464
rect 21364 27421 21373 27455
rect 21373 27421 21407 27455
rect 21407 27421 21416 27455
rect 21364 27412 21416 27421
rect 22192 27455 22244 27464
rect 22192 27421 22201 27455
rect 22201 27421 22235 27455
rect 22235 27421 22244 27455
rect 22192 27412 22244 27421
rect 1676 27276 1728 27328
rect 4068 27276 4120 27328
rect 4804 27319 4856 27328
rect 4804 27285 4813 27319
rect 4813 27285 4847 27319
rect 4847 27285 4856 27319
rect 4804 27276 4856 27285
rect 9680 27319 9732 27328
rect 9680 27285 9689 27319
rect 9689 27285 9723 27319
rect 9723 27285 9732 27319
rect 9680 27276 9732 27285
rect 10968 27344 11020 27396
rect 12164 27344 12216 27396
rect 17132 27344 17184 27396
rect 20444 27344 20496 27396
rect 22836 27412 22888 27464
rect 23388 27455 23440 27464
rect 23388 27421 23397 27455
rect 23397 27421 23431 27455
rect 23431 27421 23440 27455
rect 23388 27412 23440 27421
rect 24584 27412 24636 27464
rect 25964 27455 26016 27464
rect 19800 27276 19852 27328
rect 25412 27344 25464 27396
rect 25964 27421 25973 27455
rect 25973 27421 26007 27455
rect 26007 27421 26016 27455
rect 25964 27412 26016 27421
rect 26700 27412 26752 27464
rect 28172 27412 28224 27464
rect 28356 27412 28408 27464
rect 29092 27455 29144 27464
rect 29092 27421 29101 27455
rect 29101 27421 29135 27455
rect 29135 27421 29144 27455
rect 29092 27412 29144 27421
rect 29920 27455 29972 27464
rect 29920 27421 29929 27455
rect 29929 27421 29963 27455
rect 29963 27421 29972 27455
rect 29920 27412 29972 27421
rect 31116 27455 31168 27464
rect 31116 27421 31125 27455
rect 31125 27421 31159 27455
rect 31159 27421 31168 27455
rect 31116 27412 31168 27421
rect 31852 27412 31904 27464
rect 33692 27455 33744 27464
rect 33692 27421 33701 27455
rect 33701 27421 33735 27455
rect 33735 27421 33744 27455
rect 33692 27412 33744 27421
rect 34244 27455 34296 27464
rect 34244 27421 34253 27455
rect 34253 27421 34287 27455
rect 34287 27421 34296 27455
rect 34244 27412 34296 27421
rect 35072 27455 35124 27464
rect 35072 27421 35081 27455
rect 35081 27421 35115 27455
rect 35115 27421 35124 27455
rect 35072 27412 35124 27421
rect 35716 27455 35768 27464
rect 35716 27421 35725 27455
rect 35725 27421 35759 27455
rect 35759 27421 35768 27455
rect 35716 27412 35768 27421
rect 36820 27455 36872 27464
rect 27252 27344 27304 27396
rect 21272 27276 21324 27328
rect 25872 27276 25924 27328
rect 26056 27319 26108 27328
rect 26056 27285 26065 27319
rect 26065 27285 26099 27319
rect 26099 27285 26108 27319
rect 26056 27276 26108 27285
rect 26240 27276 26292 27328
rect 28080 27276 28132 27328
rect 28540 27276 28592 27328
rect 31944 27344 31996 27396
rect 36176 27344 36228 27396
rect 36820 27421 36829 27455
rect 36829 27421 36863 27455
rect 36863 27421 36872 27455
rect 36820 27412 36872 27421
rect 37280 27412 37332 27464
rect 37832 27412 37884 27464
rect 37924 27412 37976 27464
rect 39120 27412 39172 27464
rect 39856 27412 39908 27464
rect 40684 27412 40736 27464
rect 41604 27412 41656 27464
rect 41972 27455 42024 27464
rect 41972 27421 41981 27455
rect 41981 27421 42015 27455
rect 42015 27421 42024 27455
rect 41972 27412 42024 27421
rect 42524 27480 42576 27532
rect 86132 27480 86184 27532
rect 42708 27412 42760 27464
rect 42800 27455 42852 27464
rect 42800 27421 42809 27455
rect 42809 27421 42843 27455
rect 42843 27421 42852 27455
rect 43444 27455 43496 27464
rect 42800 27412 42852 27421
rect 43444 27421 43453 27455
rect 43453 27421 43487 27455
rect 43487 27421 43496 27455
rect 43444 27412 43496 27421
rect 43996 27455 44048 27464
rect 43996 27421 44005 27455
rect 44005 27421 44039 27455
rect 44039 27421 44048 27455
rect 43996 27412 44048 27421
rect 44548 27455 44600 27464
rect 44548 27421 44557 27455
rect 44557 27421 44591 27455
rect 44591 27421 44600 27455
rect 44548 27412 44600 27421
rect 45376 27455 45428 27464
rect 45376 27421 45385 27455
rect 45385 27421 45419 27455
rect 45419 27421 45428 27455
rect 45376 27412 45428 27421
rect 45468 27412 45520 27464
rect 46664 27455 46716 27464
rect 46664 27421 46673 27455
rect 46673 27421 46707 27455
rect 46707 27421 46716 27455
rect 46664 27412 46716 27421
rect 48596 27455 48648 27464
rect 48596 27421 48605 27455
rect 48605 27421 48639 27455
rect 48639 27421 48648 27455
rect 48596 27412 48648 27421
rect 49056 27412 49108 27464
rect 50528 27455 50580 27464
rect 50528 27421 50537 27455
rect 50537 27421 50571 27455
rect 50571 27421 50580 27455
rect 50528 27412 50580 27421
rect 51816 27455 51868 27464
rect 42616 27344 42668 27396
rect 46756 27344 46808 27396
rect 51172 27344 51224 27396
rect 51816 27421 51825 27455
rect 51825 27421 51859 27455
rect 51859 27421 51868 27455
rect 51816 27412 51868 27421
rect 52920 27455 52972 27464
rect 52920 27421 52929 27455
rect 52929 27421 52963 27455
rect 52963 27421 52972 27455
rect 52920 27412 52972 27421
rect 53564 27455 53616 27464
rect 53564 27421 53573 27455
rect 53573 27421 53607 27455
rect 53607 27421 53616 27455
rect 53564 27412 53616 27421
rect 54024 27412 54076 27464
rect 51724 27344 51776 27396
rect 52736 27344 52788 27396
rect 57060 27412 57112 27464
rect 58808 27455 58860 27464
rect 58808 27421 58817 27455
rect 58817 27421 58851 27455
rect 58851 27421 58860 27455
rect 58808 27412 58860 27421
rect 58624 27344 58676 27396
rect 59636 27412 59688 27464
rect 61292 27455 61344 27464
rect 61292 27421 61301 27455
rect 61301 27421 61335 27455
rect 61335 27421 61344 27455
rect 61292 27412 61344 27421
rect 61384 27412 61436 27464
rect 63868 27455 63920 27464
rect 60004 27344 60056 27396
rect 41052 27276 41104 27328
rect 41236 27319 41288 27328
rect 41236 27285 41245 27319
rect 41245 27285 41279 27319
rect 41279 27285 41288 27319
rect 41236 27276 41288 27285
rect 42892 27276 42944 27328
rect 43536 27276 43588 27328
rect 48320 27276 48372 27328
rect 50436 27276 50488 27328
rect 52092 27276 52144 27328
rect 52276 27276 52328 27328
rect 53196 27276 53248 27328
rect 54300 27276 54352 27328
rect 56968 27276 57020 27328
rect 58716 27276 58768 27328
rect 59268 27276 59320 27328
rect 60556 27276 60608 27328
rect 61568 27344 61620 27396
rect 63868 27421 63877 27455
rect 63877 27421 63911 27455
rect 63911 27421 63920 27455
rect 63868 27412 63920 27421
rect 64420 27412 64472 27464
rect 66260 27412 66312 27464
rect 66444 27412 66496 27464
rect 66996 27412 67048 27464
rect 67640 27412 67692 27464
rect 68652 27412 68704 27464
rect 69388 27412 69440 27464
rect 70860 27412 70912 27464
rect 71504 27455 71556 27464
rect 71504 27421 71513 27455
rect 71513 27421 71547 27455
rect 71547 27421 71556 27455
rect 71504 27412 71556 27421
rect 72056 27455 72108 27464
rect 72056 27421 72065 27455
rect 72065 27421 72099 27455
rect 72099 27421 72108 27455
rect 72056 27412 72108 27421
rect 73712 27455 73764 27464
rect 68192 27344 68244 27396
rect 67456 27276 67508 27328
rect 68652 27319 68704 27328
rect 68652 27285 68661 27319
rect 68661 27285 68695 27319
rect 68695 27285 68704 27319
rect 68652 27276 68704 27285
rect 69480 27344 69532 27396
rect 73712 27421 73721 27455
rect 73721 27421 73755 27455
rect 73755 27421 73764 27455
rect 73712 27412 73764 27421
rect 74448 27455 74500 27464
rect 74448 27421 74457 27455
rect 74457 27421 74491 27455
rect 74491 27421 74500 27455
rect 74448 27412 74500 27421
rect 76288 27455 76340 27464
rect 76288 27421 76297 27455
rect 76297 27421 76331 27455
rect 76331 27421 76340 27455
rect 76288 27412 76340 27421
rect 76380 27412 76432 27464
rect 69848 27276 69900 27328
rect 72516 27276 72568 27328
rect 75092 27344 75144 27396
rect 73804 27319 73856 27328
rect 73804 27285 73813 27319
rect 73813 27285 73847 27319
rect 73847 27285 73856 27319
rect 73804 27276 73856 27285
rect 75184 27276 75236 27328
rect 78312 27412 78364 27464
rect 79416 27455 79468 27464
rect 79416 27421 79425 27455
rect 79425 27421 79459 27455
rect 79459 27421 79468 27455
rect 79416 27412 79468 27421
rect 80060 27455 80112 27464
rect 80060 27421 80069 27455
rect 80069 27421 80103 27455
rect 80103 27421 80112 27455
rect 80060 27412 80112 27421
rect 81440 27455 81492 27464
rect 81440 27421 81449 27455
rect 81449 27421 81483 27455
rect 81483 27421 81492 27455
rect 81440 27412 81492 27421
rect 82176 27455 82228 27464
rect 82176 27421 82185 27455
rect 82185 27421 82219 27455
rect 82219 27421 82228 27455
rect 82176 27412 82228 27421
rect 82544 27455 82596 27464
rect 82544 27421 82553 27455
rect 82553 27421 82587 27455
rect 82587 27421 82596 27455
rect 82544 27412 82596 27421
rect 83832 27455 83884 27464
rect 83832 27421 83841 27455
rect 83841 27421 83875 27455
rect 83875 27421 83884 27455
rect 83832 27412 83884 27421
rect 84200 27412 84252 27464
rect 85120 27455 85172 27464
rect 85120 27421 85129 27455
rect 85129 27421 85163 27455
rect 85163 27421 85172 27455
rect 85120 27412 85172 27421
rect 86408 27455 86460 27464
rect 86408 27421 86417 27455
rect 86417 27421 86451 27455
rect 86451 27421 86460 27455
rect 86408 27412 86460 27421
rect 89536 27548 89588 27600
rect 87604 27480 87656 27532
rect 87788 27412 87840 27464
rect 78128 27344 78180 27396
rect 78956 27319 79008 27328
rect 78956 27285 78965 27319
rect 78965 27285 78999 27319
rect 78999 27285 79008 27319
rect 78956 27276 79008 27285
rect 79600 27319 79652 27328
rect 79600 27285 79609 27319
rect 79609 27285 79643 27319
rect 79643 27285 79652 27319
rect 79600 27276 79652 27285
rect 80244 27319 80296 27328
rect 80244 27285 80253 27319
rect 80253 27285 80287 27319
rect 80287 27285 80296 27319
rect 80244 27276 80296 27285
rect 81532 27319 81584 27328
rect 81532 27285 81541 27319
rect 81541 27285 81575 27319
rect 81575 27285 81584 27319
rect 81532 27276 81584 27285
rect 82728 27319 82780 27328
rect 82728 27285 82737 27319
rect 82737 27285 82771 27319
rect 82771 27285 82780 27319
rect 82728 27276 82780 27285
rect 87880 27276 87932 27328
rect 22898 27174 22950 27226
rect 22962 27174 23014 27226
rect 23026 27174 23078 27226
rect 23090 27174 23142 27226
rect 23154 27174 23206 27226
rect 44846 27174 44898 27226
rect 44910 27174 44962 27226
rect 44974 27174 45026 27226
rect 45038 27174 45090 27226
rect 45102 27174 45154 27226
rect 66794 27174 66846 27226
rect 66858 27174 66910 27226
rect 66922 27174 66974 27226
rect 66986 27174 67038 27226
rect 67050 27174 67102 27226
rect 20 27072 72 27124
rect 3056 27072 3108 27124
rect 3976 27115 4028 27124
rect 3976 27081 3985 27115
rect 3985 27081 4019 27115
rect 4019 27081 4028 27115
rect 3976 27072 4028 27081
rect 7288 27115 7340 27124
rect 7288 27081 7297 27115
rect 7297 27081 7331 27115
rect 7331 27081 7340 27115
rect 7288 27072 7340 27081
rect 10416 27115 10468 27124
rect 10416 27081 10425 27115
rect 10425 27081 10459 27115
rect 10459 27081 10468 27115
rect 10416 27072 10468 27081
rect 13636 27115 13688 27124
rect 13636 27081 13645 27115
rect 13645 27081 13679 27115
rect 13679 27081 13688 27115
rect 13636 27072 13688 27081
rect 18788 27072 18840 27124
rect 20352 27115 20404 27124
rect 20352 27081 20361 27115
rect 20361 27081 20395 27115
rect 20395 27081 20404 27115
rect 20352 27072 20404 27081
rect 20444 27072 20496 27124
rect 32956 27115 33008 27124
rect 1768 27047 1820 27056
rect 1768 27013 1777 27047
rect 1777 27013 1811 27047
rect 1811 27013 1820 27047
rect 1768 27004 1820 27013
rect 6736 27047 6788 27056
rect 6736 27013 6745 27047
rect 6745 27013 6779 27047
rect 6779 27013 6788 27047
rect 6736 27004 6788 27013
rect 10508 27004 10560 27056
rect 13544 27004 13596 27056
rect 2872 26936 2924 26988
rect 4160 26979 4212 26988
rect 4160 26945 4169 26979
rect 4169 26945 4203 26979
rect 4203 26945 4212 26979
rect 4160 26936 4212 26945
rect 7472 26979 7524 26988
rect 7472 26945 7481 26979
rect 7481 26945 7515 26979
rect 7515 26945 7524 26979
rect 7472 26936 7524 26945
rect 10600 26979 10652 26988
rect 10600 26945 10609 26979
rect 10609 26945 10643 26979
rect 10643 26945 10652 26979
rect 10600 26936 10652 26945
rect 12348 26979 12400 26988
rect 12348 26945 12357 26979
rect 12357 26945 12391 26979
rect 12391 26945 12400 26979
rect 12348 26936 12400 26945
rect 15660 27004 15712 27056
rect 15752 27004 15804 27056
rect 32680 27004 32732 27056
rect 32956 27081 32965 27115
rect 32965 27081 32999 27115
rect 32999 27081 33008 27115
rect 32956 27072 33008 27081
rect 33048 27072 33100 27124
rect 37556 27072 37608 27124
rect 37924 27115 37976 27124
rect 37924 27081 37933 27115
rect 37933 27081 37967 27115
rect 37967 27081 37976 27115
rect 37924 27072 37976 27081
rect 38016 27072 38068 27124
rect 40684 27115 40736 27124
rect 40684 27081 40693 27115
rect 40693 27081 40727 27115
rect 40727 27081 40736 27115
rect 40684 27072 40736 27081
rect 35532 27004 35584 27056
rect 14740 26979 14792 26988
rect 2044 26800 2096 26852
rect 6920 26843 6972 26852
rect 6920 26809 6929 26843
rect 6929 26809 6963 26843
rect 6963 26809 6972 26843
rect 6920 26800 6972 26809
rect 9680 26800 9732 26852
rect 14740 26945 14749 26979
rect 14749 26945 14783 26979
rect 14783 26945 14792 26979
rect 14740 26936 14792 26945
rect 17040 26979 17092 26988
rect 17040 26945 17049 26979
rect 17049 26945 17083 26979
rect 17083 26945 17092 26979
rect 17040 26936 17092 26945
rect 18052 26936 18104 26988
rect 19432 26936 19484 26988
rect 19984 26979 20036 26988
rect 19984 26945 19993 26979
rect 19993 26945 20027 26979
rect 20027 26945 20036 26979
rect 19984 26936 20036 26945
rect 20444 26936 20496 26988
rect 22192 26936 22244 26988
rect 23940 26936 23992 26988
rect 24124 26979 24176 26988
rect 24124 26945 24133 26979
rect 24133 26945 24167 26979
rect 24167 26945 24176 26979
rect 24124 26936 24176 26945
rect 26240 26936 26292 26988
rect 26516 26936 26568 26988
rect 27528 26936 27580 26988
rect 27712 26936 27764 26988
rect 28724 26936 28776 26988
rect 30380 26979 30432 26988
rect 30380 26945 30389 26979
rect 30389 26945 30423 26979
rect 30423 26945 30432 26979
rect 30380 26936 30432 26945
rect 12532 26775 12584 26784
rect 12532 26741 12541 26775
rect 12541 26741 12575 26775
rect 12575 26741 12584 26775
rect 12532 26732 12584 26741
rect 28264 26868 28316 26920
rect 28816 26868 28868 26920
rect 32864 26936 32916 26988
rect 33232 26936 33284 26988
rect 35256 26936 35308 26988
rect 38016 26936 38068 26988
rect 38108 26979 38160 26988
rect 38108 26945 38117 26979
rect 38117 26945 38151 26979
rect 38151 26945 38160 26979
rect 38108 26936 38160 26945
rect 38568 27004 38620 27056
rect 42524 27072 42576 27124
rect 43444 27072 43496 27124
rect 45284 27072 45336 27124
rect 50804 27072 50856 27124
rect 52736 27072 52788 27124
rect 52828 27072 52880 27124
rect 40776 26936 40828 26988
rect 40960 26936 41012 26988
rect 41052 26936 41104 26988
rect 41420 26936 41472 26988
rect 15660 26800 15712 26852
rect 21272 26800 21324 26852
rect 28172 26843 28224 26852
rect 16856 26775 16908 26784
rect 16856 26741 16865 26775
rect 16865 26741 16899 26775
rect 16899 26741 16908 26775
rect 16856 26732 16908 26741
rect 17132 26732 17184 26784
rect 23940 26775 23992 26784
rect 23940 26741 23949 26775
rect 23949 26741 23983 26775
rect 23983 26741 23992 26775
rect 23940 26732 23992 26741
rect 24032 26732 24084 26784
rect 26424 26732 26476 26784
rect 27436 26732 27488 26784
rect 28172 26809 28181 26843
rect 28181 26809 28215 26843
rect 28215 26809 28224 26843
rect 28172 26800 28224 26809
rect 29920 26800 29972 26852
rect 30012 26800 30064 26852
rect 33416 26868 33468 26920
rect 30748 26800 30800 26852
rect 38292 26868 38344 26920
rect 57060 27072 57112 27124
rect 57980 27072 58032 27124
rect 60648 27115 60700 27124
rect 60648 27081 60657 27115
rect 60657 27081 60691 27115
rect 60691 27081 60700 27115
rect 60648 27072 60700 27081
rect 53196 27004 53248 27056
rect 64880 27115 64932 27124
rect 64880 27081 64889 27115
rect 64889 27081 64923 27115
rect 64923 27081 64932 27115
rect 64880 27072 64932 27081
rect 66444 27072 66496 27124
rect 69388 27072 69440 27124
rect 71504 27072 71556 27124
rect 73160 27072 73212 27124
rect 75092 27072 75144 27124
rect 75460 27115 75512 27124
rect 75460 27081 75469 27115
rect 75469 27081 75503 27115
rect 75503 27081 75512 27115
rect 75460 27072 75512 27081
rect 83832 27072 83884 27124
rect 86316 27115 86368 27124
rect 86316 27081 86325 27115
rect 86325 27081 86359 27115
rect 86359 27081 86368 27115
rect 86316 27072 86368 27081
rect 86960 27072 87012 27124
rect 41696 26936 41748 26988
rect 44180 26936 44232 26988
rect 44732 26979 44784 26988
rect 44732 26945 44741 26979
rect 44741 26945 44775 26979
rect 44775 26945 44784 26979
rect 44732 26936 44784 26945
rect 44824 26936 44876 26988
rect 48780 26936 48832 26988
rect 49700 26936 49752 26988
rect 53932 26936 53984 26988
rect 54208 26979 54260 26988
rect 54208 26945 54217 26979
rect 54217 26945 54251 26979
rect 54251 26945 54260 26979
rect 54208 26936 54260 26945
rect 55496 26936 55548 26988
rect 58440 26979 58492 26988
rect 58440 26945 58449 26979
rect 58449 26945 58483 26979
rect 58483 26945 58492 26979
rect 58440 26936 58492 26945
rect 58992 26979 59044 26988
rect 58992 26945 59001 26979
rect 59001 26945 59035 26979
rect 59035 26945 59044 26979
rect 58992 26936 59044 26945
rect 64512 26979 64564 26988
rect 64512 26945 64521 26979
rect 64521 26945 64555 26979
rect 64555 26945 64564 26979
rect 64512 26936 64564 26945
rect 68468 27004 68520 27056
rect 81532 27004 81584 27056
rect 65616 26979 65668 26988
rect 65616 26945 65625 26979
rect 65625 26945 65659 26979
rect 65659 26945 65668 26979
rect 65616 26936 65668 26945
rect 70124 26936 70176 26988
rect 73528 26979 73580 26988
rect 73528 26945 73537 26979
rect 73537 26945 73571 26979
rect 73571 26945 73580 26979
rect 73528 26936 73580 26945
rect 73896 26936 73948 26988
rect 75644 26979 75696 26988
rect 75644 26945 75653 26979
rect 75653 26945 75687 26979
rect 75687 26945 75696 26979
rect 75644 26936 75696 26945
rect 41788 26868 41840 26920
rect 54300 26868 54352 26920
rect 54484 26911 54536 26920
rect 54484 26877 54493 26911
rect 54493 26877 54527 26911
rect 54527 26877 54536 26911
rect 54484 26868 54536 26877
rect 56968 26868 57020 26920
rect 69204 26868 69256 26920
rect 84384 26936 84436 26988
rect 85120 26936 85172 26988
rect 76748 26868 76800 26920
rect 44824 26800 44876 26852
rect 87236 26936 87288 26988
rect 87420 26911 87472 26920
rect 87420 26877 87429 26911
rect 87429 26877 87463 26911
rect 87463 26877 87472 26911
rect 87420 26868 87472 26877
rect 30472 26732 30524 26784
rect 30656 26732 30708 26784
rect 32864 26775 32916 26784
rect 32864 26741 32873 26775
rect 32873 26741 32907 26775
rect 32907 26741 32916 26775
rect 32864 26732 32916 26741
rect 41052 26732 41104 26784
rect 41420 26732 41472 26784
rect 42616 26732 42668 26784
rect 42708 26732 42760 26784
rect 49332 26732 49384 26784
rect 50344 26732 50396 26784
rect 86592 26800 86644 26852
rect 59636 26732 59688 26784
rect 68560 26732 68612 26784
rect 75644 26732 75696 26784
rect 85396 26775 85448 26784
rect 85396 26741 85405 26775
rect 85405 26741 85439 26775
rect 85439 26741 85448 26775
rect 85396 26732 85448 26741
rect 11924 26630 11976 26682
rect 11988 26630 12040 26682
rect 12052 26630 12104 26682
rect 12116 26630 12168 26682
rect 12180 26630 12232 26682
rect 33872 26630 33924 26682
rect 33936 26630 33988 26682
rect 34000 26630 34052 26682
rect 34064 26630 34116 26682
rect 34128 26630 34180 26682
rect 55820 26630 55872 26682
rect 55884 26630 55936 26682
rect 55948 26630 56000 26682
rect 56012 26630 56064 26682
rect 56076 26630 56128 26682
rect 77768 26630 77820 26682
rect 77832 26630 77884 26682
rect 77896 26630 77948 26682
rect 77960 26630 78012 26682
rect 78024 26630 78076 26682
rect 2228 26528 2280 26580
rect 12532 26528 12584 26580
rect 42708 26528 42760 26580
rect 42800 26528 42852 26580
rect 54760 26528 54812 26580
rect 55680 26528 55732 26580
rect 65064 26528 65116 26580
rect 65616 26528 65668 26580
rect 88248 26528 88300 26580
rect 14464 26460 14516 26512
rect 20076 26460 20128 26512
rect 20444 26460 20496 26512
rect 26700 26503 26752 26512
rect 18236 26392 18288 26444
rect 22008 26392 22060 26444
rect 26700 26469 26709 26503
rect 26709 26469 26743 26503
rect 26743 26469 26752 26503
rect 26700 26460 26752 26469
rect 27252 26503 27304 26512
rect 27252 26469 27261 26503
rect 27261 26469 27295 26503
rect 27295 26469 27304 26503
rect 27252 26460 27304 26469
rect 31760 26460 31812 26512
rect 35348 26460 35400 26512
rect 38292 26460 38344 26512
rect 40684 26460 40736 26512
rect 40960 26503 41012 26512
rect 40960 26469 40969 26503
rect 40969 26469 41003 26503
rect 41003 26469 41012 26503
rect 40960 26460 41012 26469
rect 41052 26460 41104 26512
rect 68560 26460 68612 26512
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 1860 26324 1912 26376
rect 3056 26367 3108 26376
rect 3056 26333 3065 26367
rect 3065 26333 3099 26367
rect 3099 26333 3108 26367
rect 3056 26324 3108 26333
rect 3976 26367 4028 26376
rect 3976 26333 3985 26367
rect 3985 26333 4019 26367
rect 4019 26333 4028 26367
rect 3976 26324 4028 26333
rect 16856 26324 16908 26376
rect 25964 26324 26016 26376
rect 27712 26392 27764 26444
rect 27436 26367 27488 26376
rect 27436 26333 27445 26367
rect 27445 26333 27479 26367
rect 27479 26333 27488 26367
rect 27436 26324 27488 26333
rect 27804 26324 27856 26376
rect 29184 26324 29236 26376
rect 29460 26324 29512 26376
rect 29644 26324 29696 26376
rect 35532 26392 35584 26444
rect 39396 26392 39448 26444
rect 43260 26392 43312 26444
rect 44824 26392 44876 26444
rect 58992 26392 59044 26444
rect 68928 26392 68980 26444
rect 82728 26392 82780 26444
rect 85396 26392 85448 26444
rect 30380 26324 30432 26376
rect 30656 26367 30708 26376
rect 30656 26333 30665 26367
rect 30665 26333 30699 26367
rect 30699 26333 30708 26367
rect 30656 26324 30708 26333
rect 31024 26367 31076 26376
rect 31024 26333 31033 26367
rect 31033 26333 31067 26367
rect 31067 26333 31076 26367
rect 31024 26324 31076 26333
rect 31300 26367 31352 26376
rect 31300 26333 31309 26367
rect 31309 26333 31343 26367
rect 31343 26333 31352 26367
rect 31300 26324 31352 26333
rect 38200 26324 38252 26376
rect 40684 26324 40736 26376
rect 40868 26324 40920 26376
rect 42616 26324 42668 26376
rect 45284 26324 45336 26376
rect 45376 26324 45428 26376
rect 55588 26324 55640 26376
rect 70124 26324 70176 26376
rect 85120 26324 85172 26376
rect 87052 26367 87104 26376
rect 87052 26333 87061 26367
rect 87061 26333 87095 26367
rect 87095 26333 87104 26367
rect 87052 26324 87104 26333
rect 87972 26367 88024 26376
rect 87972 26333 87981 26367
rect 87981 26333 88015 26367
rect 88015 26333 88024 26367
rect 87972 26324 88024 26333
rect 13544 26256 13596 26308
rect 20352 26256 20404 26308
rect 3792 26231 3844 26240
rect 3792 26197 3801 26231
rect 3801 26197 3835 26231
rect 3835 26197 3844 26231
rect 3792 26188 3844 26197
rect 19432 26188 19484 26240
rect 23388 26256 23440 26308
rect 23940 26256 23992 26308
rect 26700 26256 26752 26308
rect 25504 26188 25556 26240
rect 30012 26188 30064 26240
rect 30472 26231 30524 26240
rect 30472 26197 30481 26231
rect 30481 26197 30515 26231
rect 30515 26197 30524 26231
rect 30472 26188 30524 26197
rect 58440 26256 58492 26308
rect 40868 26188 40920 26240
rect 42064 26188 42116 26240
rect 46664 26188 46716 26240
rect 88892 26256 88944 26308
rect 88156 26231 88208 26240
rect 88156 26197 88165 26231
rect 88165 26197 88199 26231
rect 88199 26197 88208 26231
rect 88156 26188 88208 26197
rect 22898 26086 22950 26138
rect 22962 26086 23014 26138
rect 23026 26086 23078 26138
rect 23090 26086 23142 26138
rect 23154 26086 23206 26138
rect 44846 26086 44898 26138
rect 44910 26086 44962 26138
rect 44974 26086 45026 26138
rect 45038 26086 45090 26138
rect 45102 26086 45154 26138
rect 66794 26086 66846 26138
rect 66858 26086 66910 26138
rect 66922 26086 66974 26138
rect 66986 26086 67038 26138
rect 67050 26086 67102 26138
rect 1492 25984 1544 26036
rect 2780 26027 2832 26036
rect 2780 25993 2789 26027
rect 2789 25993 2823 26027
rect 2823 25993 2832 26027
rect 2780 25984 2832 25993
rect 26700 25984 26752 26036
rect 32220 25984 32272 26036
rect 44732 25984 44784 26036
rect 86132 25984 86184 26036
rect 86776 26027 86828 26036
rect 86776 25993 86785 26027
rect 86785 25993 86819 26027
rect 86819 25993 86828 26027
rect 86776 25984 86828 25993
rect 87512 26027 87564 26036
rect 87512 25993 87521 26027
rect 87521 25993 87555 26027
rect 87555 25993 87564 26027
rect 87512 25984 87564 25993
rect 87696 25984 87748 26036
rect 2596 25848 2648 25900
rect 2688 25891 2740 25900
rect 2688 25857 2697 25891
rect 2697 25857 2731 25891
rect 2731 25857 2740 25891
rect 2688 25848 2740 25857
rect 3792 25848 3844 25900
rect 88156 25916 88208 25968
rect 44640 25848 44692 25900
rect 86776 25848 86828 25900
rect 26792 25780 26844 25832
rect 35348 25780 35400 25832
rect 43260 25780 43312 25832
rect 664 25712 716 25764
rect 13084 25712 13136 25764
rect 32864 25712 32916 25764
rect 33692 25712 33744 25764
rect 58532 25712 58584 25764
rect 3148 25644 3200 25696
rect 21088 25644 21140 25696
rect 26608 25644 26660 25696
rect 87144 25687 87196 25696
rect 87144 25653 87153 25687
rect 87153 25653 87187 25687
rect 87187 25653 87196 25687
rect 87144 25644 87196 25653
rect 11924 25542 11976 25594
rect 11988 25542 12040 25594
rect 12052 25542 12104 25594
rect 12116 25542 12168 25594
rect 12180 25542 12232 25594
rect 33872 25542 33924 25594
rect 33936 25542 33988 25594
rect 34000 25542 34052 25594
rect 34064 25542 34116 25594
rect 34128 25542 34180 25594
rect 55820 25542 55872 25594
rect 55884 25542 55936 25594
rect 55948 25542 56000 25594
rect 56012 25542 56064 25594
rect 56076 25542 56128 25594
rect 77768 25542 77820 25594
rect 77832 25542 77884 25594
rect 77896 25542 77948 25594
rect 77960 25542 78012 25594
rect 78024 25542 78076 25594
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 17960 25168 18012 25220
rect 87880 25211 87932 25220
rect 87880 25177 87889 25211
rect 87889 25177 87923 25211
rect 87923 25177 87932 25211
rect 87880 25168 87932 25177
rect 87972 25143 88024 25152
rect 87972 25109 87981 25143
rect 87981 25109 88015 25143
rect 88015 25109 88024 25143
rect 87972 25100 88024 25109
rect 22898 24998 22950 25050
rect 22962 24998 23014 25050
rect 23026 24998 23078 25050
rect 23090 24998 23142 25050
rect 23154 24998 23206 25050
rect 44846 24998 44898 25050
rect 44910 24998 44962 25050
rect 44974 24998 45026 25050
rect 45038 24998 45090 25050
rect 45102 24998 45154 25050
rect 66794 24998 66846 25050
rect 66858 24998 66910 25050
rect 66922 24998 66974 25050
rect 66986 24998 67038 25050
rect 67050 24998 67102 25050
rect 88248 24803 88300 24812
rect 88248 24769 88257 24803
rect 88257 24769 88291 24803
rect 88291 24769 88300 24803
rect 88248 24760 88300 24769
rect 1400 24735 1452 24744
rect 1400 24701 1409 24735
rect 1409 24701 1443 24735
rect 1443 24701 1452 24735
rect 1400 24692 1452 24701
rect 22744 24624 22796 24676
rect 88064 24599 88116 24608
rect 88064 24565 88073 24599
rect 88073 24565 88107 24599
rect 88107 24565 88116 24599
rect 88064 24556 88116 24565
rect 11924 24454 11976 24506
rect 11988 24454 12040 24506
rect 12052 24454 12104 24506
rect 12116 24454 12168 24506
rect 12180 24454 12232 24506
rect 33872 24454 33924 24506
rect 33936 24454 33988 24506
rect 34000 24454 34052 24506
rect 34064 24454 34116 24506
rect 34128 24454 34180 24506
rect 55820 24454 55872 24506
rect 55884 24454 55936 24506
rect 55948 24454 56000 24506
rect 56012 24454 56064 24506
rect 56076 24454 56128 24506
rect 77768 24454 77820 24506
rect 77832 24454 77884 24506
rect 77896 24454 77948 24506
rect 77960 24454 78012 24506
rect 78024 24454 78076 24506
rect 53932 24216 53984 24268
rect 63408 24216 63460 24268
rect 35716 24148 35768 24200
rect 64328 24148 64380 24200
rect 86776 24148 86828 24200
rect 10600 24080 10652 24132
rect 56692 24080 56744 24132
rect 88064 24055 88116 24064
rect 88064 24021 88073 24055
rect 88073 24021 88107 24055
rect 88107 24021 88116 24055
rect 88064 24012 88116 24021
rect 22898 23910 22950 23962
rect 22962 23910 23014 23962
rect 23026 23910 23078 23962
rect 23090 23910 23142 23962
rect 23154 23910 23206 23962
rect 44846 23910 44898 23962
rect 44910 23910 44962 23962
rect 44974 23910 45026 23962
rect 45038 23910 45090 23962
rect 45102 23910 45154 23962
rect 66794 23910 66846 23962
rect 66858 23910 66910 23962
rect 66922 23910 66974 23962
rect 66986 23910 67038 23962
rect 67050 23910 67102 23962
rect 86776 23851 86828 23860
rect 86776 23817 86785 23851
rect 86785 23817 86819 23851
rect 86819 23817 86828 23851
rect 86776 23808 86828 23817
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 17960 23672 18012 23724
rect 36820 23536 36872 23588
rect 22284 23468 22336 23520
rect 73988 23468 74040 23520
rect 74448 23468 74500 23520
rect 86500 23604 86552 23656
rect 88064 23511 88116 23520
rect 88064 23477 88073 23511
rect 88073 23477 88107 23511
rect 88107 23477 88116 23511
rect 88064 23468 88116 23477
rect 11924 23366 11976 23418
rect 11988 23366 12040 23418
rect 12052 23366 12104 23418
rect 12116 23366 12168 23418
rect 12180 23366 12232 23418
rect 33872 23366 33924 23418
rect 33936 23366 33988 23418
rect 34000 23366 34052 23418
rect 34064 23366 34116 23418
rect 34128 23366 34180 23418
rect 55820 23366 55872 23418
rect 55884 23366 55936 23418
rect 55948 23366 56000 23418
rect 56012 23366 56064 23418
rect 56076 23366 56128 23418
rect 77768 23366 77820 23418
rect 77832 23366 77884 23418
rect 77896 23366 77948 23418
rect 77960 23366 78012 23418
rect 78024 23366 78076 23418
rect 4804 22924 4856 22976
rect 32312 22924 32364 22976
rect 35072 22924 35124 22976
rect 56324 22924 56376 22976
rect 22898 22822 22950 22874
rect 22962 22822 23014 22874
rect 23026 22822 23078 22874
rect 23090 22822 23142 22874
rect 23154 22822 23206 22874
rect 44846 22822 44898 22874
rect 44910 22822 44962 22874
rect 44974 22822 45026 22874
rect 45038 22822 45090 22874
rect 45102 22822 45154 22874
rect 66794 22822 66846 22874
rect 66858 22822 66910 22874
rect 66922 22822 66974 22874
rect 66986 22822 67038 22874
rect 67050 22822 67102 22874
rect 6920 22720 6972 22772
rect 36360 22720 36412 22772
rect 54484 22720 54536 22772
rect 71228 22720 71280 22772
rect 36176 22584 36228 22636
rect 38568 22584 38620 22636
rect 73436 22584 73488 22636
rect 88064 22627 88116 22636
rect 88064 22593 88073 22627
rect 88073 22593 88107 22627
rect 88107 22593 88116 22627
rect 88064 22584 88116 22593
rect 1584 22559 1636 22568
rect 1584 22525 1593 22559
rect 1593 22525 1627 22559
rect 1627 22525 1636 22559
rect 1584 22516 1636 22525
rect 86500 22380 86552 22432
rect 88156 22423 88208 22432
rect 88156 22389 88165 22423
rect 88165 22389 88199 22423
rect 88199 22389 88208 22423
rect 88156 22380 88208 22389
rect 11924 22278 11976 22330
rect 11988 22278 12040 22330
rect 12052 22278 12104 22330
rect 12116 22278 12168 22330
rect 12180 22278 12232 22330
rect 33872 22278 33924 22330
rect 33936 22278 33988 22330
rect 34000 22278 34052 22330
rect 34064 22278 34116 22330
rect 34128 22278 34180 22330
rect 55820 22278 55872 22330
rect 55884 22278 55936 22330
rect 55948 22278 56000 22330
rect 56012 22278 56064 22330
rect 56076 22278 56128 22330
rect 77768 22278 77820 22330
rect 77832 22278 77884 22330
rect 77896 22278 77948 22330
rect 77960 22278 78012 22330
rect 78024 22278 78076 22330
rect 16488 21972 16540 22024
rect 1400 21879 1452 21888
rect 1400 21845 1409 21879
rect 1409 21845 1443 21879
rect 1443 21845 1452 21879
rect 1400 21836 1452 21845
rect 87604 21836 87656 21888
rect 88064 21879 88116 21888
rect 88064 21845 88073 21879
rect 88073 21845 88107 21879
rect 88107 21845 88116 21879
rect 88064 21836 88116 21845
rect 22898 21734 22950 21786
rect 22962 21734 23014 21786
rect 23026 21734 23078 21786
rect 23090 21734 23142 21786
rect 23154 21734 23206 21786
rect 44846 21734 44898 21786
rect 44910 21734 44962 21786
rect 44974 21734 45026 21786
rect 45038 21734 45090 21786
rect 45102 21734 45154 21786
rect 66794 21734 66846 21786
rect 66858 21734 66910 21786
rect 66922 21734 66974 21786
rect 66986 21734 67038 21786
rect 67050 21734 67102 21786
rect 3976 21632 4028 21684
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 3976 21539 4028 21548
rect 3976 21505 3985 21539
rect 3985 21505 4019 21539
rect 4019 21505 4028 21539
rect 3976 21496 4028 21505
rect 4804 21428 4856 21480
rect 2596 21360 2648 21412
rect 19892 21360 19944 21412
rect 43996 21360 44048 21412
rect 63224 21360 63276 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 87512 21292 87564 21344
rect 88064 21335 88116 21344
rect 88064 21301 88073 21335
rect 88073 21301 88107 21335
rect 88107 21301 88116 21335
rect 88064 21292 88116 21301
rect 11924 21190 11976 21242
rect 11988 21190 12040 21242
rect 12052 21190 12104 21242
rect 12116 21190 12168 21242
rect 12180 21190 12232 21242
rect 33872 21190 33924 21242
rect 33936 21190 33988 21242
rect 34000 21190 34052 21242
rect 34064 21190 34116 21242
rect 34128 21190 34180 21242
rect 55820 21190 55872 21242
rect 55884 21190 55936 21242
rect 55948 21190 56000 21242
rect 56012 21190 56064 21242
rect 56076 21190 56128 21242
rect 77768 21190 77820 21242
rect 77832 21190 77884 21242
rect 77896 21190 77948 21242
rect 77960 21190 78012 21242
rect 78024 21190 78076 21242
rect 1584 21088 1636 21140
rect 57060 21088 57112 21140
rect 84844 20952 84896 21004
rect 87420 20927 87472 20936
rect 87420 20893 87429 20927
rect 87429 20893 87463 20927
rect 87463 20893 87472 20927
rect 87420 20884 87472 20893
rect 1400 20791 1452 20800
rect 1400 20757 1409 20791
rect 1409 20757 1443 20791
rect 1443 20757 1452 20791
rect 1400 20748 1452 20757
rect 1952 20791 2004 20800
rect 1952 20757 1961 20791
rect 1961 20757 1995 20791
rect 1995 20757 2004 20791
rect 1952 20748 2004 20757
rect 36820 20748 36872 20800
rect 37740 20748 37792 20800
rect 22898 20646 22950 20698
rect 22962 20646 23014 20698
rect 23026 20646 23078 20698
rect 23090 20646 23142 20698
rect 23154 20646 23206 20698
rect 44846 20646 44898 20698
rect 44910 20646 44962 20698
rect 44974 20646 45026 20698
rect 45038 20646 45090 20698
rect 45102 20646 45154 20698
rect 66794 20646 66846 20698
rect 66858 20646 66910 20698
rect 66922 20646 66974 20698
rect 66986 20646 67038 20698
rect 67050 20646 67102 20698
rect 22008 20544 22060 20596
rect 22468 20476 22520 20528
rect 25872 20476 25924 20528
rect 23756 20408 23808 20460
rect 30932 20408 30984 20460
rect 24768 20340 24820 20392
rect 88248 20204 88300 20256
rect 11924 20102 11976 20154
rect 11988 20102 12040 20154
rect 12052 20102 12104 20154
rect 12116 20102 12168 20154
rect 12180 20102 12232 20154
rect 33872 20102 33924 20154
rect 33936 20102 33988 20154
rect 34000 20102 34052 20154
rect 34064 20102 34116 20154
rect 34128 20102 34180 20154
rect 55820 20102 55872 20154
rect 55884 20102 55936 20154
rect 55948 20102 56000 20154
rect 56012 20102 56064 20154
rect 56076 20102 56128 20154
rect 77768 20102 77820 20154
rect 77832 20102 77884 20154
rect 77896 20102 77948 20154
rect 77960 20102 78012 20154
rect 78024 20102 78076 20154
rect 57152 20000 57204 20052
rect 59268 20000 59320 20052
rect 88156 20000 88208 20052
rect 38384 19932 38436 19984
rect 83740 19932 83792 19984
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 87696 19703 87748 19712
rect 87696 19669 87705 19703
rect 87705 19669 87739 19703
rect 87739 19669 87748 19703
rect 87696 19660 87748 19669
rect 88064 19703 88116 19712
rect 88064 19669 88073 19703
rect 88073 19669 88107 19703
rect 88107 19669 88116 19703
rect 88064 19660 88116 19669
rect 22898 19558 22950 19610
rect 22962 19558 23014 19610
rect 23026 19558 23078 19610
rect 23090 19558 23142 19610
rect 23154 19558 23206 19610
rect 44846 19558 44898 19610
rect 44910 19558 44962 19610
rect 44974 19558 45026 19610
rect 45038 19558 45090 19610
rect 45102 19558 45154 19610
rect 66794 19558 66846 19610
rect 66858 19558 66910 19610
rect 66922 19558 66974 19610
rect 66986 19558 67038 19610
rect 67050 19558 67102 19610
rect 63868 19456 63920 19508
rect 87696 19456 87748 19508
rect 25872 19388 25924 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 22468 19320 22520 19372
rect 24952 19320 25004 19372
rect 27988 19388 28040 19440
rect 31392 19320 31444 19372
rect 38108 19320 38160 19372
rect 56508 19363 56560 19372
rect 56508 19329 56517 19363
rect 56517 19329 56551 19363
rect 56551 19329 56560 19363
rect 56508 19320 56560 19329
rect 56600 19320 56652 19372
rect 56324 19295 56376 19304
rect 56324 19261 56333 19295
rect 56333 19261 56367 19295
rect 56367 19261 56376 19295
rect 56324 19252 56376 19261
rect 2596 19184 2648 19236
rect 27804 19184 27856 19236
rect 28080 19184 28132 19236
rect 57152 19320 57204 19372
rect 64972 19320 65024 19372
rect 4160 19116 4212 19168
rect 27896 19116 27948 19168
rect 28264 19116 28316 19168
rect 57152 19159 57204 19168
rect 57152 19125 57161 19159
rect 57161 19125 57195 19159
rect 57195 19125 57204 19159
rect 57152 19116 57204 19125
rect 88064 19159 88116 19168
rect 88064 19125 88073 19159
rect 88073 19125 88107 19159
rect 88107 19125 88116 19159
rect 88064 19116 88116 19125
rect 11924 19014 11976 19066
rect 11988 19014 12040 19066
rect 12052 19014 12104 19066
rect 12116 19014 12168 19066
rect 12180 19014 12232 19066
rect 33872 19014 33924 19066
rect 33936 19014 33988 19066
rect 34000 19014 34052 19066
rect 34064 19014 34116 19066
rect 34128 19014 34180 19066
rect 55820 19014 55872 19066
rect 55884 19014 55936 19066
rect 55948 19014 56000 19066
rect 56012 19014 56064 19066
rect 56076 19014 56128 19066
rect 77768 19014 77820 19066
rect 77832 19014 77884 19066
rect 77896 19014 77948 19066
rect 77960 19014 78012 19066
rect 78024 19014 78076 19066
rect 24584 18955 24636 18964
rect 24584 18921 24593 18955
rect 24593 18921 24627 18955
rect 24627 18921 24636 18955
rect 24584 18912 24636 18921
rect 26240 18912 26292 18964
rect 27068 18912 27120 18964
rect 33692 18912 33744 18964
rect 34520 18912 34572 18964
rect 56692 18955 56744 18964
rect 56692 18921 56701 18955
rect 56701 18921 56735 18955
rect 56735 18921 56744 18955
rect 56692 18912 56744 18921
rect 24492 18776 24544 18828
rect 34336 18844 34388 18896
rect 57704 18844 57756 18896
rect 70676 18844 70728 18896
rect 22008 18708 22060 18760
rect 24768 18751 24820 18760
rect 24768 18717 24777 18751
rect 24777 18717 24811 18751
rect 24811 18717 24820 18751
rect 24768 18708 24820 18717
rect 24952 18751 25004 18760
rect 24952 18717 24961 18751
rect 24961 18717 24995 18751
rect 24995 18717 25004 18751
rect 24952 18708 25004 18717
rect 27804 18776 27856 18828
rect 27712 18708 27764 18760
rect 48228 18776 48280 18828
rect 35992 18708 36044 18760
rect 48044 18708 48096 18760
rect 55956 18708 56008 18760
rect 56508 18708 56560 18760
rect 56968 18708 57020 18760
rect 73528 18708 73580 18760
rect 88248 18751 88300 18760
rect 88248 18717 88257 18751
rect 88257 18717 88291 18751
rect 88291 18717 88300 18751
rect 88248 18708 88300 18717
rect 1400 18615 1452 18624
rect 1400 18581 1409 18615
rect 1409 18581 1443 18615
rect 1443 18581 1452 18615
rect 1400 18572 1452 18581
rect 27896 18572 27948 18624
rect 28264 18572 28316 18624
rect 35716 18572 35768 18624
rect 39120 18640 39172 18692
rect 50160 18640 50212 18692
rect 59176 18640 59228 18692
rect 41236 18572 41288 18624
rect 47676 18572 47728 18624
rect 56232 18572 56284 18624
rect 56600 18572 56652 18624
rect 68008 18640 68060 18692
rect 71964 18640 72016 18692
rect 78956 18572 79008 18624
rect 88064 18615 88116 18624
rect 88064 18581 88073 18615
rect 88073 18581 88107 18615
rect 88107 18581 88116 18615
rect 88064 18572 88116 18581
rect 22898 18470 22950 18522
rect 22962 18470 23014 18522
rect 23026 18470 23078 18522
rect 23090 18470 23142 18522
rect 23154 18470 23206 18522
rect 44846 18470 44898 18522
rect 44910 18470 44962 18522
rect 44974 18470 45026 18522
rect 45038 18470 45090 18522
rect 45102 18470 45154 18522
rect 66794 18470 66846 18522
rect 66858 18470 66910 18522
rect 66922 18470 66974 18522
rect 66986 18470 67038 18522
rect 67050 18470 67102 18522
rect 25964 18368 26016 18420
rect 1860 18300 1912 18352
rect 12348 18232 12400 18284
rect 20812 18232 20864 18284
rect 23756 18232 23808 18284
rect 26976 18300 27028 18352
rect 27436 18232 27488 18284
rect 28540 18368 28592 18420
rect 35992 18411 36044 18420
rect 28080 18232 28132 18284
rect 28356 18275 28408 18284
rect 28356 18241 28365 18275
rect 28365 18241 28399 18275
rect 28399 18241 28408 18275
rect 28356 18232 28408 18241
rect 26240 18164 26292 18216
rect 27712 18164 27764 18216
rect 27896 18164 27948 18216
rect 35992 18377 36001 18411
rect 36001 18377 36035 18411
rect 36035 18377 36044 18411
rect 35992 18368 36044 18377
rect 43536 18368 43588 18420
rect 48044 18411 48096 18420
rect 48044 18377 48053 18411
rect 48053 18377 48087 18411
rect 48087 18377 48096 18411
rect 48044 18368 48096 18377
rect 48228 18368 48280 18420
rect 49148 18368 49200 18420
rect 49332 18411 49384 18420
rect 49332 18377 49341 18411
rect 49341 18377 49375 18411
rect 49375 18377 49384 18411
rect 49332 18368 49384 18377
rect 52920 18368 52972 18420
rect 56232 18368 56284 18420
rect 67456 18411 67508 18420
rect 67456 18377 67465 18411
rect 67465 18377 67499 18411
rect 67499 18377 67508 18411
rect 67456 18368 67508 18377
rect 36452 18343 36504 18352
rect 36452 18309 36461 18343
rect 36461 18309 36495 18343
rect 36495 18309 36504 18343
rect 36452 18300 36504 18309
rect 39488 18300 39540 18352
rect 41512 18300 41564 18352
rect 46204 18300 46256 18352
rect 34336 18275 34388 18284
rect 34336 18241 34345 18275
rect 34345 18241 34379 18275
rect 34379 18241 34388 18275
rect 34336 18232 34388 18241
rect 28632 18207 28684 18216
rect 28632 18173 28641 18207
rect 28641 18173 28675 18207
rect 28675 18173 28684 18207
rect 28632 18164 28684 18173
rect 34520 18207 34572 18216
rect 34520 18173 34529 18207
rect 34529 18173 34563 18207
rect 34563 18173 34572 18207
rect 34520 18164 34572 18173
rect 35992 18232 36044 18284
rect 36820 18232 36872 18284
rect 42432 18232 42484 18284
rect 44548 18232 44600 18284
rect 47768 18232 47820 18284
rect 48228 18232 48280 18284
rect 48872 18232 48924 18284
rect 49332 18232 49384 18284
rect 51816 18232 51868 18284
rect 54760 18300 54812 18352
rect 76380 18368 76432 18420
rect 55128 18275 55180 18284
rect 36268 18164 36320 18216
rect 36728 18164 36780 18216
rect 44272 18164 44324 18216
rect 51172 18164 51224 18216
rect 55128 18241 55137 18275
rect 55137 18241 55171 18275
rect 55171 18241 55180 18275
rect 55128 18232 55180 18241
rect 55404 18275 55456 18284
rect 55404 18241 55413 18275
rect 55413 18241 55447 18275
rect 55447 18241 55456 18275
rect 78128 18300 78180 18352
rect 55404 18232 55456 18241
rect 55956 18275 56008 18284
rect 55956 18241 55965 18275
rect 55965 18241 55999 18275
rect 55999 18241 56008 18275
rect 55956 18232 56008 18241
rect 56324 18232 56376 18284
rect 64880 18232 64932 18284
rect 69204 18232 69256 18284
rect 69756 18232 69808 18284
rect 70492 18275 70544 18284
rect 70492 18241 70501 18275
rect 70501 18241 70535 18275
rect 70535 18241 70544 18275
rect 70492 18232 70544 18241
rect 55680 18164 55732 18216
rect 7472 18096 7524 18148
rect 49608 18096 49660 18148
rect 51080 18096 51132 18148
rect 53840 18096 53892 18148
rect 1400 18071 1452 18080
rect 1400 18037 1409 18071
rect 1409 18037 1443 18071
rect 1443 18037 1452 18071
rect 1400 18028 1452 18037
rect 24952 18028 25004 18080
rect 26240 18028 26292 18080
rect 27620 18028 27672 18080
rect 27804 18028 27856 18080
rect 34980 18028 35032 18080
rect 36636 18028 36688 18080
rect 41788 18028 41840 18080
rect 45192 18028 45244 18080
rect 54392 18071 54444 18080
rect 54392 18037 54401 18071
rect 54401 18037 54435 18071
rect 54435 18037 54444 18071
rect 54392 18028 54444 18037
rect 55128 18096 55180 18148
rect 60372 18164 60424 18216
rect 60556 18164 60608 18216
rect 61384 18164 61436 18216
rect 69296 18164 69348 18216
rect 70032 18164 70084 18216
rect 70676 18207 70728 18216
rect 70676 18173 70685 18207
rect 70685 18173 70719 18207
rect 70719 18173 70728 18207
rect 70676 18164 70728 18173
rect 88064 18164 88116 18216
rect 57980 18096 58032 18148
rect 58716 18096 58768 18148
rect 67364 18096 67416 18148
rect 70216 18096 70268 18148
rect 70860 18096 70912 18148
rect 56324 18028 56376 18080
rect 62764 18028 62816 18080
rect 68100 18028 68152 18080
rect 69020 18071 69072 18080
rect 69020 18037 69029 18071
rect 69029 18037 69063 18071
rect 69063 18037 69072 18071
rect 69020 18028 69072 18037
rect 70952 18028 71004 18080
rect 11924 17926 11976 17978
rect 11988 17926 12040 17978
rect 12052 17926 12104 17978
rect 12116 17926 12168 17978
rect 12180 17926 12232 17978
rect 33872 17926 33924 17978
rect 33936 17926 33988 17978
rect 34000 17926 34052 17978
rect 34064 17926 34116 17978
rect 34128 17926 34180 17978
rect 55820 17926 55872 17978
rect 55884 17926 55936 17978
rect 55948 17926 56000 17978
rect 56012 17926 56064 17978
rect 56076 17926 56128 17978
rect 77768 17926 77820 17978
rect 77832 17926 77884 17978
rect 77896 17926 77948 17978
rect 77960 17926 78012 17978
rect 78024 17926 78076 17978
rect 1952 17824 2004 17876
rect 12532 17824 12584 17876
rect 2872 17756 2924 17808
rect 29000 17824 29052 17876
rect 2044 17688 2096 17740
rect 12440 17688 12492 17740
rect 2688 17620 2740 17672
rect 12532 17620 12584 17672
rect 12624 17620 12676 17672
rect 24952 17663 25004 17672
rect 4068 17552 4120 17604
rect 24676 17552 24728 17604
rect 12716 17484 12768 17536
rect 24584 17484 24636 17536
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 25780 17688 25832 17740
rect 27344 17731 27396 17740
rect 27344 17697 27353 17731
rect 27353 17697 27387 17731
rect 27387 17697 27396 17731
rect 27620 17731 27672 17740
rect 27344 17688 27396 17697
rect 27620 17697 27629 17731
rect 27629 17697 27663 17731
rect 27663 17697 27672 17731
rect 27620 17688 27672 17697
rect 27160 17620 27212 17672
rect 28448 17756 28500 17808
rect 31760 17756 31812 17808
rect 31944 17824 31996 17876
rect 28540 17688 28592 17740
rect 31116 17688 31168 17740
rect 31208 17688 31260 17740
rect 32404 17688 32456 17740
rect 26976 17595 27028 17604
rect 26976 17561 26985 17595
rect 26985 17561 27019 17595
rect 27019 17561 27028 17595
rect 26976 17552 27028 17561
rect 26332 17484 26384 17536
rect 28080 17484 28132 17536
rect 33600 17663 33652 17672
rect 33600 17629 33609 17663
rect 33609 17629 33643 17663
rect 33643 17629 33652 17663
rect 33600 17620 33652 17629
rect 34428 17620 34480 17672
rect 28356 17552 28408 17604
rect 31944 17552 31996 17604
rect 32128 17552 32180 17604
rect 36268 17756 36320 17808
rect 37556 17756 37608 17808
rect 40500 17756 40552 17808
rect 41512 17824 41564 17876
rect 46204 17824 46256 17876
rect 46296 17824 46348 17876
rect 48780 17867 48832 17876
rect 37832 17688 37884 17740
rect 40684 17688 40736 17740
rect 44548 17799 44600 17808
rect 41420 17688 41472 17740
rect 34704 17663 34756 17672
rect 34704 17629 34713 17663
rect 34713 17629 34747 17663
rect 34747 17629 34756 17663
rect 34704 17620 34756 17629
rect 36636 17620 36688 17672
rect 30012 17484 30064 17536
rect 30840 17484 30892 17536
rect 32496 17484 32548 17536
rect 33784 17527 33836 17536
rect 33784 17493 33793 17527
rect 33793 17493 33827 17527
rect 33827 17493 33836 17527
rect 33784 17484 33836 17493
rect 34796 17552 34848 17604
rect 34980 17595 35032 17604
rect 34980 17561 35014 17595
rect 35014 17561 35032 17595
rect 34980 17552 35032 17561
rect 41328 17620 41380 17672
rect 41512 17663 41564 17672
rect 41512 17629 41521 17663
rect 41521 17629 41555 17663
rect 41555 17629 41564 17663
rect 41512 17620 41564 17629
rect 35164 17484 35216 17536
rect 38200 17484 38252 17536
rect 40224 17484 40276 17536
rect 41420 17552 41472 17604
rect 41788 17595 41840 17604
rect 41788 17561 41822 17595
rect 41822 17561 41840 17595
rect 41788 17552 41840 17561
rect 42800 17620 42852 17672
rect 44548 17765 44557 17799
rect 44557 17765 44591 17799
rect 44591 17765 44600 17799
rect 44548 17756 44600 17765
rect 45468 17799 45520 17808
rect 45468 17765 45477 17799
rect 45477 17765 45511 17799
rect 45511 17765 45520 17799
rect 45468 17756 45520 17765
rect 48780 17833 48789 17867
rect 48789 17833 48823 17867
rect 48823 17833 48832 17867
rect 48780 17824 48832 17833
rect 50160 17867 50212 17876
rect 50160 17833 50169 17867
rect 50169 17833 50203 17867
rect 50203 17833 50212 17867
rect 50160 17824 50212 17833
rect 51080 17824 51132 17876
rect 60556 17824 60608 17876
rect 62764 17824 62816 17876
rect 70216 17824 70268 17876
rect 43444 17688 43496 17740
rect 43352 17620 43404 17672
rect 44272 17663 44324 17672
rect 44272 17629 44281 17663
rect 44281 17629 44315 17663
rect 44315 17629 44324 17663
rect 44272 17620 44324 17629
rect 48872 17688 48924 17740
rect 54300 17756 54352 17808
rect 55312 17756 55364 17808
rect 45652 17663 45704 17672
rect 45652 17629 45661 17663
rect 45661 17629 45695 17663
rect 45695 17629 45704 17663
rect 45652 17620 45704 17629
rect 45928 17663 45980 17672
rect 45928 17629 45937 17663
rect 45937 17629 45971 17663
rect 45971 17629 45980 17663
rect 45928 17620 45980 17629
rect 46940 17663 46992 17672
rect 46940 17629 46949 17663
rect 46949 17629 46983 17663
rect 46983 17629 46992 17663
rect 46940 17620 46992 17629
rect 47216 17663 47268 17672
rect 47216 17629 47225 17663
rect 47225 17629 47259 17663
rect 47259 17629 47268 17663
rect 47216 17620 47268 17629
rect 48136 17663 48188 17672
rect 46572 17552 46624 17604
rect 41696 17484 41748 17536
rect 47860 17552 47912 17604
rect 48136 17629 48145 17663
rect 48145 17629 48179 17663
rect 48179 17629 48188 17663
rect 48136 17620 48188 17629
rect 48228 17620 48280 17672
rect 49148 17663 49200 17672
rect 49148 17629 49157 17663
rect 49157 17629 49191 17663
rect 49191 17629 49200 17663
rect 49148 17620 49200 17629
rect 49240 17663 49292 17672
rect 49240 17629 49249 17663
rect 49249 17629 49283 17663
rect 49283 17629 49292 17663
rect 53012 17688 53064 17740
rect 53104 17688 53156 17740
rect 55404 17688 55456 17740
rect 49240 17620 49292 17629
rect 50528 17620 50580 17672
rect 52184 17620 52236 17672
rect 53288 17663 53340 17672
rect 53288 17629 53297 17663
rect 53297 17629 53331 17663
rect 53331 17629 53340 17663
rect 53288 17620 53340 17629
rect 53932 17620 53984 17672
rect 54116 17663 54168 17672
rect 54116 17629 54125 17663
rect 54125 17629 54159 17663
rect 54159 17629 54168 17663
rect 54116 17620 54168 17629
rect 54576 17620 54628 17672
rect 54668 17620 54720 17672
rect 55312 17663 55364 17672
rect 55312 17629 55321 17663
rect 55321 17629 55355 17663
rect 55355 17629 55364 17663
rect 55312 17620 55364 17629
rect 56416 17756 56468 17808
rect 60464 17756 60516 17808
rect 60648 17756 60700 17808
rect 61016 17756 61068 17808
rect 61108 17756 61160 17808
rect 64512 17756 64564 17808
rect 65524 17756 65576 17808
rect 68468 17756 68520 17808
rect 55680 17731 55732 17740
rect 55680 17697 55689 17731
rect 55689 17697 55723 17731
rect 55723 17697 55732 17731
rect 55680 17688 55732 17697
rect 55588 17620 55640 17672
rect 56048 17663 56100 17672
rect 56048 17629 56057 17663
rect 56057 17629 56091 17663
rect 56091 17629 56100 17663
rect 56048 17620 56100 17629
rect 56324 17620 56376 17672
rect 53104 17552 53156 17604
rect 58716 17663 58768 17672
rect 58716 17629 58725 17663
rect 58725 17629 58759 17663
rect 58759 17629 58768 17663
rect 58716 17620 58768 17629
rect 58992 17663 59044 17672
rect 58992 17629 59001 17663
rect 59001 17629 59035 17663
rect 59035 17629 59044 17663
rect 58992 17620 59044 17629
rect 59268 17620 59320 17672
rect 59912 17620 59964 17672
rect 60832 17688 60884 17740
rect 61568 17620 61620 17672
rect 62764 17688 62816 17740
rect 62396 17663 62448 17672
rect 62396 17629 62405 17663
rect 62405 17629 62439 17663
rect 62439 17629 62448 17663
rect 62396 17620 62448 17629
rect 62488 17620 62540 17672
rect 65156 17663 65208 17672
rect 65156 17629 65165 17663
rect 65165 17629 65199 17663
rect 65199 17629 65208 17663
rect 65156 17620 65208 17629
rect 68100 17663 68152 17672
rect 68100 17629 68109 17663
rect 68109 17629 68143 17663
rect 68143 17629 68152 17663
rect 68100 17620 68152 17629
rect 68468 17620 68520 17672
rect 69204 17688 69256 17740
rect 69664 17620 69716 17672
rect 70952 17663 71004 17672
rect 70952 17629 70961 17663
rect 70961 17629 70995 17663
rect 70995 17629 71004 17663
rect 70952 17620 71004 17629
rect 47400 17484 47452 17536
rect 48964 17484 49016 17536
rect 49148 17484 49200 17536
rect 53380 17527 53432 17536
rect 53380 17493 53395 17527
rect 53395 17493 53429 17527
rect 53429 17493 53432 17527
rect 53380 17484 53432 17493
rect 53564 17484 53616 17536
rect 53656 17484 53708 17536
rect 56416 17484 56468 17536
rect 56600 17484 56652 17536
rect 59084 17484 59136 17536
rect 59360 17552 59412 17604
rect 60648 17552 60700 17604
rect 60832 17595 60884 17604
rect 60832 17561 60841 17595
rect 60841 17561 60875 17595
rect 60875 17561 60884 17595
rect 60832 17552 60884 17561
rect 59728 17484 59780 17536
rect 60372 17484 60424 17536
rect 60924 17527 60976 17536
rect 60924 17493 60933 17527
rect 60933 17493 60967 17527
rect 60967 17493 60976 17527
rect 60924 17484 60976 17493
rect 61016 17484 61068 17536
rect 62120 17552 62172 17604
rect 62580 17527 62632 17536
rect 62580 17493 62589 17527
rect 62589 17493 62623 17527
rect 62623 17493 62632 17527
rect 62580 17484 62632 17493
rect 65524 17552 65576 17604
rect 66720 17484 66772 17536
rect 68284 17552 68336 17604
rect 68560 17552 68612 17604
rect 75184 17552 75236 17604
rect 69572 17484 69624 17536
rect 70492 17484 70544 17536
rect 70768 17527 70820 17536
rect 70768 17493 70777 17527
rect 70777 17493 70811 17527
rect 70811 17493 70820 17527
rect 70768 17484 70820 17493
rect 22898 17382 22950 17434
rect 22962 17382 23014 17434
rect 23026 17382 23078 17434
rect 23090 17382 23142 17434
rect 23154 17382 23206 17434
rect 44846 17382 44898 17434
rect 44910 17382 44962 17434
rect 44974 17382 45026 17434
rect 45038 17382 45090 17434
rect 45102 17382 45154 17434
rect 66794 17382 66846 17434
rect 66858 17382 66910 17434
rect 66922 17382 66974 17434
rect 66986 17382 67038 17434
rect 67050 17382 67102 17434
rect 12440 17280 12492 17332
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 22376 17212 22428 17264
rect 22744 17280 22796 17332
rect 28356 17280 28408 17332
rect 30012 17280 30064 17332
rect 24676 17212 24728 17264
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 24952 17187 25004 17196
rect 24952 17153 24961 17187
rect 24961 17153 24995 17187
rect 24995 17153 25004 17187
rect 24952 17144 25004 17153
rect 26240 17187 26292 17196
rect 26240 17153 26249 17187
rect 26249 17153 26283 17187
rect 26283 17153 26292 17187
rect 26240 17144 26292 17153
rect 27804 17212 27856 17264
rect 32128 17212 32180 17264
rect 32220 17212 32272 17264
rect 32772 17212 32824 17264
rect 35716 17255 35768 17264
rect 28080 17144 28132 17196
rect 24216 17119 24268 17128
rect 24216 17085 24225 17119
rect 24225 17085 24259 17119
rect 24259 17085 24268 17119
rect 24676 17119 24728 17128
rect 24216 17076 24268 17085
rect 24676 17085 24685 17119
rect 24685 17085 24719 17119
rect 24719 17085 24728 17119
rect 24676 17076 24728 17085
rect 26976 17076 27028 17128
rect 27252 17119 27304 17128
rect 27252 17085 27261 17119
rect 27261 17085 27295 17119
rect 27295 17085 27304 17119
rect 27252 17076 27304 17085
rect 24952 17008 25004 17060
rect 28356 17076 28408 17128
rect 31760 17076 31812 17128
rect 32680 17144 32732 17196
rect 33600 17187 33652 17196
rect 33600 17153 33609 17187
rect 33609 17153 33643 17187
rect 33643 17153 33652 17187
rect 33600 17144 33652 17153
rect 33784 17187 33836 17196
rect 33784 17153 33793 17187
rect 33793 17153 33827 17187
rect 33827 17153 33836 17187
rect 33784 17144 33836 17153
rect 35716 17221 35750 17255
rect 35750 17221 35768 17255
rect 35716 17212 35768 17221
rect 37832 17255 37884 17264
rect 37832 17221 37841 17255
rect 37841 17221 37875 17255
rect 37875 17221 37884 17255
rect 37832 17212 37884 17221
rect 32036 17076 32088 17128
rect 25688 16940 25740 16992
rect 26240 16940 26292 16992
rect 28540 16940 28592 16992
rect 31484 16983 31536 16992
rect 31484 16949 31493 16983
rect 31493 16949 31527 16983
rect 31527 16949 31536 16983
rect 31484 16940 31536 16949
rect 32404 17076 32456 17128
rect 32772 17119 32824 17128
rect 32772 17085 32781 17119
rect 32781 17085 32815 17119
rect 32815 17085 32824 17119
rect 32772 17076 32824 17085
rect 37556 17144 37608 17196
rect 37648 17187 37700 17196
rect 37648 17153 37657 17187
rect 37657 17153 37691 17187
rect 37691 17153 37700 17187
rect 39488 17212 39540 17264
rect 38200 17187 38252 17196
rect 37648 17144 37700 17153
rect 38200 17153 38209 17187
rect 38209 17153 38243 17187
rect 38243 17153 38252 17187
rect 38200 17144 38252 17153
rect 41512 17212 41564 17264
rect 41880 17212 41932 17264
rect 42892 17255 42944 17264
rect 42892 17221 42901 17255
rect 42901 17221 42935 17255
rect 42935 17221 42944 17255
rect 42892 17212 42944 17221
rect 40132 17144 40184 17196
rect 41236 17187 41288 17196
rect 41236 17153 41245 17187
rect 41245 17153 41279 17187
rect 41279 17153 41288 17187
rect 41788 17187 41840 17196
rect 41236 17144 41288 17153
rect 41788 17153 41797 17187
rect 41797 17153 41831 17187
rect 41831 17153 41840 17187
rect 41788 17144 41840 17153
rect 42248 17144 42300 17196
rect 42800 17187 42852 17196
rect 34336 17076 34388 17128
rect 35440 17119 35492 17128
rect 35440 17085 35449 17119
rect 35449 17085 35483 17119
rect 35483 17085 35492 17119
rect 35440 17076 35492 17085
rect 33048 17008 33100 17060
rect 34704 17008 34756 17060
rect 36452 17008 36504 17060
rect 39580 17008 39632 17060
rect 41420 17008 41472 17060
rect 41696 17076 41748 17128
rect 42800 17153 42809 17187
rect 42809 17153 42843 17187
rect 42843 17153 42852 17187
rect 42800 17144 42852 17153
rect 43628 17144 43680 17196
rect 44732 17212 44784 17264
rect 45744 17212 45796 17264
rect 45100 17187 45152 17196
rect 45100 17153 45134 17187
rect 45134 17153 45152 17187
rect 42432 17051 42484 17060
rect 36820 16983 36872 16992
rect 36820 16949 36829 16983
rect 36829 16949 36863 16983
rect 36863 16949 36872 16983
rect 36820 16940 36872 16949
rect 40316 16940 40368 16992
rect 41512 16940 41564 16992
rect 42432 17017 42441 17051
rect 42441 17017 42475 17051
rect 42475 17017 42484 17051
rect 42432 17008 42484 17017
rect 43076 17076 43128 17128
rect 45100 17144 45152 17153
rect 46572 17187 46624 17196
rect 46572 17153 46581 17187
rect 46581 17153 46615 17187
rect 46615 17153 46624 17187
rect 46572 17144 46624 17153
rect 46756 17187 46808 17196
rect 46756 17153 46765 17187
rect 46765 17153 46799 17187
rect 46799 17153 46808 17187
rect 46756 17144 46808 17153
rect 47032 17187 47084 17196
rect 47032 17153 47041 17187
rect 47041 17153 47075 17187
rect 47075 17153 47084 17187
rect 47952 17212 48004 17264
rect 53656 17255 53708 17264
rect 47032 17144 47084 17153
rect 47676 17144 47728 17196
rect 48320 17144 48372 17196
rect 48780 17144 48832 17196
rect 49700 17187 49752 17196
rect 49700 17153 49709 17187
rect 49709 17153 49743 17187
rect 49743 17153 49752 17187
rect 49700 17144 49752 17153
rect 49884 17187 49936 17196
rect 49884 17153 49893 17187
rect 49893 17153 49927 17187
rect 49927 17153 49936 17187
rect 49884 17144 49936 17153
rect 50528 17144 50580 17196
rect 50804 17187 50856 17196
rect 50804 17153 50813 17187
rect 50813 17153 50847 17187
rect 50847 17153 50856 17187
rect 50804 17144 50856 17153
rect 43352 16940 43404 16992
rect 43628 16940 43680 16992
rect 43812 17008 43864 17060
rect 44824 17008 44876 17060
rect 46296 17008 46348 17060
rect 46848 16940 46900 16992
rect 49424 17076 49476 17128
rect 50160 17076 50212 17128
rect 51080 17076 51132 17128
rect 48964 17051 49016 17060
rect 48964 17017 48973 17051
rect 48973 17017 49007 17051
rect 49007 17017 49016 17051
rect 48964 17008 49016 17017
rect 49608 17008 49660 17060
rect 49976 17008 50028 17060
rect 50804 16940 50856 16992
rect 50988 16940 51040 16992
rect 51356 16983 51408 16992
rect 51356 16949 51365 16983
rect 51365 16949 51399 16983
rect 51399 16949 51408 16983
rect 53656 17221 53665 17255
rect 53665 17221 53699 17255
rect 53699 17221 53708 17255
rect 53656 17212 53708 17221
rect 53472 17187 53524 17196
rect 53472 17153 53481 17187
rect 53481 17153 53515 17187
rect 53515 17153 53524 17187
rect 54208 17212 54260 17264
rect 54392 17255 54444 17264
rect 54392 17221 54426 17255
rect 54426 17221 54444 17255
rect 54392 17212 54444 17221
rect 54484 17212 54536 17264
rect 53472 17144 53524 17153
rect 53932 17144 53984 17196
rect 53748 17008 53800 17060
rect 53840 17008 53892 17060
rect 51356 16940 51408 16949
rect 53932 16940 53984 16992
rect 55312 17076 55364 17128
rect 56048 17076 56100 17128
rect 56324 17187 56376 17196
rect 56324 17153 56333 17187
rect 56333 17153 56367 17187
rect 56367 17153 56376 17187
rect 56324 17144 56376 17153
rect 56784 17144 56836 17196
rect 57704 17144 57756 17196
rect 57888 17187 57940 17196
rect 57888 17153 57897 17187
rect 57897 17153 57931 17187
rect 57931 17153 57940 17187
rect 57888 17144 57940 17153
rect 58072 17187 58124 17196
rect 58072 17153 58081 17187
rect 58081 17153 58115 17187
rect 58115 17153 58124 17187
rect 58072 17144 58124 17153
rect 58164 17187 58216 17196
rect 58164 17153 58173 17187
rect 58173 17153 58207 17187
rect 58207 17153 58216 17187
rect 58532 17212 58584 17264
rect 59912 17255 59964 17264
rect 59912 17221 59921 17255
rect 59921 17221 59955 17255
rect 59955 17221 59964 17255
rect 59912 17212 59964 17221
rect 58164 17144 58216 17153
rect 58808 17144 58860 17196
rect 58900 17187 58952 17196
rect 58900 17153 58909 17187
rect 58909 17153 58943 17187
rect 58943 17153 58952 17187
rect 58900 17144 58952 17153
rect 58624 17076 58676 17128
rect 59268 17076 59320 17128
rect 59544 17119 59596 17128
rect 59544 17085 59553 17119
rect 59553 17085 59587 17119
rect 59587 17085 59596 17119
rect 59544 17076 59596 17085
rect 59728 17187 59780 17196
rect 59728 17153 59737 17187
rect 59737 17153 59771 17187
rect 59771 17153 59780 17187
rect 62672 17212 62724 17264
rect 64420 17212 64472 17264
rect 59728 17144 59780 17153
rect 60372 17144 60424 17196
rect 62120 17187 62172 17196
rect 62120 17153 62129 17187
rect 62129 17153 62163 17187
rect 62163 17153 62172 17187
rect 62120 17144 62172 17153
rect 62396 17144 62448 17196
rect 63500 17187 63552 17196
rect 63500 17153 63509 17187
rect 63509 17153 63543 17187
rect 63543 17153 63552 17187
rect 63500 17144 63552 17153
rect 63684 17144 63736 17196
rect 64788 17144 64840 17196
rect 64972 17187 65024 17196
rect 64972 17153 64981 17187
rect 64981 17153 65015 17187
rect 65015 17153 65024 17187
rect 64972 17144 65024 17153
rect 59820 17076 59872 17128
rect 60004 17076 60056 17128
rect 61384 17076 61436 17128
rect 64696 17076 64748 17128
rect 69388 17212 69440 17264
rect 70676 17212 70728 17264
rect 66720 17144 66772 17196
rect 66996 17187 67048 17196
rect 66996 17153 67005 17187
rect 67005 17153 67039 17187
rect 67039 17153 67048 17187
rect 66996 17144 67048 17153
rect 69020 17144 69072 17196
rect 69112 17144 69164 17196
rect 55128 17008 55180 17060
rect 56324 17008 56376 17060
rect 60280 17008 60332 17060
rect 66444 17119 66496 17128
rect 55220 16940 55272 16992
rect 55312 16940 55364 16992
rect 56508 16983 56560 16992
rect 56508 16949 56517 16983
rect 56517 16949 56551 16983
rect 56551 16949 56560 16983
rect 56508 16940 56560 16949
rect 59268 16940 59320 16992
rect 60648 16940 60700 16992
rect 65156 17008 65208 17060
rect 66444 17085 66453 17119
rect 66453 17085 66487 17119
rect 66487 17085 66496 17119
rect 66444 17076 66496 17085
rect 66536 17076 66588 17128
rect 69664 17119 69716 17128
rect 61660 16983 61712 16992
rect 61660 16949 61669 16983
rect 61669 16949 61703 16983
rect 61703 16949 61712 16983
rect 61660 16940 61712 16949
rect 62580 16940 62632 16992
rect 64236 16940 64288 16992
rect 65340 16940 65392 16992
rect 68560 17008 68612 17060
rect 68652 17008 68704 17060
rect 69664 17085 69673 17119
rect 69673 17085 69707 17119
rect 69707 17085 69716 17119
rect 69664 17076 69716 17085
rect 70768 17144 70820 17196
rect 87604 17212 87656 17264
rect 70400 17076 70452 17128
rect 70584 17076 70636 17128
rect 71320 17076 71372 17128
rect 87052 17008 87104 17060
rect 88064 17051 88116 17060
rect 88064 17017 88073 17051
rect 88073 17017 88107 17051
rect 88107 17017 88116 17051
rect 88064 17008 88116 17017
rect 11924 16838 11976 16890
rect 11988 16838 12040 16890
rect 12052 16838 12104 16890
rect 12116 16838 12168 16890
rect 12180 16838 12232 16890
rect 33872 16838 33924 16890
rect 33936 16838 33988 16890
rect 34000 16838 34052 16890
rect 34064 16838 34116 16890
rect 34128 16838 34180 16890
rect 55820 16838 55872 16890
rect 55884 16838 55936 16890
rect 55948 16838 56000 16890
rect 56012 16838 56064 16890
rect 56076 16838 56128 16890
rect 77768 16838 77820 16890
rect 77832 16838 77884 16890
rect 77896 16838 77948 16890
rect 77960 16838 78012 16890
rect 78024 16838 78076 16890
rect 20076 16779 20128 16788
rect 20076 16745 20085 16779
rect 20085 16745 20119 16779
rect 20119 16745 20128 16779
rect 20076 16736 20128 16745
rect 21088 16736 21140 16788
rect 21640 16736 21692 16788
rect 61384 16736 61436 16788
rect 61568 16736 61620 16788
rect 62396 16736 62448 16788
rect 63500 16736 63552 16788
rect 64328 16736 64380 16788
rect 28724 16668 28776 16720
rect 32772 16668 32824 16720
rect 36452 16668 36504 16720
rect 2964 16532 3016 16584
rect 20536 16575 20588 16584
rect 20536 16541 20545 16575
rect 20545 16541 20579 16575
rect 20579 16541 20588 16575
rect 25780 16600 25832 16652
rect 28172 16600 28224 16652
rect 32864 16600 32916 16652
rect 21364 16575 21416 16584
rect 20536 16532 20588 16541
rect 21364 16541 21373 16575
rect 21373 16541 21407 16575
rect 21407 16541 21416 16575
rect 21364 16532 21416 16541
rect 21640 16575 21692 16584
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 25964 16532 26016 16584
rect 26332 16575 26384 16584
rect 26332 16541 26366 16575
rect 26366 16541 26384 16575
rect 26332 16532 26384 16541
rect 28448 16575 28500 16584
rect 28448 16541 28457 16575
rect 28457 16541 28491 16575
rect 28491 16541 28500 16575
rect 28448 16532 28500 16541
rect 30840 16575 30892 16584
rect 30840 16541 30849 16575
rect 30849 16541 30883 16575
rect 30883 16541 30892 16575
rect 30840 16532 30892 16541
rect 31116 16532 31168 16584
rect 33324 16532 33376 16584
rect 33784 16600 33836 16652
rect 36360 16643 36412 16652
rect 36360 16609 36369 16643
rect 36369 16609 36403 16643
rect 36403 16609 36412 16643
rect 36360 16600 36412 16609
rect 36728 16668 36780 16720
rect 36820 16600 36872 16652
rect 35900 16532 35952 16584
rect 38200 16532 38252 16584
rect 26148 16464 26200 16516
rect 1400 16439 1452 16448
rect 1400 16405 1409 16439
rect 1409 16405 1443 16439
rect 1443 16405 1452 16439
rect 1400 16396 1452 16405
rect 25320 16396 25372 16448
rect 25596 16396 25648 16448
rect 28632 16464 28684 16516
rect 31484 16507 31536 16516
rect 31484 16473 31518 16507
rect 31518 16473 31536 16507
rect 31484 16464 31536 16473
rect 27436 16439 27488 16448
rect 27436 16405 27445 16439
rect 27445 16405 27479 16439
rect 27479 16405 27488 16439
rect 27436 16396 27488 16405
rect 29184 16396 29236 16448
rect 29736 16396 29788 16448
rect 30656 16439 30708 16448
rect 30656 16405 30665 16439
rect 30665 16405 30699 16439
rect 30699 16405 30708 16439
rect 30656 16396 30708 16405
rect 30748 16396 30800 16448
rect 32864 16464 32916 16516
rect 34704 16464 34756 16516
rect 38752 16600 38804 16652
rect 40132 16668 40184 16720
rect 40316 16668 40368 16720
rect 41696 16668 41748 16720
rect 42984 16668 43036 16720
rect 45928 16668 45980 16720
rect 46940 16668 46992 16720
rect 47768 16711 47820 16720
rect 47768 16677 47777 16711
rect 47777 16677 47811 16711
rect 47811 16677 47820 16711
rect 47768 16668 47820 16677
rect 47860 16668 47912 16720
rect 50068 16668 50120 16720
rect 51264 16668 51316 16720
rect 52828 16668 52880 16720
rect 55128 16668 55180 16720
rect 58716 16668 58768 16720
rect 59268 16668 59320 16720
rect 62028 16668 62080 16720
rect 63040 16668 63092 16720
rect 64144 16668 64196 16720
rect 64788 16668 64840 16720
rect 40224 16575 40276 16584
rect 40224 16541 40233 16575
rect 40233 16541 40267 16575
rect 40267 16541 40276 16575
rect 40224 16532 40276 16541
rect 41512 16575 41564 16584
rect 41512 16541 41521 16575
rect 41521 16541 41555 16575
rect 41555 16541 41564 16575
rect 41512 16532 41564 16541
rect 41696 16532 41748 16584
rect 41880 16575 41932 16584
rect 41880 16541 41889 16575
rect 41889 16541 41923 16575
rect 41923 16541 41932 16575
rect 41880 16532 41932 16541
rect 42708 16532 42760 16584
rect 47032 16600 47084 16652
rect 48228 16600 48280 16652
rect 49792 16600 49844 16652
rect 51172 16600 51224 16652
rect 53472 16600 53524 16652
rect 32680 16396 32732 16448
rect 33140 16439 33192 16448
rect 33140 16405 33149 16439
rect 33149 16405 33183 16439
rect 33183 16405 33192 16439
rect 33140 16396 33192 16405
rect 35532 16396 35584 16448
rect 35992 16396 36044 16448
rect 37556 16396 37608 16448
rect 38660 16439 38712 16448
rect 38660 16405 38669 16439
rect 38669 16405 38703 16439
rect 38703 16405 38712 16439
rect 38660 16396 38712 16405
rect 46756 16532 46808 16584
rect 46848 16575 46900 16584
rect 46848 16541 46857 16575
rect 46857 16541 46891 16575
rect 46891 16541 46900 16575
rect 47216 16575 47268 16584
rect 46848 16532 46900 16541
rect 47216 16541 47225 16575
rect 47225 16541 47259 16575
rect 47259 16541 47268 16575
rect 47216 16532 47268 16541
rect 47400 16575 47452 16584
rect 47400 16541 47409 16575
rect 47409 16541 47443 16575
rect 47443 16541 47452 16575
rect 47400 16532 47452 16541
rect 47584 16575 47636 16584
rect 47584 16541 47598 16575
rect 47598 16541 47632 16575
rect 47632 16541 47636 16575
rect 47584 16532 47636 16541
rect 50252 16532 50304 16584
rect 51356 16532 51408 16584
rect 52368 16575 52420 16584
rect 52368 16541 52377 16575
rect 52377 16541 52411 16575
rect 52411 16541 52420 16575
rect 52368 16532 52420 16541
rect 52552 16575 52604 16584
rect 52552 16541 52561 16575
rect 52561 16541 52595 16575
rect 52595 16541 52604 16575
rect 52552 16532 52604 16541
rect 52736 16575 52788 16584
rect 52736 16541 52750 16575
rect 52750 16541 52784 16575
rect 52784 16541 52788 16575
rect 53380 16575 53432 16584
rect 52736 16532 52788 16541
rect 53380 16541 53389 16575
rect 53389 16541 53423 16575
rect 53423 16541 53432 16575
rect 53380 16532 53432 16541
rect 41788 16396 41840 16448
rect 43168 16396 43220 16448
rect 43352 16396 43404 16448
rect 44732 16464 44784 16516
rect 47124 16464 47176 16516
rect 47308 16464 47360 16516
rect 50896 16464 50948 16516
rect 50988 16464 51040 16516
rect 51080 16464 51132 16516
rect 44824 16396 44876 16448
rect 46664 16396 46716 16448
rect 47768 16396 47820 16448
rect 48228 16396 48280 16448
rect 50252 16396 50304 16448
rect 50344 16396 50396 16448
rect 51448 16396 51500 16448
rect 52000 16464 52052 16516
rect 52460 16464 52512 16516
rect 53104 16464 53156 16516
rect 51632 16396 51684 16448
rect 53932 16532 53984 16584
rect 54760 16575 54812 16584
rect 54116 16464 54168 16516
rect 54392 16464 54444 16516
rect 54760 16541 54769 16575
rect 54769 16541 54803 16575
rect 54803 16541 54812 16575
rect 54760 16532 54812 16541
rect 55220 16600 55272 16652
rect 58900 16600 58952 16652
rect 59912 16600 59964 16652
rect 56508 16532 56560 16584
rect 55312 16464 55364 16516
rect 56600 16464 56652 16516
rect 56876 16464 56928 16516
rect 57888 16464 57940 16516
rect 58440 16507 58492 16516
rect 54300 16396 54352 16448
rect 56416 16396 56468 16448
rect 56784 16396 56836 16448
rect 57336 16396 57388 16448
rect 58440 16473 58449 16507
rect 58449 16473 58483 16507
rect 58483 16473 58492 16507
rect 58440 16464 58492 16473
rect 58532 16439 58584 16448
rect 58532 16405 58547 16439
rect 58547 16405 58581 16439
rect 58581 16405 58584 16439
rect 58532 16396 58584 16405
rect 60832 16532 60884 16584
rect 61016 16532 61068 16584
rect 61108 16575 61160 16584
rect 61108 16541 61117 16575
rect 61117 16541 61151 16575
rect 61151 16541 61160 16575
rect 61108 16532 61160 16541
rect 59084 16464 59136 16516
rect 59268 16464 59320 16516
rect 60096 16464 60148 16516
rect 60740 16464 60792 16516
rect 61200 16464 61252 16516
rect 62580 16532 62632 16584
rect 62764 16575 62816 16584
rect 62764 16541 62773 16575
rect 62773 16541 62807 16575
rect 62807 16541 62816 16575
rect 62764 16532 62816 16541
rect 65248 16600 65300 16652
rect 65524 16600 65576 16652
rect 68560 16736 68612 16788
rect 87328 16736 87380 16788
rect 69388 16668 69440 16720
rect 77116 16668 77168 16720
rect 71136 16643 71188 16652
rect 60188 16396 60240 16448
rect 60648 16439 60700 16448
rect 60648 16405 60657 16439
rect 60657 16405 60691 16439
rect 60691 16405 60700 16439
rect 61660 16464 61712 16516
rect 63132 16464 63184 16516
rect 65340 16532 65392 16584
rect 71136 16609 71145 16643
rect 71145 16609 71179 16643
rect 71179 16609 71188 16643
rect 71136 16600 71188 16609
rect 73068 16600 73120 16652
rect 68928 16532 68980 16584
rect 70768 16532 70820 16584
rect 71320 16575 71372 16584
rect 71320 16541 71329 16575
rect 71329 16541 71363 16575
rect 71363 16541 71372 16575
rect 71320 16532 71372 16541
rect 87880 16532 87932 16584
rect 68652 16507 68704 16516
rect 63316 16439 63368 16448
rect 60648 16396 60700 16405
rect 63316 16405 63325 16439
rect 63325 16405 63359 16439
rect 63359 16405 63368 16439
rect 63316 16396 63368 16405
rect 65340 16396 65392 16448
rect 65984 16396 66036 16448
rect 68652 16473 68686 16507
rect 68686 16473 68704 16507
rect 68652 16464 68704 16473
rect 68376 16396 68428 16448
rect 68560 16396 68612 16448
rect 69756 16439 69808 16448
rect 69756 16405 69765 16439
rect 69765 16405 69799 16439
rect 69799 16405 69808 16439
rect 69756 16396 69808 16405
rect 70124 16439 70176 16448
rect 70124 16405 70133 16439
rect 70133 16405 70167 16439
rect 70167 16405 70176 16439
rect 70124 16396 70176 16405
rect 88064 16439 88116 16448
rect 88064 16405 88073 16439
rect 88073 16405 88107 16439
rect 88107 16405 88116 16439
rect 88064 16396 88116 16405
rect 22898 16294 22950 16346
rect 22962 16294 23014 16346
rect 23026 16294 23078 16346
rect 23090 16294 23142 16346
rect 23154 16294 23206 16346
rect 44846 16294 44898 16346
rect 44910 16294 44962 16346
rect 44974 16294 45026 16346
rect 45038 16294 45090 16346
rect 45102 16294 45154 16346
rect 66794 16294 66846 16346
rect 66858 16294 66910 16346
rect 66922 16294 66974 16346
rect 66986 16294 67038 16346
rect 67050 16294 67102 16346
rect 2964 16235 3016 16244
rect 2964 16201 2973 16235
rect 2973 16201 3007 16235
rect 3007 16201 3016 16235
rect 2964 16192 3016 16201
rect 20260 16192 20312 16244
rect 22560 16192 22612 16244
rect 24584 16192 24636 16244
rect 25596 16192 25648 16244
rect 26240 16192 26292 16244
rect 30748 16192 30800 16244
rect 34704 16235 34756 16244
rect 21364 16124 21416 16176
rect 25320 16167 25372 16176
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 21916 16056 21968 16108
rect 22192 16099 22244 16108
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22192 16056 22244 16065
rect 22744 16056 22796 16108
rect 24768 16056 24820 16108
rect 25044 16099 25096 16108
rect 25044 16065 25053 16099
rect 25053 16065 25087 16099
rect 25087 16065 25096 16099
rect 25044 16056 25096 16065
rect 25320 16133 25354 16167
rect 25354 16133 25372 16167
rect 25320 16124 25372 16133
rect 30472 16124 30524 16176
rect 30840 16124 30892 16176
rect 31576 16124 31628 16176
rect 26884 16056 26936 16108
rect 27712 16056 27764 16108
rect 30104 16056 30156 16108
rect 33140 16124 33192 16176
rect 34704 16201 34713 16235
rect 34713 16201 34747 16235
rect 34747 16201 34756 16235
rect 34704 16192 34756 16201
rect 23296 15988 23348 16040
rect 24584 16031 24636 16040
rect 24584 15997 24593 16031
rect 24593 15997 24627 16031
rect 24627 15997 24636 16031
rect 24584 15988 24636 15997
rect 26976 16031 27028 16040
rect 26976 15997 26985 16031
rect 26985 15997 27019 16031
rect 27019 15997 27028 16031
rect 26976 15988 27028 15997
rect 29184 16031 29236 16040
rect 29184 15997 29193 16031
rect 29193 15997 29227 16031
rect 29227 15997 29236 16031
rect 29184 15988 29236 15997
rect 32404 16056 32456 16108
rect 32864 16099 32916 16108
rect 32864 16065 32873 16099
rect 32873 16065 32907 16099
rect 32907 16065 32916 16099
rect 32864 16056 32916 16065
rect 32128 15988 32180 16040
rect 32220 15988 32272 16040
rect 33048 16056 33100 16108
rect 33140 15988 33192 16040
rect 36544 16192 36596 16244
rect 35716 16056 35768 16108
rect 37832 16192 37884 16244
rect 38660 16192 38712 16244
rect 43076 16192 43128 16244
rect 43168 16235 43220 16244
rect 43168 16201 43185 16235
rect 43185 16201 43219 16235
rect 43219 16201 43220 16235
rect 43168 16192 43220 16201
rect 43352 16124 43404 16176
rect 37556 16056 37608 16108
rect 37740 16099 37792 16108
rect 37740 16065 37749 16099
rect 37749 16065 37783 16099
rect 37783 16065 37792 16099
rect 37740 16056 37792 16065
rect 41420 16056 41472 16108
rect 42616 16099 42668 16108
rect 42616 16065 42625 16099
rect 42625 16065 42659 16099
rect 42659 16065 42668 16099
rect 42616 16056 42668 16065
rect 42892 16099 42944 16108
rect 42892 16065 42901 16099
rect 42901 16065 42935 16099
rect 42935 16065 42944 16099
rect 42892 16056 42944 16065
rect 42984 16099 43036 16108
rect 42984 16065 42998 16099
rect 42998 16065 43032 16099
rect 43032 16065 43036 16099
rect 42984 16056 43036 16065
rect 37832 15988 37884 16040
rect 51356 16192 51408 16244
rect 52000 16192 52052 16244
rect 52460 16192 52512 16244
rect 53104 16192 53156 16244
rect 53196 16192 53248 16244
rect 60740 16192 60792 16244
rect 65984 16192 66036 16244
rect 66076 16192 66128 16244
rect 72424 16192 72476 16244
rect 43628 16099 43680 16108
rect 43628 16065 43637 16099
rect 43637 16065 43671 16099
rect 43671 16065 43680 16099
rect 43628 16056 43680 16065
rect 43904 16099 43956 16108
rect 43904 16065 43913 16099
rect 43913 16065 43947 16099
rect 43947 16065 43956 16099
rect 43904 16056 43956 16065
rect 43996 16099 44048 16108
rect 43996 16065 44010 16099
rect 44010 16065 44044 16099
rect 44044 16065 44048 16099
rect 43996 16056 44048 16065
rect 44732 16056 44784 16108
rect 45008 16099 45060 16108
rect 45008 16065 45017 16099
rect 45017 16065 45051 16099
rect 45051 16065 45060 16099
rect 45008 16056 45060 16065
rect 45928 16124 45980 16176
rect 46480 16167 46532 16176
rect 46480 16133 46489 16167
rect 46489 16133 46523 16167
rect 46523 16133 46532 16167
rect 46480 16124 46532 16133
rect 46848 16124 46900 16176
rect 47400 16124 47452 16176
rect 45376 16056 45428 16108
rect 46204 16056 46256 16108
rect 46388 16056 46440 16108
rect 47124 16056 47176 16108
rect 47768 16099 47820 16108
rect 47492 15988 47544 16040
rect 47768 16065 47777 16099
rect 47777 16065 47811 16099
rect 47811 16065 47820 16099
rect 47768 16056 47820 16065
rect 47676 15988 47728 16040
rect 50804 16124 50856 16176
rect 50896 16124 50948 16176
rect 51172 16124 51224 16176
rect 48228 16099 48280 16108
rect 48228 16065 48237 16099
rect 48237 16065 48271 16099
rect 48271 16065 48280 16099
rect 48412 16099 48464 16108
rect 48228 16056 48280 16065
rect 48412 16065 48421 16099
rect 48421 16065 48455 16099
rect 48455 16065 48464 16099
rect 48412 16056 48464 16065
rect 48044 15988 48096 16040
rect 48596 16056 48648 16108
rect 49976 16056 50028 16108
rect 50160 16056 50212 16108
rect 29092 15920 29144 15972
rect 31944 15920 31996 15972
rect 32864 15920 32916 15972
rect 33324 15920 33376 15972
rect 35348 15920 35400 15972
rect 40684 15920 40736 15972
rect 42984 15920 43036 15972
rect 25228 15852 25280 15904
rect 26976 15852 27028 15904
rect 27712 15852 27764 15904
rect 34244 15852 34296 15904
rect 36360 15852 36412 15904
rect 37464 15852 37516 15904
rect 44456 15852 44508 15904
rect 45652 15895 45704 15904
rect 45652 15861 45661 15895
rect 45661 15861 45695 15895
rect 45695 15861 45704 15895
rect 45652 15852 45704 15861
rect 46664 15852 46716 15904
rect 47216 15920 47268 15972
rect 48136 15920 48188 15972
rect 49608 15988 49660 16040
rect 49700 15988 49752 16040
rect 49884 15988 49936 16040
rect 50344 16099 50396 16108
rect 50344 16065 50353 16099
rect 50353 16065 50387 16099
rect 50387 16065 50396 16099
rect 50344 16056 50396 16065
rect 50620 16056 50672 16108
rect 51540 16056 51592 16108
rect 51908 16056 51960 16108
rect 52460 16056 52512 16108
rect 50528 15988 50580 16040
rect 52644 15988 52696 16040
rect 52828 16056 52880 16108
rect 53748 16124 53800 16176
rect 54944 16124 54996 16176
rect 58440 16124 58492 16176
rect 58624 16124 58676 16176
rect 53196 16099 53248 16108
rect 53196 16065 53199 16099
rect 53199 16065 53248 16099
rect 53196 16056 53248 16065
rect 53932 16056 53984 16108
rect 54576 16056 54628 16108
rect 55220 16056 55272 16108
rect 56784 16056 56836 16108
rect 47768 15852 47820 15904
rect 50160 15920 50212 15972
rect 49884 15895 49936 15904
rect 49884 15861 49893 15895
rect 49893 15861 49927 15895
rect 49927 15861 49936 15895
rect 49884 15852 49936 15861
rect 50712 15852 50764 15904
rect 54208 15988 54260 16040
rect 56324 15988 56376 16040
rect 57888 16056 57940 16108
rect 58256 16099 58308 16108
rect 58256 16065 58265 16099
rect 58265 16065 58299 16099
rect 58299 16065 58308 16099
rect 58256 16056 58308 16065
rect 58348 16099 58400 16108
rect 58348 16065 58357 16099
rect 58357 16065 58391 16099
rect 58391 16065 58400 16099
rect 58348 16056 58400 16065
rect 58532 16056 58584 16108
rect 58992 16099 59044 16108
rect 58992 16065 59001 16099
rect 59001 16065 59035 16099
rect 59035 16065 59044 16099
rect 58992 16056 59044 16065
rect 59176 16099 59228 16108
rect 59176 16065 59179 16099
rect 59179 16065 59228 16099
rect 59176 16056 59228 16065
rect 57980 15988 58032 16040
rect 60004 16056 60056 16108
rect 60464 16056 60516 16108
rect 55036 15920 55088 15972
rect 60280 15988 60332 16040
rect 60372 15988 60424 16040
rect 62120 16099 62172 16108
rect 62120 16065 62129 16099
rect 62129 16065 62163 16099
rect 62163 16065 62172 16099
rect 62120 16056 62172 16065
rect 62396 16056 62448 16108
rect 62764 16056 62816 16108
rect 62212 15988 62264 16040
rect 63040 16099 63092 16108
rect 63040 16065 63049 16099
rect 63049 16065 63083 16099
rect 63083 16065 63092 16099
rect 63040 16056 63092 16065
rect 63224 16099 63276 16108
rect 63224 16065 63233 16099
rect 63233 16065 63267 16099
rect 63267 16065 63276 16099
rect 63224 16056 63276 16065
rect 64604 16056 64656 16108
rect 64880 16099 64932 16108
rect 64880 16065 64889 16099
rect 64889 16065 64923 16099
rect 64923 16065 64932 16099
rect 64880 16056 64932 16065
rect 65708 16056 65760 16108
rect 69756 16124 69808 16176
rect 73068 16124 73120 16176
rect 66444 15988 66496 16040
rect 68100 15988 68152 16040
rect 69940 16056 69992 16108
rect 71872 16056 71924 16108
rect 68928 15988 68980 16040
rect 71504 15988 71556 16040
rect 86592 15988 86644 16040
rect 58164 15920 58216 15972
rect 53840 15852 53892 15904
rect 56600 15852 56652 15904
rect 58716 15852 58768 15904
rect 58992 15852 59044 15904
rect 63776 15895 63828 15904
rect 63776 15861 63785 15895
rect 63785 15861 63819 15895
rect 63819 15861 63828 15895
rect 63776 15852 63828 15861
rect 64972 15852 65024 15904
rect 65616 15852 65668 15904
rect 69480 15920 69532 15972
rect 68744 15852 68796 15904
rect 72056 15852 72108 15904
rect 88064 15895 88116 15904
rect 88064 15861 88073 15895
rect 88073 15861 88107 15895
rect 88107 15861 88116 15895
rect 88064 15852 88116 15861
rect 11924 15750 11976 15802
rect 11988 15750 12040 15802
rect 12052 15750 12104 15802
rect 12116 15750 12168 15802
rect 12180 15750 12232 15802
rect 33872 15750 33924 15802
rect 33936 15750 33988 15802
rect 34000 15750 34052 15802
rect 34064 15750 34116 15802
rect 34128 15750 34180 15802
rect 55820 15750 55872 15802
rect 55884 15750 55936 15802
rect 55948 15750 56000 15802
rect 56012 15750 56064 15802
rect 56076 15750 56128 15802
rect 77768 15750 77820 15802
rect 77832 15750 77884 15802
rect 77896 15750 77948 15802
rect 77960 15750 78012 15802
rect 78024 15750 78076 15802
rect 22192 15648 22244 15700
rect 25596 15648 25648 15700
rect 25964 15648 26016 15700
rect 27804 15648 27856 15700
rect 32220 15648 32272 15700
rect 32496 15648 32548 15700
rect 27620 15580 27672 15632
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 20904 15512 20956 15564
rect 21916 15512 21968 15564
rect 21088 15444 21140 15496
rect 22652 15444 22704 15496
rect 25412 15512 25464 15564
rect 27896 15555 27948 15564
rect 27896 15521 27905 15555
rect 27905 15521 27939 15555
rect 27939 15521 27948 15555
rect 27896 15512 27948 15521
rect 30564 15580 30616 15632
rect 29000 15512 29052 15564
rect 33048 15648 33100 15700
rect 34428 15648 34480 15700
rect 35440 15580 35492 15632
rect 43996 15648 44048 15700
rect 45008 15648 45060 15700
rect 45376 15691 45428 15700
rect 45376 15657 45385 15691
rect 45385 15657 45419 15691
rect 45419 15657 45428 15691
rect 45376 15648 45428 15657
rect 46664 15648 46716 15700
rect 46756 15648 46808 15700
rect 48228 15648 48280 15700
rect 50252 15648 50304 15700
rect 51448 15648 51500 15700
rect 52368 15648 52420 15700
rect 53380 15648 53432 15700
rect 57244 15648 57296 15700
rect 58256 15648 58308 15700
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 26148 15444 26200 15496
rect 26976 15444 27028 15496
rect 28264 15444 28316 15496
rect 29552 15444 29604 15496
rect 31116 15444 31168 15496
rect 32036 15444 32088 15496
rect 32496 15444 32548 15496
rect 35072 15487 35124 15496
rect 35072 15453 35081 15487
rect 35081 15453 35115 15487
rect 35115 15453 35124 15487
rect 35072 15444 35124 15453
rect 35900 15512 35952 15564
rect 35348 15487 35400 15496
rect 35348 15453 35357 15487
rect 35357 15453 35391 15487
rect 35391 15453 35400 15487
rect 37372 15512 37424 15564
rect 38384 15555 38436 15564
rect 38384 15521 38393 15555
rect 38393 15521 38427 15555
rect 38427 15521 38436 15555
rect 38384 15512 38436 15521
rect 35348 15444 35400 15453
rect 37280 15444 37332 15496
rect 37648 15444 37700 15496
rect 42340 15487 42392 15496
rect 42340 15453 42349 15487
rect 42349 15453 42383 15487
rect 42383 15453 42392 15487
rect 42340 15444 42392 15453
rect 20720 15419 20772 15428
rect 20720 15385 20729 15419
rect 20729 15385 20763 15419
rect 20763 15385 20772 15419
rect 20720 15376 20772 15385
rect 22192 15376 22244 15428
rect 23940 15376 23992 15428
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 12348 15308 12400 15360
rect 22560 15308 22612 15360
rect 25136 15308 25188 15360
rect 25688 15376 25740 15428
rect 29184 15376 29236 15428
rect 30196 15419 30248 15428
rect 30196 15385 30205 15419
rect 30205 15385 30239 15419
rect 30239 15385 30248 15419
rect 30196 15376 30248 15385
rect 30656 15376 30708 15428
rect 36360 15419 36412 15428
rect 36360 15385 36394 15419
rect 36394 15385 36412 15419
rect 36360 15376 36412 15385
rect 26056 15308 26108 15360
rect 27344 15308 27396 15360
rect 28080 15308 28132 15360
rect 32496 15308 32548 15360
rect 35348 15308 35400 15360
rect 35624 15308 35676 15360
rect 37832 15376 37884 15428
rect 38568 15376 38620 15428
rect 41696 15376 41748 15428
rect 37556 15308 37608 15360
rect 41512 15308 41564 15360
rect 42432 15308 42484 15360
rect 45744 15555 45796 15564
rect 45744 15521 45753 15555
rect 45753 15521 45787 15555
rect 45787 15521 45796 15555
rect 45744 15512 45796 15521
rect 42708 15487 42760 15496
rect 42708 15453 42717 15487
rect 42717 15453 42751 15487
rect 42751 15453 42760 15487
rect 42708 15444 42760 15453
rect 45100 15487 45152 15496
rect 45100 15453 45109 15487
rect 45109 15453 45143 15487
rect 45143 15453 45152 15487
rect 45100 15444 45152 15453
rect 45376 15444 45428 15496
rect 45652 15444 45704 15496
rect 44088 15376 44140 15428
rect 47492 15512 47544 15564
rect 47676 15487 47728 15496
rect 47676 15453 47685 15487
rect 47685 15453 47719 15487
rect 47719 15453 47728 15487
rect 47676 15444 47728 15453
rect 49332 15580 49384 15632
rect 49424 15623 49476 15632
rect 49424 15589 49433 15623
rect 49433 15589 49467 15623
rect 49467 15589 49476 15623
rect 49424 15580 49476 15589
rect 53104 15580 53156 15632
rect 54116 15580 54168 15632
rect 55404 15580 55456 15632
rect 58348 15580 58400 15632
rect 53748 15555 53800 15564
rect 53748 15521 53757 15555
rect 53757 15521 53791 15555
rect 53791 15521 53800 15555
rect 53748 15512 53800 15521
rect 44272 15308 44324 15360
rect 44364 15308 44416 15360
rect 45100 15308 45152 15360
rect 45836 15308 45888 15360
rect 45928 15308 45980 15360
rect 48274 15376 48326 15428
rect 48688 15444 48740 15496
rect 50252 15444 50304 15496
rect 51080 15444 51132 15496
rect 51264 15487 51316 15496
rect 51264 15453 51273 15487
rect 51273 15453 51307 15487
rect 51307 15453 51316 15487
rect 51264 15444 51316 15453
rect 51448 15444 51500 15496
rect 51908 15487 51960 15496
rect 51908 15453 51917 15487
rect 51917 15453 51951 15487
rect 51951 15453 51960 15487
rect 51908 15444 51960 15453
rect 52276 15487 52328 15496
rect 52276 15453 52285 15487
rect 52285 15453 52319 15487
rect 52319 15453 52328 15487
rect 52276 15444 52328 15453
rect 52552 15487 52604 15496
rect 52552 15453 52561 15487
rect 52561 15453 52595 15487
rect 52595 15453 52604 15487
rect 52552 15444 52604 15453
rect 53288 15444 53340 15496
rect 58164 15512 58216 15564
rect 58256 15555 58308 15564
rect 58256 15521 58265 15555
rect 58265 15521 58299 15555
rect 58299 15521 58308 15555
rect 58256 15512 58308 15521
rect 55680 15444 55732 15496
rect 56232 15487 56284 15496
rect 56232 15453 56241 15487
rect 56241 15453 56275 15487
rect 56275 15453 56284 15487
rect 56232 15444 56284 15453
rect 56508 15444 56560 15496
rect 57520 15444 57572 15496
rect 58992 15648 59044 15700
rect 60004 15691 60056 15700
rect 60004 15657 60013 15691
rect 60013 15657 60047 15691
rect 60047 15657 60056 15691
rect 60004 15648 60056 15657
rect 60280 15648 60332 15700
rect 60832 15648 60884 15700
rect 65616 15691 65668 15700
rect 58624 15555 58676 15564
rect 58624 15521 58633 15555
rect 58633 15521 58667 15555
rect 58667 15521 58676 15555
rect 58624 15512 58676 15521
rect 60280 15512 60332 15564
rect 62396 15580 62448 15632
rect 62856 15580 62908 15632
rect 65616 15657 65625 15691
rect 65625 15657 65659 15691
rect 65659 15657 65668 15691
rect 65616 15648 65668 15657
rect 62580 15512 62632 15564
rect 62672 15512 62724 15564
rect 64144 15512 64196 15564
rect 65340 15512 65392 15564
rect 58716 15444 58768 15496
rect 60372 15444 60424 15496
rect 63040 15444 63092 15496
rect 63776 15444 63828 15496
rect 64880 15487 64932 15496
rect 64880 15453 64889 15487
rect 64889 15453 64923 15487
rect 64923 15453 64932 15487
rect 64880 15444 64932 15453
rect 65248 15444 65300 15496
rect 65800 15487 65852 15496
rect 65800 15453 65809 15487
rect 65809 15453 65843 15487
rect 65843 15453 65852 15487
rect 65800 15444 65852 15453
rect 67272 15512 67324 15564
rect 71872 15691 71924 15700
rect 71872 15657 71881 15691
rect 71881 15657 71915 15691
rect 71915 15657 71924 15691
rect 71872 15648 71924 15657
rect 69940 15580 69992 15632
rect 71228 15555 71280 15564
rect 71228 15521 71237 15555
rect 71237 15521 71271 15555
rect 71271 15521 71280 15555
rect 71228 15512 71280 15521
rect 71504 15512 71556 15564
rect 68928 15487 68980 15496
rect 50160 15419 50212 15428
rect 50160 15385 50169 15419
rect 50169 15385 50203 15419
rect 50203 15385 50212 15419
rect 50160 15376 50212 15385
rect 50804 15376 50856 15428
rect 48044 15308 48096 15360
rect 49700 15308 49752 15360
rect 49976 15308 50028 15360
rect 50436 15308 50488 15360
rect 52000 15376 52052 15428
rect 53564 15376 53616 15428
rect 53748 15376 53800 15428
rect 55128 15376 55180 15428
rect 54760 15308 54812 15360
rect 56784 15376 56836 15428
rect 57980 15376 58032 15428
rect 61844 15419 61896 15428
rect 61844 15385 61853 15419
rect 61853 15385 61887 15419
rect 61887 15385 61896 15419
rect 61844 15376 61896 15385
rect 55404 15308 55456 15360
rect 57336 15351 57388 15360
rect 57336 15317 57345 15351
rect 57345 15317 57379 15351
rect 57379 15317 57388 15351
rect 57336 15308 57388 15317
rect 57428 15308 57480 15360
rect 60556 15308 60608 15360
rect 60924 15308 60976 15360
rect 62396 15376 62448 15428
rect 62120 15308 62172 15360
rect 62672 15308 62724 15360
rect 64144 15308 64196 15360
rect 64328 15351 64380 15360
rect 64328 15317 64337 15351
rect 64337 15317 64371 15351
rect 64371 15317 64380 15351
rect 64328 15308 64380 15317
rect 64604 15308 64656 15360
rect 67824 15351 67876 15360
rect 67824 15317 67833 15351
rect 67833 15317 67867 15351
rect 67867 15317 67876 15351
rect 67824 15308 67876 15317
rect 68928 15453 68937 15487
rect 68937 15453 68971 15487
rect 68971 15453 68980 15487
rect 68928 15444 68980 15453
rect 70124 15444 70176 15496
rect 72056 15487 72108 15496
rect 72056 15453 72065 15487
rect 72065 15453 72099 15487
rect 72099 15453 72108 15487
rect 72056 15444 72108 15453
rect 72424 15487 72476 15496
rect 72424 15453 72433 15487
rect 72433 15453 72467 15487
rect 72467 15453 72476 15487
rect 72424 15444 72476 15453
rect 88064 15419 88116 15428
rect 88064 15385 88073 15419
rect 88073 15385 88107 15419
rect 88107 15385 88116 15419
rect 88064 15376 88116 15385
rect 70308 15351 70360 15360
rect 70308 15317 70317 15351
rect 70317 15317 70351 15351
rect 70351 15317 70360 15351
rect 70308 15308 70360 15317
rect 70400 15308 70452 15360
rect 88156 15351 88208 15360
rect 88156 15317 88165 15351
rect 88165 15317 88199 15351
rect 88199 15317 88208 15351
rect 88156 15308 88208 15317
rect 22898 15206 22950 15258
rect 22962 15206 23014 15258
rect 23026 15206 23078 15258
rect 23090 15206 23142 15258
rect 23154 15206 23206 15258
rect 44846 15206 44898 15258
rect 44910 15206 44962 15258
rect 44974 15206 45026 15258
rect 45038 15206 45090 15258
rect 45102 15206 45154 15258
rect 66794 15206 66846 15258
rect 66858 15206 66910 15258
rect 66922 15206 66974 15258
rect 66986 15206 67038 15258
rect 67050 15206 67102 15258
rect 11704 15104 11756 15156
rect 16488 15104 16540 15156
rect 19892 15104 19944 15156
rect 20720 15104 20772 15156
rect 12716 15036 12768 15088
rect 20904 15104 20956 15156
rect 22100 15104 22152 15156
rect 22468 15104 22520 15156
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 19064 15011 19116 15020
rect 19064 14977 19073 15011
rect 19073 14977 19107 15011
rect 19107 14977 19116 15011
rect 19064 14968 19116 14977
rect 22008 14968 22060 15020
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 23388 15036 23440 15088
rect 24308 15104 24360 15156
rect 24860 15104 24912 15156
rect 25504 15104 25556 15156
rect 25596 15104 25648 15156
rect 24676 15036 24728 15088
rect 27344 15104 27396 15156
rect 27528 15104 27580 15156
rect 31944 15104 31996 15156
rect 32128 15147 32180 15156
rect 32128 15113 32137 15147
rect 32137 15113 32171 15147
rect 32171 15113 32180 15147
rect 32128 15104 32180 15113
rect 32312 15104 32364 15156
rect 33232 15147 33284 15156
rect 33232 15113 33241 15147
rect 33241 15113 33275 15147
rect 33275 15113 33284 15147
rect 33232 15104 33284 15113
rect 33324 15104 33376 15156
rect 22744 15011 22796 15020
rect 22376 14968 22428 14977
rect 22744 14977 22753 15011
rect 22753 14977 22787 15011
rect 22787 14977 22796 15011
rect 22744 14968 22796 14977
rect 23296 14968 23348 15020
rect 20628 14900 20680 14952
rect 24216 14968 24268 15020
rect 24308 15011 24360 15020
rect 24308 14977 24317 15011
rect 24317 14977 24351 15011
rect 24351 14977 24360 15011
rect 24308 14968 24360 14977
rect 25044 15011 25096 15020
rect 24124 14900 24176 14952
rect 24400 14900 24452 14952
rect 25044 14977 25053 15011
rect 25053 14977 25087 15011
rect 25087 14977 25096 15011
rect 25044 14968 25096 14977
rect 25136 14968 25188 15020
rect 26516 14968 26568 15020
rect 27252 14968 27304 15020
rect 26240 14900 26292 14952
rect 26792 14900 26844 14952
rect 27712 14968 27764 15020
rect 27436 14900 27488 14952
rect 27528 14943 27580 14952
rect 27528 14909 27537 14943
rect 27537 14909 27571 14943
rect 27571 14909 27580 14943
rect 28908 15036 28960 15088
rect 32496 15079 32548 15088
rect 28540 15011 28592 15020
rect 28540 14977 28549 15011
rect 28549 14977 28583 15011
rect 28583 14977 28592 15011
rect 28540 14968 28592 14977
rect 29000 14968 29052 15020
rect 29184 15011 29236 15020
rect 29184 14977 29193 15011
rect 29193 14977 29227 15011
rect 29227 14977 29236 15011
rect 29184 14968 29236 14977
rect 30104 14968 30156 15020
rect 27528 14900 27580 14909
rect 28908 14900 28960 14952
rect 31300 15011 31352 15020
rect 31300 14977 31309 15011
rect 31309 14977 31343 15011
rect 31343 14977 31352 15011
rect 31300 14968 31352 14977
rect 32496 15045 32505 15079
rect 32505 15045 32539 15079
rect 32539 15045 32548 15079
rect 32496 15036 32548 15045
rect 32680 15036 32732 15088
rect 32588 14968 32640 15020
rect 33508 14968 33560 15020
rect 33600 14968 33652 15020
rect 33968 14968 34020 15020
rect 34244 15036 34296 15088
rect 35256 15011 35308 15020
rect 35256 14977 35265 15011
rect 35265 14977 35299 15011
rect 35299 14977 35308 15011
rect 35256 14968 35308 14977
rect 35440 15011 35492 15020
rect 35440 14977 35449 15011
rect 35449 14977 35483 15011
rect 35483 14977 35492 15011
rect 35440 14968 35492 14977
rect 41512 15104 41564 15156
rect 42432 15104 42484 15156
rect 53104 15104 53156 15156
rect 34520 14900 34572 14952
rect 36176 15011 36228 15020
rect 36176 14977 36185 15011
rect 36185 14977 36219 15011
rect 36219 14977 36228 15011
rect 36176 14968 36228 14977
rect 36268 14900 36320 14952
rect 36452 15011 36504 15020
rect 36452 14977 36461 15011
rect 36461 14977 36495 15011
rect 36495 14977 36504 15011
rect 36452 14968 36504 14977
rect 37096 14968 37148 15020
rect 37832 14968 37884 15020
rect 39948 14968 40000 15020
rect 41696 15011 41748 15020
rect 41696 14977 41705 15011
rect 41705 14977 41739 15011
rect 41739 14977 41748 15011
rect 41696 14968 41748 14977
rect 37280 14943 37332 14952
rect 37280 14909 37289 14943
rect 37289 14909 37323 14943
rect 37323 14909 37332 14943
rect 37280 14900 37332 14909
rect 39396 14943 39448 14952
rect 39396 14909 39405 14943
rect 39405 14909 39439 14943
rect 39439 14909 39448 14943
rect 39396 14900 39448 14909
rect 21180 14807 21232 14816
rect 21180 14773 21189 14807
rect 21189 14773 21223 14807
rect 21223 14773 21232 14807
rect 21180 14764 21232 14773
rect 21364 14807 21416 14816
rect 21364 14773 21373 14807
rect 21373 14773 21407 14807
rect 21407 14773 21416 14807
rect 21364 14764 21416 14773
rect 22100 14764 22152 14816
rect 23112 14764 23164 14816
rect 23848 14764 23900 14816
rect 24308 14807 24360 14816
rect 24308 14773 24317 14807
rect 24317 14773 24351 14807
rect 24351 14773 24360 14807
rect 24308 14764 24360 14773
rect 26424 14807 26476 14816
rect 26424 14773 26433 14807
rect 26433 14773 26467 14807
rect 26467 14773 26476 14807
rect 26424 14764 26476 14773
rect 26516 14764 26568 14816
rect 27068 14764 27120 14816
rect 27528 14764 27580 14816
rect 27988 14764 28040 14816
rect 28540 14764 28592 14816
rect 30840 14764 30892 14816
rect 31760 14764 31812 14816
rect 31852 14764 31904 14816
rect 32128 14764 32180 14816
rect 33232 14764 33284 14816
rect 34520 14764 34572 14816
rect 34704 14807 34756 14816
rect 34704 14773 34713 14807
rect 34713 14773 34747 14807
rect 34747 14773 34756 14807
rect 34704 14764 34756 14773
rect 35900 14764 35952 14816
rect 38568 14764 38620 14816
rect 40776 14807 40828 14816
rect 40776 14773 40785 14807
rect 40785 14773 40819 14807
rect 40819 14773 40828 14807
rect 40776 14764 40828 14773
rect 41788 14832 41840 14884
rect 41972 14832 42024 14884
rect 42892 14764 42944 14816
rect 43076 14943 43128 14952
rect 43076 14909 43085 14943
rect 43085 14909 43119 14943
rect 43119 14909 43128 14943
rect 43076 14900 43128 14909
rect 44364 15011 44416 15020
rect 44364 14977 44373 15011
rect 44373 14977 44407 15011
rect 44407 14977 44416 15011
rect 44364 14968 44416 14977
rect 44548 15011 44600 15020
rect 44548 14977 44557 15011
rect 44557 14977 44591 15011
rect 44591 14977 44600 15011
rect 44548 14968 44600 14977
rect 48320 14968 48372 15020
rect 48596 14968 48648 15020
rect 50436 15036 50488 15088
rect 51080 15036 51132 15088
rect 51540 15036 51592 15088
rect 43444 14900 43496 14952
rect 44088 14900 44140 14952
rect 45652 14943 45704 14952
rect 45652 14909 45661 14943
rect 45661 14909 45695 14943
rect 45695 14909 45704 14943
rect 45652 14900 45704 14909
rect 45836 14900 45888 14952
rect 46848 14900 46900 14952
rect 48872 14943 48924 14952
rect 48872 14909 48881 14943
rect 48881 14909 48915 14943
rect 48915 14909 48924 14943
rect 48872 14900 48924 14909
rect 44088 14764 44140 14816
rect 45744 14832 45796 14884
rect 46756 14832 46808 14884
rect 46940 14832 46992 14884
rect 45560 14764 45612 14816
rect 48596 14764 48648 14816
rect 49792 14764 49844 14816
rect 52920 15036 52972 15088
rect 54300 15104 54352 15156
rect 62948 15104 63000 15156
rect 64328 15104 64380 15156
rect 53840 15036 53892 15088
rect 54944 15036 54996 15088
rect 55128 15036 55180 15088
rect 53288 15011 53340 15020
rect 53288 14977 53297 15011
rect 53297 14977 53331 15011
rect 53331 14977 53340 15011
rect 53288 14968 53340 14977
rect 53472 14968 53524 15020
rect 54208 14968 54260 15020
rect 54484 15011 54536 15020
rect 54484 14977 54493 15011
rect 54493 14977 54527 15011
rect 54527 14977 54536 15011
rect 56324 15036 56376 15088
rect 58164 15036 58216 15088
rect 58256 15036 58308 15088
rect 54484 14968 54536 14977
rect 55680 14968 55732 15020
rect 56692 14968 56744 15020
rect 56876 15011 56928 15020
rect 56876 14977 56885 15011
rect 56885 14977 56919 15011
rect 56919 14977 56928 15011
rect 56876 14968 56928 14977
rect 59360 15036 59412 15088
rect 59544 14968 59596 15020
rect 61752 14968 61804 15020
rect 62028 15011 62080 15020
rect 62028 14977 62037 15011
rect 62037 14977 62071 15011
rect 62071 14977 62080 15011
rect 62028 14968 62080 14977
rect 50988 14832 51040 14884
rect 52644 14832 52696 14884
rect 55036 14875 55088 14884
rect 55036 14841 55045 14875
rect 55045 14841 55079 14875
rect 55079 14841 55088 14875
rect 55036 14832 55088 14841
rect 51080 14764 51132 14816
rect 51356 14764 51408 14816
rect 54300 14764 54352 14816
rect 54668 14807 54720 14816
rect 54668 14773 54677 14807
rect 54677 14773 54711 14807
rect 54711 14773 54720 14807
rect 54668 14764 54720 14773
rect 54852 14764 54904 14816
rect 56968 14900 57020 14952
rect 58072 14943 58124 14952
rect 58072 14909 58081 14943
rect 58081 14909 58115 14943
rect 58115 14909 58124 14943
rect 58072 14900 58124 14909
rect 58716 14900 58768 14952
rect 59360 14900 59412 14952
rect 60832 14900 60884 14952
rect 61844 14900 61896 14952
rect 65524 15104 65576 15156
rect 67272 15147 67324 15156
rect 67272 15113 67281 15147
rect 67281 15113 67315 15147
rect 67315 15113 67324 15147
rect 67272 15104 67324 15113
rect 62304 15011 62356 15020
rect 62304 14977 62313 15011
rect 62313 14977 62347 15011
rect 62347 14977 62356 15011
rect 62304 14968 62356 14977
rect 62396 15011 62448 15020
rect 62396 14977 62405 15011
rect 62405 14977 62439 15011
rect 62439 14977 62448 15011
rect 63592 15011 63644 15020
rect 62396 14968 62448 14977
rect 63592 14977 63601 15011
rect 63601 14977 63635 15011
rect 63635 14977 63644 15011
rect 63592 14968 63644 14977
rect 65248 15036 65300 15088
rect 68008 15036 68060 15088
rect 64604 15011 64656 15020
rect 64604 14977 64638 15011
rect 64638 14977 64656 15011
rect 62764 14900 62816 14952
rect 64604 14968 64656 14977
rect 65708 14968 65760 15020
rect 66444 14968 66496 15020
rect 65800 14900 65852 14952
rect 69204 15104 69256 15156
rect 69296 15147 69348 15156
rect 69296 15113 69305 15147
rect 69305 15113 69339 15147
rect 69339 15113 69348 15147
rect 69296 15104 69348 15113
rect 69664 15104 69716 15156
rect 70860 15104 70912 15156
rect 68744 15011 68796 15020
rect 68744 14977 68753 15011
rect 68753 14977 68787 15011
rect 68787 14977 68796 15011
rect 68744 14968 68796 14977
rect 68652 14900 68704 14952
rect 69204 14968 69256 15020
rect 71964 15036 72016 15088
rect 88248 15036 88300 15088
rect 69480 14968 69532 15020
rect 69756 14968 69808 15020
rect 88156 14968 88208 15020
rect 57980 14832 58032 14884
rect 63960 14832 64012 14884
rect 65340 14832 65392 14884
rect 68928 14832 68980 14884
rect 70676 14900 70728 14952
rect 58348 14764 58400 14816
rect 63224 14764 63276 14816
rect 63592 14764 63644 14816
rect 63868 14764 63920 14816
rect 64604 14764 64656 14816
rect 68744 14764 68796 14816
rect 69204 14764 69256 14816
rect 74816 14832 74868 14884
rect 71228 14764 71280 14816
rect 72056 14764 72108 14816
rect 11924 14662 11976 14714
rect 11988 14662 12040 14714
rect 12052 14662 12104 14714
rect 12116 14662 12168 14714
rect 12180 14662 12232 14714
rect 33872 14662 33924 14714
rect 33936 14662 33988 14714
rect 34000 14662 34052 14714
rect 34064 14662 34116 14714
rect 34128 14662 34180 14714
rect 55820 14662 55872 14714
rect 55884 14662 55936 14714
rect 55948 14662 56000 14714
rect 56012 14662 56064 14714
rect 56076 14662 56128 14714
rect 77768 14662 77820 14714
rect 77832 14662 77884 14714
rect 77896 14662 77948 14714
rect 77960 14662 78012 14714
rect 78024 14662 78076 14714
rect 21180 14560 21232 14612
rect 21640 14560 21692 14612
rect 22744 14560 22796 14612
rect 6644 14492 6696 14544
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 20352 14356 20404 14408
rect 22192 14492 22244 14544
rect 22560 14492 22612 14544
rect 23296 14560 23348 14612
rect 26056 14560 26108 14612
rect 26884 14560 26936 14612
rect 27068 14560 27120 14612
rect 28816 14560 28868 14612
rect 31300 14560 31352 14612
rect 31852 14560 31904 14612
rect 31944 14560 31996 14612
rect 37096 14603 37148 14612
rect 24768 14492 24820 14544
rect 24952 14492 25004 14544
rect 21732 14424 21784 14476
rect 26608 14492 26660 14544
rect 20904 14288 20956 14340
rect 22100 14356 22152 14408
rect 22284 14399 22336 14408
rect 22284 14365 22293 14399
rect 22293 14365 22327 14399
rect 22327 14365 22336 14399
rect 22284 14356 22336 14365
rect 22560 14331 22612 14340
rect 22560 14297 22569 14331
rect 22569 14297 22603 14331
rect 22603 14297 22612 14331
rect 24400 14399 24452 14408
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 22560 14288 22612 14297
rect 23940 14288 23992 14340
rect 18236 14220 18288 14272
rect 20260 14220 20312 14272
rect 20628 14220 20680 14272
rect 21548 14220 21600 14272
rect 22468 14220 22520 14272
rect 22744 14220 22796 14272
rect 24676 14331 24728 14340
rect 24676 14297 24685 14331
rect 24685 14297 24719 14331
rect 24719 14297 24728 14331
rect 25596 14356 25648 14408
rect 25780 14399 25832 14408
rect 25780 14365 25789 14399
rect 25789 14365 25823 14399
rect 25823 14365 25832 14399
rect 25780 14356 25832 14365
rect 26516 14356 26568 14408
rect 26700 14399 26752 14408
rect 26700 14365 26709 14399
rect 26709 14365 26743 14399
rect 26743 14365 26752 14399
rect 26700 14356 26752 14365
rect 27252 14356 27304 14408
rect 27896 14424 27948 14476
rect 31484 14492 31536 14544
rect 34520 14492 34572 14544
rect 35072 14492 35124 14544
rect 37096 14569 37105 14603
rect 37105 14569 37139 14603
rect 37139 14569 37148 14603
rect 37096 14560 37148 14569
rect 37832 14560 37884 14612
rect 45008 14560 45060 14612
rect 45192 14560 45244 14612
rect 50896 14560 50948 14612
rect 51632 14560 51684 14612
rect 53288 14560 53340 14612
rect 54392 14560 54444 14612
rect 30472 14424 30524 14476
rect 31668 14424 31720 14476
rect 32036 14467 32088 14476
rect 32036 14433 32045 14467
rect 32045 14433 32079 14467
rect 32079 14433 32088 14467
rect 32036 14424 32088 14433
rect 28908 14399 28960 14408
rect 28908 14365 28917 14399
rect 28917 14365 28951 14399
rect 28951 14365 28960 14399
rect 28908 14356 28960 14365
rect 29276 14356 29328 14408
rect 29644 14356 29696 14408
rect 30196 14356 30248 14408
rect 31116 14356 31168 14408
rect 31852 14356 31904 14408
rect 32772 14356 32824 14408
rect 35624 14424 35676 14476
rect 33876 14356 33928 14408
rect 34704 14356 34756 14408
rect 34980 14399 35032 14408
rect 34980 14365 34989 14399
rect 34989 14365 35023 14399
rect 35023 14365 35032 14399
rect 34980 14356 35032 14365
rect 24676 14288 24728 14297
rect 24860 14220 24912 14272
rect 25228 14220 25280 14272
rect 27068 14288 27120 14340
rect 27528 14288 27580 14340
rect 27712 14288 27764 14340
rect 28816 14288 28868 14340
rect 30748 14288 30800 14340
rect 31576 14288 31628 14340
rect 26056 14220 26108 14272
rect 27896 14220 27948 14272
rect 30012 14220 30064 14272
rect 31208 14220 31260 14272
rect 34244 14288 34296 14340
rect 34888 14288 34940 14340
rect 35440 14288 35492 14340
rect 34152 14220 34204 14272
rect 34428 14220 34480 14272
rect 35808 14331 35860 14340
rect 35808 14297 35817 14331
rect 35817 14297 35851 14331
rect 35851 14297 35860 14331
rect 38568 14424 38620 14476
rect 39396 14492 39448 14544
rect 37556 14356 37608 14408
rect 37924 14399 37976 14408
rect 37924 14365 37933 14399
rect 37933 14365 37967 14399
rect 37967 14365 37976 14399
rect 37924 14356 37976 14365
rect 38292 14399 38344 14408
rect 38292 14365 38301 14399
rect 38301 14365 38335 14399
rect 38335 14365 38344 14399
rect 38292 14356 38344 14365
rect 38476 14399 38528 14408
rect 38476 14365 38485 14399
rect 38485 14365 38519 14399
rect 38519 14365 38528 14399
rect 38476 14356 38528 14365
rect 39396 14399 39448 14408
rect 39396 14365 39405 14399
rect 39405 14365 39439 14399
rect 39439 14365 39448 14399
rect 39396 14356 39448 14365
rect 39764 14424 39816 14476
rect 41328 14492 41380 14544
rect 42800 14492 42852 14544
rect 44180 14535 44232 14544
rect 44180 14501 44189 14535
rect 44189 14501 44223 14535
rect 44223 14501 44232 14535
rect 44180 14492 44232 14501
rect 45284 14492 45336 14544
rect 45560 14535 45612 14544
rect 45560 14501 45569 14535
rect 45569 14501 45603 14535
rect 45603 14501 45612 14535
rect 45560 14492 45612 14501
rect 42156 14424 42208 14476
rect 43536 14424 43588 14476
rect 40592 14356 40644 14408
rect 41880 14399 41932 14408
rect 41880 14365 41889 14399
rect 41889 14365 41923 14399
rect 41923 14365 41932 14399
rect 41880 14356 41932 14365
rect 44824 14424 44876 14476
rect 43904 14399 43956 14408
rect 35808 14288 35860 14297
rect 36176 14288 36228 14340
rect 39948 14288 40000 14340
rect 40224 14288 40276 14340
rect 43904 14365 43913 14399
rect 43913 14365 43947 14399
rect 43947 14365 43956 14399
rect 43904 14356 43956 14365
rect 43996 14356 44048 14408
rect 44548 14356 44600 14408
rect 45284 14356 45336 14408
rect 43628 14288 43680 14340
rect 47768 14399 47820 14408
rect 47768 14365 47777 14399
rect 47777 14365 47811 14399
rect 47811 14365 47820 14399
rect 47768 14356 47820 14365
rect 50988 14492 51040 14544
rect 48596 14356 48648 14408
rect 49148 14399 49200 14408
rect 49148 14365 49157 14399
rect 49157 14365 49191 14399
rect 49191 14365 49200 14399
rect 49148 14356 49200 14365
rect 52000 14424 52052 14476
rect 50896 14356 50948 14408
rect 51080 14399 51132 14408
rect 51080 14365 51089 14399
rect 51089 14365 51123 14399
rect 51123 14365 51132 14399
rect 51080 14356 51132 14365
rect 52184 14424 52236 14476
rect 56416 14492 56468 14544
rect 58348 14492 58400 14544
rect 59636 14492 59688 14544
rect 61844 14492 61896 14544
rect 62028 14492 62080 14544
rect 70400 14492 70452 14544
rect 70768 14535 70820 14544
rect 70768 14501 70777 14535
rect 70777 14501 70811 14535
rect 70811 14501 70820 14535
rect 70768 14492 70820 14501
rect 73436 14492 73488 14544
rect 87236 14492 87288 14544
rect 54484 14424 54536 14476
rect 54852 14424 54904 14476
rect 54944 14424 54996 14476
rect 52920 14399 52972 14408
rect 50436 14288 50488 14340
rect 52920 14365 52929 14399
rect 52929 14365 52963 14399
rect 52963 14365 52972 14399
rect 52920 14356 52972 14365
rect 54116 14399 54168 14408
rect 54116 14365 54125 14399
rect 54125 14365 54159 14399
rect 54159 14365 54168 14399
rect 54116 14356 54168 14365
rect 54668 14356 54720 14408
rect 56508 14424 56560 14476
rect 58164 14424 58216 14476
rect 58440 14424 58492 14476
rect 58624 14467 58676 14476
rect 58624 14433 58633 14467
rect 58633 14433 58667 14467
rect 58667 14433 58676 14467
rect 58624 14424 58676 14433
rect 59912 14424 59964 14476
rect 57980 14356 58032 14408
rect 58072 14399 58124 14408
rect 58072 14365 58081 14399
rect 58081 14365 58115 14399
rect 58115 14365 58124 14399
rect 60464 14399 60516 14408
rect 58072 14356 58124 14365
rect 60464 14365 60473 14399
rect 60473 14365 60507 14399
rect 60507 14365 60516 14399
rect 60464 14356 60516 14365
rect 37004 14220 37056 14272
rect 37096 14220 37148 14272
rect 40776 14220 40828 14272
rect 42984 14220 43036 14272
rect 47492 14220 47544 14272
rect 47676 14263 47728 14272
rect 47676 14229 47685 14263
rect 47685 14229 47719 14263
rect 47719 14229 47728 14263
rect 47676 14220 47728 14229
rect 48412 14263 48464 14272
rect 48412 14229 48421 14263
rect 48421 14229 48455 14263
rect 48455 14229 48464 14263
rect 48412 14220 48464 14229
rect 48504 14220 48556 14272
rect 49056 14220 49108 14272
rect 49516 14220 49568 14272
rect 53932 14288 53984 14340
rect 55220 14288 55272 14340
rect 56600 14288 56652 14340
rect 56784 14331 56836 14340
rect 56784 14297 56793 14331
rect 56793 14297 56827 14331
rect 56827 14297 56836 14331
rect 56784 14288 56836 14297
rect 56968 14288 57020 14340
rect 57796 14288 57848 14340
rect 58164 14288 58216 14340
rect 59084 14288 59136 14340
rect 50620 14220 50672 14272
rect 55680 14220 55732 14272
rect 57244 14220 57296 14272
rect 60372 14288 60424 14340
rect 60924 14399 60976 14408
rect 60924 14365 60927 14399
rect 60927 14365 60976 14399
rect 60924 14356 60976 14365
rect 61292 14356 61344 14408
rect 62120 14424 62172 14476
rect 64604 14424 64656 14476
rect 61752 14356 61804 14408
rect 62028 14356 62080 14408
rect 62672 14399 62724 14408
rect 62672 14365 62681 14399
rect 62681 14365 62715 14399
rect 62715 14365 62724 14399
rect 62672 14356 62724 14365
rect 63776 14399 63828 14408
rect 63776 14365 63785 14399
rect 63785 14365 63819 14399
rect 63819 14365 63828 14399
rect 63960 14399 64012 14408
rect 63776 14356 63828 14365
rect 63960 14365 63969 14399
rect 63969 14365 64003 14399
rect 64003 14365 64012 14399
rect 63960 14356 64012 14365
rect 64052 14399 64104 14408
rect 64052 14365 64061 14399
rect 64061 14365 64095 14399
rect 64095 14365 64104 14399
rect 64420 14399 64472 14408
rect 64052 14356 64104 14365
rect 64420 14365 64429 14399
rect 64429 14365 64463 14399
rect 64463 14365 64472 14399
rect 64420 14356 64472 14365
rect 64972 14424 65024 14476
rect 65340 14424 65392 14476
rect 67456 14424 67508 14476
rect 68928 14467 68980 14476
rect 66536 14356 66588 14408
rect 66720 14399 66772 14408
rect 66720 14365 66754 14399
rect 66754 14365 66772 14399
rect 66720 14356 66772 14365
rect 68928 14433 68937 14467
rect 68937 14433 68971 14467
rect 68971 14433 68980 14467
rect 68928 14424 68980 14433
rect 70032 14424 70084 14476
rect 61384 14220 61436 14272
rect 63592 14263 63644 14272
rect 63592 14229 63601 14263
rect 63601 14229 63635 14263
rect 63635 14229 63644 14263
rect 63592 14220 63644 14229
rect 64144 14220 64196 14272
rect 68652 14288 68704 14340
rect 69204 14331 69256 14340
rect 69204 14297 69238 14331
rect 69238 14297 69256 14331
rect 69204 14288 69256 14297
rect 64972 14263 65024 14272
rect 64972 14229 64981 14263
rect 64981 14229 65015 14263
rect 65015 14229 65024 14263
rect 64972 14220 65024 14229
rect 68376 14220 68428 14272
rect 68468 14263 68520 14272
rect 68468 14229 68477 14263
rect 68477 14229 68511 14263
rect 68511 14229 68520 14263
rect 70308 14356 70360 14408
rect 82820 14424 82872 14476
rect 74816 14356 74868 14408
rect 84844 14356 84896 14408
rect 69480 14288 69532 14340
rect 72056 14331 72108 14340
rect 72056 14297 72065 14331
rect 72065 14297 72099 14331
rect 72099 14297 72108 14331
rect 72056 14288 72108 14297
rect 88064 14331 88116 14340
rect 88064 14297 88073 14331
rect 88073 14297 88107 14331
rect 88107 14297 88116 14331
rect 88064 14288 88116 14297
rect 68468 14220 68520 14229
rect 73712 14220 73764 14272
rect 88156 14263 88208 14272
rect 88156 14229 88165 14263
rect 88165 14229 88199 14263
rect 88199 14229 88208 14263
rect 88156 14220 88208 14229
rect 22898 14118 22950 14170
rect 22962 14118 23014 14170
rect 23026 14118 23078 14170
rect 23090 14118 23142 14170
rect 23154 14118 23206 14170
rect 44846 14118 44898 14170
rect 44910 14118 44962 14170
rect 44974 14118 45026 14170
rect 45038 14118 45090 14170
rect 45102 14118 45154 14170
rect 66794 14118 66846 14170
rect 66858 14118 66910 14170
rect 66922 14118 66974 14170
rect 66986 14118 67038 14170
rect 67050 14118 67102 14170
rect 21180 14016 21232 14068
rect 23480 14016 23532 14068
rect 23664 14016 23716 14068
rect 24308 14016 24360 14068
rect 24400 14016 24452 14068
rect 24952 14016 25004 14068
rect 26424 14016 26476 14068
rect 26516 14016 26568 14068
rect 29092 14059 29144 14068
rect 29092 14025 29101 14059
rect 29101 14025 29135 14059
rect 29135 14025 29144 14059
rect 29092 14016 29144 14025
rect 29368 14016 29420 14068
rect 29644 14016 29696 14068
rect 20444 13948 20496 14000
rect 18236 13880 18288 13932
rect 19800 13923 19852 13932
rect 19800 13889 19809 13923
rect 19809 13889 19843 13923
rect 19843 13889 19852 13923
rect 19800 13880 19852 13889
rect 21364 13948 21416 14000
rect 21548 13948 21600 14000
rect 22744 13880 22796 13932
rect 22836 13880 22888 13932
rect 23848 13923 23900 13932
rect 19616 13812 19668 13864
rect 21180 13812 21232 13864
rect 22192 13812 22244 13864
rect 22284 13812 22336 13864
rect 23848 13889 23857 13923
rect 23857 13889 23891 13923
rect 23891 13889 23900 13923
rect 23848 13880 23900 13889
rect 24676 13923 24728 13932
rect 24676 13889 24685 13923
rect 24685 13889 24719 13923
rect 24719 13889 24728 13923
rect 24676 13880 24728 13889
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 23296 13812 23348 13864
rect 20812 13787 20864 13796
rect 20812 13753 20821 13787
rect 20821 13753 20855 13787
rect 20855 13753 20864 13787
rect 20812 13744 20864 13753
rect 1400 13719 1452 13728
rect 1400 13685 1409 13719
rect 1409 13685 1443 13719
rect 1443 13685 1452 13719
rect 1400 13676 1452 13685
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 19156 13719 19208 13728
rect 19156 13685 19165 13719
rect 19165 13685 19199 13719
rect 19199 13685 19208 13719
rect 19156 13676 19208 13685
rect 19524 13676 19576 13728
rect 22100 13744 22152 13796
rect 22560 13744 22612 13796
rect 23572 13787 23624 13796
rect 23572 13753 23581 13787
rect 23581 13753 23615 13787
rect 23615 13753 23624 13787
rect 23572 13744 23624 13753
rect 24584 13812 24636 13864
rect 26240 13923 26292 13932
rect 26240 13889 26249 13923
rect 26249 13889 26283 13923
rect 26283 13889 26292 13923
rect 26240 13880 26292 13889
rect 26332 13923 26384 13932
rect 26332 13889 26341 13923
rect 26341 13889 26375 13923
rect 26375 13889 26384 13923
rect 26608 13948 26660 14000
rect 28080 13991 28132 14000
rect 28080 13957 28089 13991
rect 28089 13957 28123 13991
rect 28123 13957 28132 13991
rect 28080 13948 28132 13957
rect 29184 13948 29236 14000
rect 30840 13948 30892 14000
rect 31484 13991 31536 14000
rect 31484 13957 31493 13991
rect 31493 13957 31527 13991
rect 31527 13957 31536 13991
rect 31484 13948 31536 13957
rect 31668 13948 31720 14000
rect 32312 13948 32364 14000
rect 33416 13948 33468 14000
rect 33692 13948 33744 14000
rect 34796 14016 34848 14068
rect 35440 14016 35492 14068
rect 36176 14016 36228 14068
rect 37924 14016 37976 14068
rect 38752 14016 38804 14068
rect 39304 14059 39356 14068
rect 38844 13948 38896 14000
rect 26332 13880 26384 13889
rect 26700 13880 26752 13932
rect 26884 13880 26936 13932
rect 27252 13880 27304 13932
rect 24492 13744 24544 13796
rect 25780 13812 25832 13864
rect 27436 13855 27488 13864
rect 21272 13719 21324 13728
rect 21272 13685 21281 13719
rect 21281 13685 21315 13719
rect 21315 13685 21324 13719
rect 21272 13676 21324 13685
rect 21732 13676 21784 13728
rect 22468 13719 22520 13728
rect 22468 13685 22477 13719
rect 22477 13685 22511 13719
rect 22511 13685 22520 13719
rect 22468 13676 22520 13685
rect 22744 13719 22796 13728
rect 22744 13685 22753 13719
rect 22753 13685 22787 13719
rect 22787 13685 22796 13719
rect 22744 13676 22796 13685
rect 23664 13676 23716 13728
rect 23756 13676 23808 13728
rect 24032 13719 24084 13728
rect 24032 13685 24041 13719
rect 24041 13685 24075 13719
rect 24075 13685 24084 13719
rect 24032 13676 24084 13685
rect 26608 13744 26660 13796
rect 26884 13744 26936 13796
rect 27436 13821 27445 13855
rect 27445 13821 27479 13855
rect 27479 13821 27488 13855
rect 27436 13812 27488 13821
rect 28080 13812 28132 13864
rect 27620 13744 27672 13796
rect 25688 13676 25740 13728
rect 26424 13676 26476 13728
rect 28724 13744 28776 13796
rect 30104 13880 30156 13932
rect 31116 13880 31168 13932
rect 32496 13923 32548 13932
rect 32496 13889 32505 13923
rect 32505 13889 32539 13923
rect 32539 13889 32548 13923
rect 32496 13880 32548 13889
rect 33140 13880 33192 13932
rect 34428 13923 34480 13932
rect 29828 13744 29880 13796
rect 31116 13744 31168 13796
rect 34428 13889 34437 13923
rect 34437 13889 34471 13923
rect 34471 13889 34480 13923
rect 34428 13880 34480 13889
rect 34888 13880 34940 13932
rect 35072 13923 35124 13932
rect 35072 13889 35081 13923
rect 35081 13889 35115 13923
rect 35115 13889 35124 13923
rect 35072 13880 35124 13889
rect 35256 13923 35308 13932
rect 35256 13889 35265 13923
rect 35265 13889 35299 13923
rect 35299 13889 35308 13923
rect 35256 13880 35308 13889
rect 33324 13744 33376 13796
rect 33416 13744 33468 13796
rect 35164 13744 35216 13796
rect 35440 13923 35492 13932
rect 35440 13889 35477 13923
rect 35477 13889 35492 13923
rect 35440 13880 35492 13889
rect 35900 13880 35952 13932
rect 37556 13923 37608 13932
rect 37556 13889 37565 13923
rect 37565 13889 37599 13923
rect 37599 13889 37608 13923
rect 37556 13880 37608 13889
rect 37740 13923 37792 13932
rect 37740 13889 37743 13923
rect 37743 13889 37792 13923
rect 37740 13880 37792 13889
rect 38292 13923 38344 13932
rect 38292 13889 38301 13923
rect 38301 13889 38335 13923
rect 38335 13889 38344 13923
rect 38292 13880 38344 13889
rect 38384 13880 38436 13932
rect 39304 14025 39313 14059
rect 39313 14025 39347 14059
rect 39347 14025 39356 14059
rect 39304 14016 39356 14025
rect 39396 14016 39448 14068
rect 41420 14016 41472 14068
rect 41512 14016 41564 14068
rect 42524 13948 42576 14000
rect 42708 13948 42760 14000
rect 41328 13880 41380 13932
rect 41696 13923 41748 13932
rect 41696 13889 41705 13923
rect 41705 13889 41739 13923
rect 41739 13889 41748 13923
rect 41696 13880 41748 13889
rect 42984 13880 43036 13932
rect 45836 13948 45888 14000
rect 47768 13948 47820 14000
rect 44364 13880 44416 13932
rect 44548 13880 44600 13932
rect 39396 13855 39448 13864
rect 35808 13744 35860 13796
rect 37556 13744 37608 13796
rect 28632 13676 28684 13728
rect 30472 13676 30524 13728
rect 30748 13676 30800 13728
rect 39396 13821 39405 13855
rect 39405 13821 39439 13855
rect 39439 13821 39448 13855
rect 39396 13812 39448 13821
rect 37924 13676 37976 13728
rect 38108 13719 38160 13728
rect 38108 13685 38117 13719
rect 38117 13685 38151 13719
rect 38151 13685 38160 13719
rect 38108 13676 38160 13685
rect 38752 13676 38804 13728
rect 39764 13812 39816 13864
rect 39948 13812 40000 13864
rect 40316 13744 40368 13796
rect 41052 13812 41104 13864
rect 42064 13812 42116 13864
rect 42892 13855 42944 13864
rect 40776 13744 40828 13796
rect 42156 13744 42208 13796
rect 42892 13821 42901 13855
rect 42901 13821 42935 13855
rect 42935 13821 42944 13855
rect 42892 13812 42944 13821
rect 45192 13812 45244 13864
rect 43168 13744 43220 13796
rect 41052 13676 41104 13728
rect 41144 13676 41196 13728
rect 45100 13676 45152 13728
rect 46020 13880 46072 13932
rect 46480 13880 46532 13932
rect 48596 13948 48648 14000
rect 48780 13948 48832 14000
rect 49240 13948 49292 14000
rect 50160 13948 50212 14000
rect 50252 13948 50304 14000
rect 50804 13948 50856 14000
rect 50988 14016 51040 14068
rect 52000 14016 52052 14068
rect 52736 13948 52788 14000
rect 48044 13880 48096 13932
rect 48964 13880 49016 13932
rect 51448 13880 51500 13932
rect 51724 13923 51776 13932
rect 51724 13889 51733 13923
rect 51733 13889 51767 13923
rect 51767 13889 51776 13923
rect 54576 13948 54628 14000
rect 55588 13948 55640 14000
rect 56232 13948 56284 14000
rect 60556 14016 60608 14068
rect 61568 14016 61620 14068
rect 61752 13948 61804 14000
rect 62304 13948 62356 14000
rect 63040 13991 63092 14000
rect 63040 13957 63049 13991
rect 63049 13957 63083 13991
rect 63083 13957 63092 13991
rect 63040 13948 63092 13957
rect 63592 13948 63644 14000
rect 64512 14016 64564 14068
rect 64880 14016 64932 14068
rect 67732 14016 67784 14068
rect 68008 14016 68060 14068
rect 67456 13948 67508 14000
rect 69480 14016 69532 14068
rect 70216 14016 70268 14068
rect 71780 14016 71832 14068
rect 73896 14059 73948 14068
rect 73896 14025 73905 14059
rect 73905 14025 73939 14059
rect 73939 14025 73948 14059
rect 73896 14016 73948 14025
rect 51724 13880 51776 13889
rect 55036 13880 55088 13932
rect 45928 13855 45980 13864
rect 45928 13821 45937 13855
rect 45937 13821 45971 13855
rect 45971 13821 45980 13855
rect 45928 13812 45980 13821
rect 46756 13812 46808 13864
rect 49792 13855 49844 13864
rect 49792 13821 49801 13855
rect 49801 13821 49835 13855
rect 49835 13821 49844 13855
rect 49792 13812 49844 13821
rect 51540 13855 51592 13864
rect 51540 13821 51549 13855
rect 51549 13821 51583 13855
rect 51583 13821 51592 13855
rect 51540 13812 51592 13821
rect 52000 13812 52052 13864
rect 54116 13812 54168 13864
rect 56784 13880 56836 13932
rect 56876 13880 56928 13932
rect 57244 13923 57296 13932
rect 57244 13889 57253 13923
rect 57253 13889 57287 13923
rect 57287 13889 57296 13923
rect 57244 13880 57296 13889
rect 57888 13923 57940 13932
rect 57888 13889 57897 13923
rect 57897 13889 57931 13923
rect 57931 13889 57940 13923
rect 57888 13880 57940 13889
rect 55220 13812 55272 13864
rect 55680 13855 55732 13864
rect 55680 13821 55689 13855
rect 55689 13821 55723 13855
rect 55723 13821 55732 13855
rect 55680 13812 55732 13821
rect 56968 13812 57020 13864
rect 57336 13812 57388 13864
rect 58348 13880 58400 13932
rect 58532 13812 58584 13864
rect 59452 13880 59504 13932
rect 61844 13923 61896 13932
rect 59176 13812 59228 13864
rect 59268 13812 59320 13864
rect 60648 13812 60700 13864
rect 61016 13812 61068 13864
rect 61844 13889 61853 13923
rect 61853 13889 61887 13923
rect 61887 13889 61896 13923
rect 61844 13880 61896 13889
rect 62028 13923 62080 13932
rect 62028 13889 62042 13923
rect 62042 13889 62076 13923
rect 62076 13889 62080 13923
rect 62028 13880 62080 13889
rect 62488 13880 62540 13932
rect 63224 13923 63276 13932
rect 63224 13889 63233 13923
rect 63233 13889 63267 13923
rect 63267 13889 63276 13923
rect 63224 13880 63276 13889
rect 63500 13923 63552 13932
rect 63500 13889 63509 13923
rect 63509 13889 63543 13923
rect 63543 13889 63552 13923
rect 63500 13880 63552 13889
rect 64052 13923 64104 13932
rect 64052 13889 64061 13923
rect 64061 13889 64095 13923
rect 64095 13889 64104 13923
rect 64052 13880 64104 13889
rect 62580 13812 62632 13864
rect 63960 13812 64012 13864
rect 64604 13880 64656 13932
rect 64972 13880 65024 13932
rect 65156 13880 65208 13932
rect 67732 13927 67784 13932
rect 67732 13893 67741 13927
rect 67741 13893 67775 13927
rect 67775 13893 67784 13927
rect 68376 13923 68428 13932
rect 67732 13880 67784 13893
rect 68376 13889 68385 13923
rect 68385 13889 68419 13923
rect 68419 13889 68428 13923
rect 68376 13880 68428 13889
rect 69112 13948 69164 14000
rect 68652 13880 68704 13932
rect 68928 13880 68980 13932
rect 70124 13880 70176 13932
rect 71872 13880 71924 13932
rect 71964 13880 72016 13932
rect 72240 13923 72292 13932
rect 72240 13889 72249 13923
rect 72249 13889 72283 13923
rect 72283 13889 72292 13923
rect 72240 13880 72292 13889
rect 72332 13880 72384 13932
rect 73712 13923 73764 13932
rect 73712 13889 73721 13923
rect 73721 13889 73755 13923
rect 73755 13889 73764 13923
rect 73712 13880 73764 13889
rect 68008 13812 68060 13864
rect 69020 13812 69072 13864
rect 69388 13855 69440 13864
rect 69388 13821 69397 13855
rect 69397 13821 69431 13855
rect 69431 13821 69440 13855
rect 69388 13812 69440 13821
rect 71228 13855 71280 13864
rect 49056 13744 49108 13796
rect 49516 13744 49568 13796
rect 51356 13744 51408 13796
rect 52920 13744 52972 13796
rect 45836 13676 45888 13728
rect 47032 13719 47084 13728
rect 47032 13685 47041 13719
rect 47041 13685 47075 13719
rect 47075 13685 47084 13719
rect 47032 13676 47084 13685
rect 47952 13676 48004 13728
rect 50160 13676 50212 13728
rect 50436 13676 50488 13728
rect 54392 13676 54444 13728
rect 54668 13676 54720 13728
rect 54944 13676 54996 13728
rect 62120 13676 62172 13728
rect 62396 13676 62448 13728
rect 63868 13719 63920 13728
rect 63868 13685 63877 13719
rect 63877 13685 63911 13719
rect 63911 13685 63920 13719
rect 63868 13676 63920 13685
rect 68192 13744 68244 13796
rect 70584 13744 70636 13796
rect 71228 13821 71237 13855
rect 71237 13821 71271 13855
rect 71271 13821 71280 13855
rect 71228 13812 71280 13821
rect 71320 13744 71372 13796
rect 71044 13676 71096 13728
rect 88064 13719 88116 13728
rect 88064 13685 88073 13719
rect 88073 13685 88107 13719
rect 88107 13685 88116 13719
rect 88064 13676 88116 13685
rect 11924 13574 11976 13626
rect 11988 13574 12040 13626
rect 12052 13574 12104 13626
rect 12116 13574 12168 13626
rect 12180 13574 12232 13626
rect 33872 13574 33924 13626
rect 33936 13574 33988 13626
rect 34000 13574 34052 13626
rect 34064 13574 34116 13626
rect 34128 13574 34180 13626
rect 55820 13574 55872 13626
rect 55884 13574 55936 13626
rect 55948 13574 56000 13626
rect 56012 13574 56064 13626
rect 56076 13574 56128 13626
rect 77768 13574 77820 13626
rect 77832 13574 77884 13626
rect 77896 13574 77948 13626
rect 77960 13574 78012 13626
rect 78024 13574 78076 13626
rect 19064 13472 19116 13524
rect 19984 13472 20036 13524
rect 20812 13472 20864 13524
rect 19892 13447 19944 13456
rect 19616 13379 19668 13388
rect 19616 13345 19625 13379
rect 19625 13345 19659 13379
rect 19659 13345 19668 13379
rect 19616 13336 19668 13345
rect 19892 13413 19901 13447
rect 19901 13413 19935 13447
rect 19935 13413 19944 13447
rect 19892 13404 19944 13413
rect 20168 13404 20220 13456
rect 21824 13472 21876 13524
rect 22560 13472 22612 13524
rect 23296 13515 23348 13524
rect 23296 13481 23305 13515
rect 23305 13481 23339 13515
rect 23339 13481 23348 13515
rect 23296 13472 23348 13481
rect 24768 13472 24820 13524
rect 26056 13472 26108 13524
rect 27528 13472 27580 13524
rect 28264 13472 28316 13524
rect 29000 13472 29052 13524
rect 30288 13515 30340 13524
rect 30288 13481 30297 13515
rect 30297 13481 30331 13515
rect 30331 13481 30340 13515
rect 30288 13472 30340 13481
rect 30472 13472 30524 13524
rect 31944 13472 31996 13524
rect 34612 13472 34664 13524
rect 37188 13472 37240 13524
rect 38844 13472 38896 13524
rect 25872 13404 25924 13456
rect 27896 13447 27948 13456
rect 23664 13336 23716 13388
rect 24584 13379 24636 13388
rect 24584 13345 24593 13379
rect 24593 13345 24627 13379
rect 24627 13345 24636 13379
rect 24584 13336 24636 13345
rect 25504 13336 25556 13388
rect 25688 13379 25740 13388
rect 25688 13345 25697 13379
rect 25697 13345 25731 13379
rect 25731 13345 25740 13379
rect 25688 13336 25740 13345
rect 26424 13336 26476 13388
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 19064 13268 19116 13320
rect 19708 13311 19760 13320
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 19984 13311 20036 13320
rect 19984 13277 19993 13311
rect 19993 13277 20027 13311
rect 20027 13277 20036 13311
rect 19984 13268 20036 13277
rect 20076 13268 20128 13320
rect 20720 13268 20772 13320
rect 21088 13268 21140 13320
rect 22008 13311 22060 13320
rect 22008 13277 22017 13311
rect 22017 13277 22051 13311
rect 22051 13277 22060 13311
rect 22008 13268 22060 13277
rect 22376 13268 22428 13320
rect 22560 13268 22612 13320
rect 24124 13268 24176 13320
rect 24216 13268 24268 13320
rect 25044 13311 25096 13320
rect 25044 13277 25053 13311
rect 25053 13277 25087 13311
rect 25087 13277 25096 13311
rect 25044 13268 25096 13277
rect 25412 13268 25464 13320
rect 26516 13311 26568 13320
rect 26516 13277 26525 13311
rect 26525 13277 26559 13311
rect 26559 13277 26568 13311
rect 26516 13268 26568 13277
rect 26608 13311 26660 13320
rect 26608 13277 26618 13311
rect 26618 13277 26652 13311
rect 26652 13277 26660 13311
rect 26608 13268 26660 13277
rect 27528 13311 27580 13320
rect 20444 13200 20496 13252
rect 23572 13200 23624 13252
rect 23664 13200 23716 13252
rect 23940 13200 23992 13252
rect 20720 13132 20772 13184
rect 22468 13132 22520 13184
rect 27528 13277 27537 13311
rect 27537 13277 27571 13311
rect 27571 13277 27580 13311
rect 27528 13268 27580 13277
rect 27896 13413 27905 13447
rect 27905 13413 27939 13447
rect 27939 13413 27948 13447
rect 27896 13404 27948 13413
rect 28448 13404 28500 13456
rect 29184 13336 29236 13388
rect 30932 13336 30984 13388
rect 31300 13336 31352 13388
rect 31852 13379 31904 13388
rect 31852 13345 31861 13379
rect 31861 13345 31895 13379
rect 31895 13345 31904 13379
rect 31852 13336 31904 13345
rect 32588 13404 32640 13456
rect 32956 13404 33008 13456
rect 33048 13404 33100 13456
rect 32772 13336 32824 13388
rect 29184 13200 29236 13252
rect 29644 13243 29696 13252
rect 29644 13209 29653 13243
rect 29653 13209 29687 13243
rect 29687 13209 29696 13243
rect 29644 13200 29696 13209
rect 30104 13311 30156 13320
rect 30104 13277 30113 13311
rect 30113 13277 30147 13311
rect 30147 13277 30156 13311
rect 30840 13311 30892 13320
rect 30104 13268 30156 13277
rect 30840 13277 30849 13311
rect 30849 13277 30883 13311
rect 30883 13277 30892 13311
rect 30840 13268 30892 13277
rect 31668 13268 31720 13320
rect 32312 13268 32364 13320
rect 34612 13336 34664 13388
rect 35716 13404 35768 13456
rect 38660 13404 38712 13456
rect 36820 13336 36872 13388
rect 38752 13336 38804 13388
rect 33784 13268 33836 13320
rect 34152 13268 34204 13320
rect 34796 13268 34848 13320
rect 41788 13472 41840 13524
rect 42432 13472 42484 13524
rect 42984 13472 43036 13524
rect 43628 13515 43680 13524
rect 43628 13481 43637 13515
rect 43637 13481 43671 13515
rect 43671 13481 43680 13515
rect 43628 13472 43680 13481
rect 44364 13515 44416 13524
rect 44364 13481 44373 13515
rect 44373 13481 44407 13515
rect 44407 13481 44416 13515
rect 44364 13472 44416 13481
rect 44456 13472 44508 13524
rect 44640 13472 44692 13524
rect 45100 13472 45152 13524
rect 50436 13472 50488 13524
rect 51264 13472 51316 13524
rect 39948 13404 40000 13456
rect 40408 13336 40460 13388
rect 30380 13200 30432 13252
rect 26056 13175 26108 13184
rect 26056 13141 26065 13175
rect 26065 13141 26099 13175
rect 26099 13141 26108 13175
rect 26056 13132 26108 13141
rect 26240 13132 26292 13184
rect 27804 13132 27856 13184
rect 29828 13132 29880 13184
rect 30656 13132 30708 13184
rect 32680 13200 32732 13252
rect 33600 13200 33652 13252
rect 38936 13200 38988 13252
rect 39304 13311 39356 13320
rect 39304 13277 39313 13311
rect 39313 13277 39347 13311
rect 39347 13277 39356 13311
rect 39304 13268 39356 13277
rect 39396 13311 39448 13320
rect 39396 13277 39405 13311
rect 39405 13277 39439 13311
rect 39439 13277 39448 13311
rect 40132 13311 40184 13320
rect 39396 13268 39448 13277
rect 40132 13277 40141 13311
rect 40141 13277 40175 13311
rect 40175 13277 40184 13311
rect 40132 13268 40184 13277
rect 40776 13336 40828 13388
rect 41512 13268 41564 13320
rect 41696 13268 41748 13320
rect 41328 13200 41380 13252
rect 42248 13311 42300 13320
rect 42248 13277 42257 13311
rect 42257 13277 42291 13311
rect 42291 13277 42300 13311
rect 42248 13268 42300 13277
rect 42800 13268 42852 13320
rect 45284 13404 45336 13456
rect 47768 13404 47820 13456
rect 47860 13404 47912 13456
rect 48688 13404 48740 13456
rect 44272 13336 44324 13388
rect 45468 13379 45520 13388
rect 45468 13345 45477 13379
rect 45477 13345 45511 13379
rect 45511 13345 45520 13379
rect 45468 13336 45520 13345
rect 45744 13336 45796 13388
rect 47676 13336 47728 13388
rect 48872 13336 48924 13388
rect 49056 13379 49108 13388
rect 49056 13345 49065 13379
rect 49065 13345 49099 13379
rect 49099 13345 49108 13379
rect 49056 13336 49108 13345
rect 49792 13404 49844 13456
rect 50344 13404 50396 13456
rect 50528 13404 50580 13456
rect 51540 13472 51592 13524
rect 51724 13472 51776 13524
rect 54944 13472 54996 13524
rect 55036 13472 55088 13524
rect 58348 13472 58400 13524
rect 61660 13472 61712 13524
rect 63592 13515 63644 13524
rect 50160 13336 50212 13388
rect 45928 13268 45980 13320
rect 42708 13200 42760 13252
rect 43076 13200 43128 13252
rect 45652 13200 45704 13252
rect 47032 13268 47084 13320
rect 47952 13268 48004 13320
rect 48136 13268 48188 13320
rect 48688 13268 48740 13320
rect 49240 13311 49292 13320
rect 49240 13277 49249 13311
rect 49249 13277 49283 13311
rect 49283 13277 49292 13311
rect 49424 13311 49476 13320
rect 49240 13268 49292 13277
rect 49424 13277 49433 13311
rect 49433 13277 49467 13311
rect 49467 13277 49476 13311
rect 49424 13268 49476 13277
rect 49516 13268 49568 13320
rect 51264 13336 51316 13388
rect 54392 13404 54444 13456
rect 50436 13311 50488 13320
rect 50436 13277 50445 13311
rect 50445 13277 50479 13311
rect 50479 13277 50488 13311
rect 50436 13268 50488 13277
rect 46388 13200 46440 13252
rect 32956 13132 33008 13184
rect 34428 13132 34480 13184
rect 34612 13132 34664 13184
rect 35900 13132 35952 13184
rect 36728 13132 36780 13184
rect 36912 13132 36964 13184
rect 41144 13132 41196 13184
rect 42340 13132 42392 13184
rect 43444 13132 43496 13184
rect 48320 13200 48372 13252
rect 52092 13336 52144 13388
rect 53472 13336 53524 13388
rect 59452 13404 59504 13456
rect 60280 13404 60332 13456
rect 60740 13404 60792 13456
rect 60832 13404 60884 13456
rect 61108 13404 61160 13456
rect 63592 13481 63601 13515
rect 63601 13481 63635 13515
rect 63635 13481 63644 13515
rect 63592 13472 63644 13481
rect 64512 13472 64564 13524
rect 69388 13472 69440 13524
rect 64420 13404 64472 13456
rect 51816 13311 51868 13320
rect 47768 13132 47820 13184
rect 48688 13132 48740 13184
rect 51816 13277 51825 13311
rect 51825 13277 51859 13311
rect 51859 13277 51868 13311
rect 51816 13268 51868 13277
rect 52184 13268 52236 13320
rect 51632 13243 51684 13252
rect 51632 13209 51641 13243
rect 51641 13209 51675 13243
rect 51675 13209 51684 13243
rect 51632 13200 51684 13209
rect 52460 13200 52512 13252
rect 52828 13311 52880 13320
rect 52828 13277 52837 13311
rect 52837 13277 52871 13311
rect 52871 13277 52880 13311
rect 52828 13268 52880 13277
rect 54116 13268 54168 13320
rect 54392 13268 54444 13320
rect 52552 13132 52604 13184
rect 53932 13200 53984 13252
rect 55128 13200 55180 13252
rect 55312 13200 55364 13252
rect 54116 13132 54168 13184
rect 54392 13175 54444 13184
rect 54392 13141 54401 13175
rect 54401 13141 54435 13175
rect 54435 13141 54444 13175
rect 54392 13132 54444 13141
rect 55404 13132 55456 13184
rect 56968 13268 57020 13320
rect 56048 13200 56100 13252
rect 57888 13268 57940 13320
rect 58164 13268 58216 13320
rect 58348 13268 58400 13320
rect 59360 13268 59412 13320
rect 59820 13311 59872 13320
rect 59820 13277 59829 13311
rect 59829 13277 59863 13311
rect 59863 13277 59872 13311
rect 59820 13268 59872 13277
rect 59268 13200 59320 13252
rect 59636 13243 59688 13252
rect 59636 13209 59645 13243
rect 59645 13209 59679 13243
rect 59679 13209 59688 13243
rect 59636 13200 59688 13209
rect 56140 13132 56192 13184
rect 57520 13132 57572 13184
rect 58900 13132 58952 13184
rect 60556 13268 60608 13320
rect 60832 13311 60884 13320
rect 60832 13277 60846 13311
rect 60846 13277 60880 13311
rect 60880 13277 60884 13311
rect 60832 13268 60884 13277
rect 61016 13268 61068 13320
rect 61660 13311 61712 13320
rect 61660 13277 61669 13311
rect 61669 13277 61703 13311
rect 61703 13277 61712 13311
rect 61660 13268 61712 13277
rect 62212 13311 62264 13320
rect 62212 13277 62221 13311
rect 62221 13277 62255 13311
rect 62255 13277 62264 13311
rect 62212 13268 62264 13277
rect 66260 13404 66312 13456
rect 68928 13404 68980 13456
rect 68468 13268 68520 13320
rect 68836 13268 68888 13320
rect 70216 13311 70268 13320
rect 60648 13243 60700 13252
rect 60648 13209 60657 13243
rect 60657 13209 60691 13243
rect 60691 13209 60700 13243
rect 60648 13200 60700 13209
rect 62672 13132 62724 13184
rect 63316 13132 63368 13184
rect 64328 13132 64380 13184
rect 64604 13175 64656 13184
rect 64604 13141 64613 13175
rect 64613 13141 64647 13175
rect 64647 13141 64656 13175
rect 64604 13132 64656 13141
rect 67640 13243 67692 13252
rect 67640 13209 67649 13243
rect 67649 13209 67683 13243
rect 67683 13209 67692 13243
rect 67640 13200 67692 13209
rect 68192 13200 68244 13252
rect 68376 13200 68428 13252
rect 68100 13132 68152 13184
rect 68560 13132 68612 13184
rect 69664 13200 69716 13252
rect 70216 13277 70225 13311
rect 70225 13277 70259 13311
rect 70259 13277 70268 13311
rect 70216 13268 70268 13277
rect 72332 13472 72384 13524
rect 71872 13404 71924 13456
rect 70768 13311 70820 13320
rect 70768 13277 70777 13311
rect 70777 13277 70811 13311
rect 70811 13277 70820 13311
rect 70768 13268 70820 13277
rect 71044 13311 71096 13320
rect 71044 13277 71078 13311
rect 71078 13277 71096 13311
rect 71044 13268 71096 13277
rect 86776 13268 86828 13320
rect 72240 13200 72292 13252
rect 69388 13132 69440 13184
rect 72516 13132 72568 13184
rect 88064 13175 88116 13184
rect 88064 13141 88073 13175
rect 88073 13141 88107 13175
rect 88107 13141 88116 13175
rect 88064 13132 88116 13141
rect 22898 13030 22950 13082
rect 22962 13030 23014 13082
rect 23026 13030 23078 13082
rect 23090 13030 23142 13082
rect 23154 13030 23206 13082
rect 44846 13030 44898 13082
rect 44910 13030 44962 13082
rect 44974 13030 45026 13082
rect 45038 13030 45090 13082
rect 45102 13030 45154 13082
rect 66794 13030 66846 13082
rect 66858 13030 66910 13082
rect 66922 13030 66974 13082
rect 66986 13030 67038 13082
rect 67050 13030 67102 13082
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 3332 12724 3384 12776
rect 3976 12724 4028 12776
rect 19524 12792 19576 12844
rect 19064 12767 19116 12776
rect 19064 12733 19073 12767
rect 19073 12733 19107 12767
rect 19107 12733 19116 12767
rect 19064 12724 19116 12733
rect 22008 12860 22060 12912
rect 19892 12792 19944 12844
rect 20168 12792 20220 12844
rect 20352 12792 20404 12844
rect 20720 12792 20772 12844
rect 22744 12928 22796 12980
rect 24492 12971 24544 12980
rect 24492 12937 24501 12971
rect 24501 12937 24535 12971
rect 24535 12937 24544 12971
rect 24492 12928 24544 12937
rect 25228 12928 25280 12980
rect 25412 12971 25464 12980
rect 25412 12937 25421 12971
rect 25421 12937 25455 12971
rect 25455 12937 25464 12971
rect 25412 12928 25464 12937
rect 25504 12928 25556 12980
rect 26516 12928 26568 12980
rect 28540 12928 28592 12980
rect 24400 12835 24452 12844
rect 19708 12724 19760 12776
rect 19800 12588 19852 12640
rect 20444 12724 20496 12776
rect 20904 12656 20956 12708
rect 20812 12588 20864 12640
rect 23480 12724 23532 12776
rect 23756 12767 23808 12776
rect 23756 12733 23765 12767
rect 23765 12733 23799 12767
rect 23799 12733 23808 12767
rect 23756 12724 23808 12733
rect 24400 12801 24409 12835
rect 24409 12801 24443 12835
rect 24443 12801 24452 12835
rect 24400 12792 24452 12801
rect 24860 12792 24912 12844
rect 26148 12860 26200 12912
rect 29184 12928 29236 12980
rect 33876 12928 33928 12980
rect 26516 12835 26568 12844
rect 26516 12801 26525 12835
rect 26525 12801 26559 12835
rect 26559 12801 26568 12835
rect 26516 12792 26568 12801
rect 32496 12860 32548 12912
rect 30380 12792 30432 12844
rect 30932 12792 30984 12844
rect 31944 12792 31996 12844
rect 32036 12792 32088 12844
rect 32404 12835 32456 12844
rect 32404 12801 32413 12835
rect 32413 12801 32447 12835
rect 32447 12801 32456 12835
rect 32404 12792 32456 12801
rect 32588 12835 32640 12844
rect 32588 12801 32597 12835
rect 32597 12801 32631 12835
rect 32631 12801 32640 12835
rect 32588 12792 32640 12801
rect 32772 12792 32824 12844
rect 33140 12792 33192 12844
rect 36452 12928 36504 12980
rect 38292 12928 38344 12980
rect 38476 12928 38528 12980
rect 41512 12928 41564 12980
rect 34244 12860 34296 12912
rect 34612 12860 34664 12912
rect 35808 12903 35860 12912
rect 35808 12869 35817 12903
rect 35817 12869 35851 12903
rect 35851 12869 35860 12903
rect 35808 12860 35860 12869
rect 37004 12860 37056 12912
rect 38384 12860 38436 12912
rect 38936 12860 38988 12912
rect 39120 12860 39172 12912
rect 40040 12860 40092 12912
rect 40960 12860 41012 12912
rect 42248 12860 42300 12912
rect 34520 12835 34572 12844
rect 34520 12801 34529 12835
rect 34529 12801 34563 12835
rect 34563 12801 34572 12835
rect 34520 12792 34572 12801
rect 34888 12835 34940 12844
rect 23940 12699 23992 12708
rect 23940 12665 23949 12699
rect 23949 12665 23983 12699
rect 23983 12665 23992 12699
rect 23940 12656 23992 12665
rect 26700 12724 26752 12776
rect 24216 12656 24268 12708
rect 23388 12588 23440 12640
rect 25228 12631 25280 12640
rect 25228 12597 25237 12631
rect 25237 12597 25271 12631
rect 25271 12597 25280 12631
rect 25228 12588 25280 12597
rect 27252 12588 27304 12640
rect 27620 12656 27672 12708
rect 28172 12656 28224 12708
rect 28448 12724 28500 12776
rect 32864 12724 32916 12776
rect 28908 12699 28960 12708
rect 28908 12665 28917 12699
rect 28917 12665 28951 12699
rect 28951 12665 28960 12699
rect 28908 12656 28960 12665
rect 33600 12724 33652 12776
rect 34888 12801 34897 12835
rect 34897 12801 34931 12835
rect 34931 12801 34940 12835
rect 34888 12792 34940 12801
rect 35440 12792 35492 12844
rect 35716 12835 35768 12844
rect 35716 12801 35725 12835
rect 35725 12801 35759 12835
rect 35759 12801 35768 12835
rect 35716 12792 35768 12801
rect 36544 12835 36596 12844
rect 36544 12801 36553 12835
rect 36553 12801 36587 12835
rect 36587 12801 36596 12835
rect 36544 12792 36596 12801
rect 37648 12792 37700 12844
rect 40408 12792 40460 12844
rect 41512 12835 41564 12844
rect 41512 12801 41521 12835
rect 41521 12801 41555 12835
rect 41555 12801 41564 12835
rect 41512 12792 41564 12801
rect 42892 12860 42944 12912
rect 29092 12588 29144 12640
rect 30012 12588 30064 12640
rect 32036 12588 32088 12640
rect 32220 12631 32272 12640
rect 32220 12597 32229 12631
rect 32229 12597 32263 12631
rect 32263 12597 32272 12631
rect 32220 12588 32272 12597
rect 32956 12588 33008 12640
rect 34428 12656 34480 12708
rect 37924 12724 37976 12776
rect 38016 12724 38068 12776
rect 42432 12835 42484 12844
rect 42432 12801 42441 12835
rect 42441 12801 42475 12835
rect 42475 12801 42484 12835
rect 42432 12792 42484 12801
rect 42616 12792 42668 12844
rect 45652 12928 45704 12980
rect 46388 12971 46440 12980
rect 46388 12937 46397 12971
rect 46397 12937 46431 12971
rect 46431 12937 46440 12971
rect 46388 12928 46440 12937
rect 48320 12971 48372 12980
rect 48320 12937 48329 12971
rect 48329 12937 48363 12971
rect 48363 12937 48372 12971
rect 48320 12928 48372 12937
rect 47676 12860 47728 12912
rect 47768 12860 47820 12912
rect 43996 12835 44048 12844
rect 43996 12801 44005 12835
rect 44005 12801 44039 12835
rect 44039 12801 44048 12835
rect 43996 12792 44048 12801
rect 44732 12835 44784 12844
rect 33508 12588 33560 12640
rect 33876 12588 33928 12640
rect 41788 12656 41840 12708
rect 35072 12631 35124 12640
rect 35072 12597 35081 12631
rect 35081 12597 35115 12631
rect 35115 12597 35124 12631
rect 35072 12588 35124 12597
rect 36544 12588 36596 12640
rect 36636 12588 36688 12640
rect 39948 12588 40000 12640
rect 40224 12588 40276 12640
rect 42984 12724 43036 12776
rect 43812 12767 43864 12776
rect 43812 12733 43821 12767
rect 43821 12733 43855 12767
rect 43855 12733 43864 12767
rect 43812 12724 43864 12733
rect 43904 12767 43956 12776
rect 43904 12733 43913 12767
rect 43913 12733 43947 12767
rect 43947 12733 43956 12767
rect 43904 12724 43956 12733
rect 44088 12767 44140 12776
rect 44088 12733 44097 12767
rect 44097 12733 44131 12767
rect 44131 12733 44140 12767
rect 44732 12801 44741 12835
rect 44741 12801 44775 12835
rect 44775 12801 44784 12835
rect 44732 12792 44784 12801
rect 44824 12835 44876 12844
rect 44824 12801 44833 12835
rect 44833 12801 44867 12835
rect 44867 12801 44876 12835
rect 44824 12792 44876 12801
rect 45652 12835 45704 12844
rect 45652 12801 45661 12835
rect 45661 12801 45695 12835
rect 45695 12801 45704 12835
rect 45652 12792 45704 12801
rect 46112 12792 46164 12844
rect 46572 12835 46624 12844
rect 46572 12801 46581 12835
rect 46581 12801 46615 12835
rect 46615 12801 46624 12835
rect 46572 12792 46624 12801
rect 46756 12835 46808 12844
rect 46756 12801 46765 12835
rect 46765 12801 46799 12835
rect 46799 12801 46808 12835
rect 46756 12792 46808 12801
rect 46848 12835 46900 12844
rect 46848 12801 46883 12835
rect 46883 12801 46900 12835
rect 47032 12835 47084 12844
rect 46848 12792 46900 12801
rect 47032 12801 47041 12835
rect 47041 12801 47075 12835
rect 47075 12801 47084 12835
rect 47032 12792 47084 12801
rect 47216 12792 47268 12844
rect 50436 12928 50488 12980
rect 51448 12928 51500 12980
rect 52828 12928 52880 12980
rect 55956 12928 56008 12980
rect 50804 12860 50856 12912
rect 52092 12860 52144 12912
rect 52184 12860 52236 12912
rect 57060 12928 57112 12980
rect 57520 12928 57572 12980
rect 57612 12928 57664 12980
rect 59084 12928 59136 12980
rect 59176 12928 59228 12980
rect 59452 12928 59504 12980
rect 61016 12928 61068 12980
rect 59820 12903 59872 12912
rect 59820 12869 59829 12903
rect 59829 12869 59863 12903
rect 59863 12869 59872 12903
rect 59820 12860 59872 12869
rect 60556 12860 60608 12912
rect 62212 12928 62264 12980
rect 61844 12860 61896 12912
rect 49148 12792 49200 12844
rect 49608 12792 49660 12844
rect 50988 12792 51040 12844
rect 44088 12724 44140 12733
rect 45284 12724 45336 12776
rect 45468 12724 45520 12776
rect 45744 12767 45796 12776
rect 45744 12733 45753 12767
rect 45753 12733 45787 12767
rect 45787 12733 45796 12767
rect 45744 12724 45796 12733
rect 46020 12724 46072 12776
rect 48044 12724 48096 12776
rect 50160 12724 50212 12776
rect 50436 12724 50488 12776
rect 50804 12724 50856 12776
rect 51816 12792 51868 12844
rect 52276 12792 52328 12844
rect 52828 12792 52880 12844
rect 53104 12835 53156 12844
rect 53104 12801 53113 12835
rect 53113 12801 53147 12835
rect 53147 12801 53156 12835
rect 53104 12792 53156 12801
rect 53196 12835 53248 12844
rect 53196 12801 53205 12835
rect 53205 12801 53239 12835
rect 53239 12801 53248 12835
rect 53196 12792 53248 12801
rect 53656 12792 53708 12844
rect 52736 12724 52788 12776
rect 53288 12724 53340 12776
rect 53840 12835 53892 12844
rect 53840 12801 53849 12835
rect 53849 12801 53883 12835
rect 53883 12801 53892 12835
rect 53840 12792 53892 12801
rect 54484 12792 54536 12844
rect 55312 12792 55364 12844
rect 55680 12792 55732 12844
rect 56416 12792 56468 12844
rect 56692 12835 56744 12844
rect 56692 12801 56701 12835
rect 56701 12801 56735 12835
rect 56735 12801 56744 12835
rect 56692 12792 56744 12801
rect 56784 12792 56836 12844
rect 54576 12724 54628 12776
rect 56140 12724 56192 12776
rect 56968 12724 57020 12776
rect 42248 12588 42300 12640
rect 43720 12588 43772 12640
rect 43904 12588 43956 12640
rect 44640 12588 44692 12640
rect 45560 12588 45612 12640
rect 45928 12588 45980 12640
rect 48044 12588 48096 12640
rect 48136 12631 48188 12640
rect 48136 12597 48145 12631
rect 48145 12597 48179 12631
rect 48179 12597 48188 12631
rect 50896 12656 50948 12708
rect 51816 12656 51868 12708
rect 52368 12656 52420 12708
rect 57336 12724 57388 12776
rect 57520 12792 57572 12844
rect 57612 12792 57664 12844
rect 57980 12792 58032 12844
rect 58716 12792 58768 12844
rect 58072 12724 58124 12776
rect 60648 12792 60700 12844
rect 63500 12928 63552 12980
rect 63960 12928 64012 12980
rect 64604 12860 64656 12912
rect 65064 12928 65116 12980
rect 66352 12928 66404 12980
rect 68376 12928 68428 12980
rect 59452 12724 59504 12776
rect 62672 12792 62724 12844
rect 65156 12792 65208 12844
rect 65340 12835 65392 12844
rect 63040 12767 63092 12776
rect 63040 12733 63049 12767
rect 63049 12733 63083 12767
rect 63083 12733 63092 12767
rect 63040 12724 63092 12733
rect 64052 12724 64104 12776
rect 65340 12801 65349 12835
rect 65349 12801 65383 12835
rect 65383 12801 65392 12835
rect 65340 12792 65392 12801
rect 67916 12860 67968 12912
rect 66260 12835 66312 12844
rect 66260 12801 66269 12835
rect 66269 12801 66303 12835
rect 66303 12801 66312 12835
rect 66260 12792 66312 12801
rect 66352 12792 66404 12844
rect 66720 12792 66772 12844
rect 67456 12792 67508 12844
rect 68928 12860 68980 12912
rect 70032 12928 70084 12980
rect 86776 12971 86828 12980
rect 86776 12937 86785 12971
rect 86785 12937 86819 12971
rect 86819 12937 86828 12971
rect 86776 12928 86828 12937
rect 69112 12792 69164 12844
rect 69388 12792 69440 12844
rect 69480 12835 69532 12844
rect 69480 12801 69489 12835
rect 69489 12801 69523 12835
rect 69523 12801 69532 12835
rect 69480 12792 69532 12801
rect 69756 12792 69808 12844
rect 70308 12860 70360 12912
rect 88156 12860 88208 12912
rect 71688 12792 71740 12844
rect 71872 12792 71924 12844
rect 72332 12835 72384 12844
rect 72332 12801 72341 12835
rect 72341 12801 72375 12835
rect 72375 12801 72384 12835
rect 72332 12792 72384 12801
rect 86960 12835 87012 12844
rect 86960 12801 86969 12835
rect 86969 12801 87003 12835
rect 87003 12801 87012 12835
rect 86960 12792 87012 12801
rect 87052 12792 87104 12844
rect 60464 12656 60516 12708
rect 60648 12656 60700 12708
rect 48872 12631 48924 12640
rect 48136 12588 48188 12597
rect 48872 12597 48881 12631
rect 48881 12597 48915 12631
rect 48915 12597 48924 12631
rect 48872 12588 48924 12597
rect 50620 12588 50672 12640
rect 52552 12588 52604 12640
rect 54392 12588 54444 12640
rect 55312 12588 55364 12640
rect 55588 12588 55640 12640
rect 55956 12588 56008 12640
rect 60004 12588 60056 12640
rect 60096 12588 60148 12640
rect 61016 12588 61068 12640
rect 64512 12656 64564 12708
rect 69664 12724 69716 12776
rect 69848 12767 69900 12776
rect 69848 12733 69857 12767
rect 69857 12733 69891 12767
rect 69891 12733 69900 12767
rect 69848 12724 69900 12733
rect 66260 12588 66312 12640
rect 69756 12656 69808 12708
rect 69296 12588 69348 12640
rect 70032 12588 70084 12640
rect 71780 12588 71832 12640
rect 72424 12631 72476 12640
rect 72424 12597 72433 12631
rect 72433 12597 72467 12631
rect 72467 12597 72476 12631
rect 72424 12588 72476 12597
rect 88064 12631 88116 12640
rect 88064 12597 88073 12631
rect 88073 12597 88107 12631
rect 88107 12597 88116 12631
rect 88064 12588 88116 12597
rect 11924 12486 11976 12538
rect 11988 12486 12040 12538
rect 12052 12486 12104 12538
rect 12116 12486 12168 12538
rect 12180 12486 12232 12538
rect 33872 12486 33924 12538
rect 33936 12486 33988 12538
rect 34000 12486 34052 12538
rect 34064 12486 34116 12538
rect 34128 12486 34180 12538
rect 55820 12486 55872 12538
rect 55884 12486 55936 12538
rect 55948 12486 56000 12538
rect 56012 12486 56064 12538
rect 56076 12486 56128 12538
rect 77768 12486 77820 12538
rect 77832 12486 77884 12538
rect 77896 12486 77948 12538
rect 77960 12486 78012 12538
rect 78024 12486 78076 12538
rect 20076 12427 20128 12436
rect 20076 12393 20085 12427
rect 20085 12393 20119 12427
rect 20119 12393 20128 12427
rect 20076 12384 20128 12393
rect 20168 12384 20220 12436
rect 18972 12316 19024 12368
rect 20812 12291 20864 12300
rect 20812 12257 20821 12291
rect 20821 12257 20855 12291
rect 20855 12257 20864 12291
rect 20812 12248 20864 12257
rect 21088 12316 21140 12368
rect 21364 12384 21416 12436
rect 25136 12384 25188 12436
rect 25228 12384 25280 12436
rect 27804 12384 27856 12436
rect 28540 12384 28592 12436
rect 28816 12384 28868 12436
rect 30932 12427 30984 12436
rect 24952 12248 25004 12300
rect 26056 12291 26108 12300
rect 26056 12257 26065 12291
rect 26065 12257 26099 12291
rect 26099 12257 26108 12291
rect 26056 12248 26108 12257
rect 28264 12316 28316 12368
rect 20720 12180 20772 12232
rect 20996 12223 21048 12232
rect 20996 12189 21005 12223
rect 21005 12189 21039 12223
rect 21039 12189 21048 12223
rect 20996 12180 21048 12189
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 21548 12180 21600 12232
rect 23480 12180 23532 12232
rect 25228 12180 25280 12232
rect 26148 12223 26200 12232
rect 1676 12044 1728 12096
rect 20168 12044 20220 12096
rect 24400 12112 24452 12164
rect 26148 12189 26157 12223
rect 26157 12189 26191 12223
rect 26191 12189 26200 12223
rect 26148 12180 26200 12189
rect 26332 12223 26384 12232
rect 26332 12189 26341 12223
rect 26341 12189 26375 12223
rect 26375 12189 26384 12223
rect 26332 12180 26384 12189
rect 26792 12180 26844 12232
rect 27620 12112 27672 12164
rect 28080 12112 28132 12164
rect 20536 12044 20588 12096
rect 21548 12044 21600 12096
rect 24952 12087 25004 12096
rect 24952 12053 24961 12087
rect 24961 12053 24995 12087
rect 24995 12053 25004 12087
rect 24952 12044 25004 12053
rect 25044 12044 25096 12096
rect 27160 12087 27212 12096
rect 27160 12053 27169 12087
rect 27169 12053 27203 12087
rect 27203 12053 27212 12087
rect 27160 12044 27212 12053
rect 27252 12044 27304 12096
rect 28632 12180 28684 12232
rect 29092 12223 29144 12232
rect 29092 12189 29101 12223
rect 29101 12189 29135 12223
rect 29135 12189 29144 12223
rect 29092 12180 29144 12189
rect 30932 12393 30941 12427
rect 30941 12393 30975 12427
rect 30975 12393 30984 12427
rect 30932 12384 30984 12393
rect 31576 12427 31628 12436
rect 31576 12393 31585 12427
rect 31585 12393 31619 12427
rect 31619 12393 31628 12427
rect 31576 12384 31628 12393
rect 33048 12384 33100 12436
rect 34520 12384 34572 12436
rect 35808 12384 35860 12436
rect 35992 12427 36044 12436
rect 35992 12393 36001 12427
rect 36001 12393 36035 12427
rect 36035 12393 36044 12427
rect 35992 12384 36044 12393
rect 36176 12384 36228 12436
rect 32128 12316 32180 12368
rect 29552 12291 29604 12300
rect 29552 12257 29561 12291
rect 29561 12257 29595 12291
rect 29595 12257 29604 12291
rect 29552 12248 29604 12257
rect 32220 12248 32272 12300
rect 32864 12316 32916 12368
rect 33508 12291 33560 12300
rect 33508 12257 33517 12291
rect 33517 12257 33551 12291
rect 33551 12257 33560 12291
rect 33508 12248 33560 12257
rect 31760 12223 31812 12232
rect 31760 12189 31769 12223
rect 31769 12189 31803 12223
rect 31803 12189 31812 12223
rect 31760 12180 31812 12189
rect 33048 12180 33100 12232
rect 33324 12223 33376 12232
rect 33324 12189 33333 12223
rect 33333 12189 33367 12223
rect 33367 12189 33376 12223
rect 33324 12180 33376 12189
rect 33784 12180 33836 12232
rect 28908 12044 28960 12096
rect 32864 12112 32916 12164
rect 34336 12248 34388 12300
rect 35256 12316 35308 12368
rect 36544 12316 36596 12368
rect 38016 12316 38068 12368
rect 39396 12427 39448 12436
rect 39396 12393 39405 12427
rect 39405 12393 39439 12427
rect 39439 12393 39448 12427
rect 39396 12384 39448 12393
rect 42248 12384 42300 12436
rect 44088 12384 44140 12436
rect 44180 12384 44232 12436
rect 45744 12384 45796 12436
rect 34612 12180 34664 12232
rect 35532 12248 35584 12300
rect 35624 12248 35676 12300
rect 36084 12248 36136 12300
rect 37556 12248 37608 12300
rect 40960 12291 41012 12300
rect 36544 12223 36596 12232
rect 35256 12155 35308 12164
rect 32220 12044 32272 12096
rect 32956 12044 33008 12096
rect 35256 12121 35265 12155
rect 35265 12121 35299 12155
rect 35299 12121 35308 12155
rect 35256 12112 35308 12121
rect 36544 12189 36553 12223
rect 36553 12189 36587 12223
rect 36587 12189 36596 12223
rect 36544 12180 36596 12189
rect 36728 12223 36780 12232
rect 36728 12189 36737 12223
rect 36737 12189 36771 12223
rect 36771 12189 36780 12223
rect 36728 12180 36780 12189
rect 36820 12223 36872 12232
rect 36820 12189 36829 12223
rect 36829 12189 36863 12223
rect 36863 12189 36872 12223
rect 36820 12180 36872 12189
rect 37096 12180 37148 12232
rect 38016 12223 38068 12232
rect 38016 12189 38025 12223
rect 38025 12189 38059 12223
rect 38059 12189 38068 12223
rect 38016 12180 38068 12189
rect 38108 12180 38160 12232
rect 38568 12180 38620 12232
rect 40040 12223 40092 12232
rect 40040 12189 40049 12223
rect 40049 12189 40083 12223
rect 40083 12189 40092 12223
rect 40040 12180 40092 12189
rect 40224 12223 40276 12232
rect 40224 12189 40233 12223
rect 40233 12189 40267 12223
rect 40267 12189 40276 12223
rect 40224 12180 40276 12189
rect 40960 12257 40969 12291
rect 40969 12257 41003 12291
rect 41003 12257 41012 12291
rect 40960 12248 41012 12257
rect 43352 12248 43404 12300
rect 46020 12316 46072 12368
rect 46296 12359 46348 12368
rect 46296 12325 46305 12359
rect 46305 12325 46339 12359
rect 46339 12325 46348 12359
rect 46296 12316 46348 12325
rect 40500 12180 40552 12232
rect 42984 12223 43036 12232
rect 42984 12189 42993 12223
rect 42993 12189 43027 12223
rect 43027 12189 43036 12223
rect 42984 12180 43036 12189
rect 44364 12223 44416 12232
rect 44364 12189 44373 12223
rect 44373 12189 44407 12223
rect 44407 12189 44416 12223
rect 44364 12180 44416 12189
rect 45468 12248 45520 12300
rect 46204 12248 46256 12300
rect 48228 12384 48280 12436
rect 48044 12316 48096 12368
rect 50988 12384 51040 12436
rect 53104 12384 53156 12436
rect 53288 12384 53340 12436
rect 53932 12384 53984 12436
rect 55404 12384 55456 12436
rect 46848 12248 46900 12300
rect 47308 12248 47360 12300
rect 45560 12223 45612 12232
rect 45560 12189 45569 12223
rect 45569 12189 45603 12223
rect 45603 12189 45612 12223
rect 45560 12180 45612 12189
rect 46572 12223 46624 12232
rect 39672 12112 39724 12164
rect 40132 12112 40184 12164
rect 34980 12044 35032 12096
rect 35164 12087 35216 12096
rect 35164 12053 35173 12087
rect 35173 12053 35207 12087
rect 35207 12053 35216 12087
rect 35164 12044 35216 12053
rect 35900 12044 35952 12096
rect 36176 12044 36228 12096
rect 36268 12044 36320 12096
rect 40592 12087 40644 12096
rect 40592 12053 40601 12087
rect 40601 12053 40635 12087
rect 40635 12053 40644 12087
rect 40592 12044 40644 12053
rect 41236 12155 41288 12164
rect 41236 12121 41270 12155
rect 41270 12121 41288 12155
rect 41236 12112 41288 12121
rect 43168 12112 43220 12164
rect 46572 12189 46581 12223
rect 46581 12189 46615 12223
rect 46615 12189 46624 12223
rect 46572 12180 46624 12189
rect 47584 12180 47636 12232
rect 48320 12180 48372 12232
rect 53380 12316 53432 12368
rect 53840 12316 53892 12368
rect 57060 12384 57112 12436
rect 57152 12384 57204 12436
rect 57520 12384 57572 12436
rect 59636 12384 59688 12436
rect 59912 12384 59964 12436
rect 61844 12427 61896 12436
rect 56600 12316 56652 12368
rect 57796 12316 57848 12368
rect 57888 12316 57940 12368
rect 61844 12393 61853 12427
rect 61853 12393 61887 12427
rect 61887 12393 61896 12427
rect 61844 12384 61896 12393
rect 63500 12384 63552 12436
rect 64788 12384 64840 12436
rect 65156 12384 65208 12436
rect 65984 12384 66036 12436
rect 67548 12384 67600 12436
rect 67916 12427 67968 12436
rect 67916 12393 67925 12427
rect 67925 12393 67959 12427
rect 67959 12393 67968 12427
rect 67916 12384 67968 12393
rect 68560 12384 68612 12436
rect 69112 12384 69164 12436
rect 69296 12384 69348 12436
rect 69480 12427 69532 12436
rect 69480 12393 69489 12427
rect 69489 12393 69523 12427
rect 69523 12393 69532 12427
rect 69480 12384 69532 12393
rect 48964 12248 49016 12300
rect 50436 12291 50488 12300
rect 48596 12223 48648 12232
rect 48596 12189 48605 12223
rect 48605 12189 48639 12223
rect 48639 12189 48648 12223
rect 48596 12180 48648 12189
rect 50436 12257 50445 12291
rect 50445 12257 50479 12291
rect 50479 12257 50488 12291
rect 50436 12248 50488 12257
rect 49700 12223 49752 12232
rect 49700 12189 49709 12223
rect 49709 12189 49743 12223
rect 49743 12189 49752 12223
rect 49700 12180 49752 12189
rect 49976 12180 50028 12232
rect 50252 12180 50304 12232
rect 50344 12180 50396 12232
rect 55128 12248 55180 12300
rect 55220 12248 55272 12300
rect 46296 12112 46348 12164
rect 47768 12112 47820 12164
rect 48228 12112 48280 12164
rect 49424 12155 49476 12164
rect 49424 12121 49433 12155
rect 49433 12121 49467 12155
rect 49467 12121 49476 12155
rect 49424 12112 49476 12121
rect 53564 12180 53616 12232
rect 54300 12223 54352 12232
rect 52092 12112 52144 12164
rect 41604 12044 41656 12096
rect 43812 12044 43864 12096
rect 47676 12044 47728 12096
rect 47860 12087 47912 12096
rect 47860 12053 47869 12087
rect 47869 12053 47903 12087
rect 47903 12053 47912 12087
rect 53748 12112 53800 12164
rect 54300 12189 54309 12223
rect 54309 12189 54343 12223
rect 54343 12189 54352 12223
rect 54300 12180 54352 12189
rect 54668 12223 54720 12232
rect 54668 12189 54677 12223
rect 54677 12189 54711 12223
rect 54711 12189 54720 12223
rect 54668 12180 54720 12189
rect 55404 12180 55456 12232
rect 56784 12248 56836 12300
rect 55588 12112 55640 12164
rect 57060 12180 57112 12232
rect 57612 12180 57664 12232
rect 57796 12180 57848 12232
rect 57980 12180 58032 12232
rect 59176 12291 59228 12300
rect 59176 12257 59185 12291
rect 59185 12257 59219 12291
rect 59219 12257 59228 12291
rect 59176 12248 59228 12257
rect 60464 12291 60516 12300
rect 60464 12257 60473 12291
rect 60473 12257 60507 12291
rect 60507 12257 60516 12291
rect 60464 12248 60516 12257
rect 58348 12112 58400 12164
rect 59176 12112 59228 12164
rect 60004 12180 60056 12232
rect 68652 12316 68704 12368
rect 69388 12316 69440 12368
rect 62304 12223 62356 12232
rect 62304 12189 62313 12223
rect 62313 12189 62347 12223
rect 62347 12189 62356 12223
rect 62304 12180 62356 12189
rect 60740 12155 60792 12164
rect 60740 12121 60774 12155
rect 60774 12121 60792 12155
rect 60740 12112 60792 12121
rect 62396 12112 62448 12164
rect 62672 12180 62724 12232
rect 63224 12223 63276 12232
rect 63224 12189 63233 12223
rect 63233 12189 63267 12223
rect 63267 12189 63276 12223
rect 63224 12180 63276 12189
rect 64052 12180 64104 12232
rect 64512 12223 64564 12232
rect 64512 12189 64521 12223
rect 64521 12189 64555 12223
rect 64555 12189 64564 12223
rect 64512 12180 64564 12189
rect 64696 12180 64748 12232
rect 64420 12112 64472 12164
rect 64880 12155 64932 12164
rect 64880 12121 64889 12155
rect 64889 12121 64923 12155
rect 64923 12121 64932 12155
rect 64880 12112 64932 12121
rect 70216 12384 70268 12436
rect 82176 12384 82228 12436
rect 72332 12316 72384 12368
rect 70768 12291 70820 12300
rect 65340 12180 65392 12232
rect 66536 12223 66588 12232
rect 66536 12189 66545 12223
rect 66545 12189 66579 12223
rect 66579 12189 66588 12223
rect 66536 12180 66588 12189
rect 67180 12112 67232 12164
rect 67272 12112 67324 12164
rect 68560 12112 68612 12164
rect 70768 12257 70777 12291
rect 70777 12257 70811 12291
rect 70811 12257 70820 12291
rect 70768 12248 70820 12257
rect 68928 12223 68980 12232
rect 68928 12189 68937 12223
rect 68937 12189 68971 12223
rect 68971 12189 68980 12223
rect 68928 12180 68980 12189
rect 69388 12112 69440 12164
rect 69664 12180 69716 12232
rect 70308 12223 70360 12232
rect 70308 12189 70317 12223
rect 70317 12189 70351 12223
rect 70351 12189 70360 12223
rect 70308 12180 70360 12189
rect 71320 12180 71372 12232
rect 70032 12155 70084 12164
rect 70032 12121 70041 12155
rect 70041 12121 70075 12155
rect 70075 12121 70084 12155
rect 70032 12112 70084 12121
rect 70124 12112 70176 12164
rect 47860 12044 47912 12053
rect 52828 12044 52880 12096
rect 53656 12044 53708 12096
rect 53932 12044 53984 12096
rect 54760 12044 54812 12096
rect 54852 12044 54904 12096
rect 56600 12044 56652 12096
rect 57796 12044 57848 12096
rect 58624 12044 58676 12096
rect 60372 12044 60424 12096
rect 60648 12044 60700 12096
rect 62764 12044 62816 12096
rect 68100 12044 68152 12096
rect 68836 12087 68888 12096
rect 68836 12053 68845 12087
rect 68845 12053 68879 12087
rect 68879 12053 68888 12087
rect 68836 12044 68888 12053
rect 68928 12044 68980 12096
rect 69756 12044 69808 12096
rect 87144 12316 87196 12368
rect 22898 11942 22950 11994
rect 22962 11942 23014 11994
rect 23026 11942 23078 11994
rect 23090 11942 23142 11994
rect 23154 11942 23206 11994
rect 44846 11942 44898 11994
rect 44910 11942 44962 11994
rect 44974 11942 45026 11994
rect 45038 11942 45090 11994
rect 45102 11942 45154 11994
rect 66794 11942 66846 11994
rect 66858 11942 66910 11994
rect 66922 11942 66974 11994
rect 66986 11942 67038 11994
rect 67050 11942 67102 11994
rect 23572 11840 23624 11892
rect 23756 11840 23808 11892
rect 26056 11840 26108 11892
rect 26424 11883 26476 11892
rect 26424 11849 26433 11883
rect 26433 11849 26467 11883
rect 26467 11849 26476 11883
rect 26424 11840 26476 11849
rect 26792 11840 26844 11892
rect 28448 11840 28500 11892
rect 30012 11840 30064 11892
rect 30104 11840 30156 11892
rect 16580 11772 16632 11824
rect 20168 11772 20220 11824
rect 21364 11772 21416 11824
rect 25320 11772 25372 11824
rect 27988 11772 28040 11824
rect 29828 11772 29880 11824
rect 18788 11747 18840 11756
rect 18788 11713 18797 11747
rect 18797 11713 18831 11747
rect 18831 11713 18840 11747
rect 18788 11704 18840 11713
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 19708 11704 19760 11756
rect 2596 11636 2648 11688
rect 1400 11611 1452 11620
rect 1400 11577 1409 11611
rect 1409 11577 1443 11611
rect 1443 11577 1452 11611
rect 1400 11568 1452 11577
rect 18604 11543 18656 11552
rect 18604 11509 18613 11543
rect 18613 11509 18647 11543
rect 18647 11509 18656 11543
rect 18604 11500 18656 11509
rect 18880 11568 18932 11620
rect 24308 11704 24360 11756
rect 24584 11704 24636 11756
rect 25780 11747 25832 11756
rect 25780 11713 25789 11747
rect 25789 11713 25823 11747
rect 25823 11713 25832 11747
rect 25780 11704 25832 11713
rect 25872 11747 25924 11756
rect 25872 11713 25882 11747
rect 25882 11713 25916 11747
rect 25916 11713 25924 11747
rect 25872 11704 25924 11713
rect 26056 11747 26108 11756
rect 26056 11713 26065 11747
rect 26065 11713 26099 11747
rect 26099 11713 26108 11747
rect 26056 11704 26108 11713
rect 26332 11704 26384 11756
rect 26516 11704 26568 11756
rect 29000 11704 29052 11756
rect 20076 11636 20128 11688
rect 20996 11636 21048 11688
rect 24216 11636 24268 11688
rect 25688 11636 25740 11688
rect 25964 11636 26016 11688
rect 27620 11636 27672 11688
rect 28172 11636 28224 11688
rect 30840 11704 30892 11756
rect 31116 11772 31168 11824
rect 31484 11747 31536 11756
rect 31484 11713 31493 11747
rect 31493 11713 31527 11747
rect 31527 11713 31536 11747
rect 31484 11704 31536 11713
rect 33048 11772 33100 11824
rect 32864 11704 32916 11756
rect 29828 11679 29880 11688
rect 29828 11645 29837 11679
rect 29837 11645 29871 11679
rect 29871 11645 29880 11679
rect 29828 11636 29880 11645
rect 20168 11500 20220 11552
rect 20720 11500 20772 11552
rect 20996 11543 21048 11552
rect 20996 11509 21005 11543
rect 21005 11509 21039 11543
rect 21039 11509 21048 11543
rect 20996 11500 21048 11509
rect 26792 11568 26844 11620
rect 24308 11500 24360 11552
rect 25596 11500 25648 11552
rect 25780 11500 25832 11552
rect 31116 11568 31168 11620
rect 31668 11611 31720 11620
rect 31668 11577 31677 11611
rect 31677 11577 31711 11611
rect 31711 11577 31720 11611
rect 33600 11747 33652 11756
rect 33600 11713 33634 11747
rect 33634 11713 33652 11747
rect 33600 11704 33652 11713
rect 33876 11772 33928 11824
rect 35808 11704 35860 11756
rect 36452 11747 36504 11756
rect 33324 11679 33376 11688
rect 33324 11645 33333 11679
rect 33333 11645 33367 11679
rect 33367 11645 33376 11679
rect 36452 11713 36461 11747
rect 36461 11713 36495 11747
rect 36495 11713 36504 11747
rect 36452 11704 36504 11713
rect 36728 11747 36780 11756
rect 36728 11713 36737 11747
rect 36737 11713 36771 11747
rect 36771 11713 36780 11747
rect 37372 11840 37424 11892
rect 37280 11815 37332 11824
rect 37280 11781 37289 11815
rect 37289 11781 37323 11815
rect 37323 11781 37332 11815
rect 37280 11772 37332 11781
rect 43812 11840 43864 11892
rect 38384 11772 38436 11824
rect 36728 11704 36780 11713
rect 36268 11679 36320 11688
rect 33324 11636 33376 11645
rect 31668 11568 31720 11577
rect 29184 11500 29236 11552
rect 32588 11543 32640 11552
rect 32588 11509 32597 11543
rect 32597 11509 32631 11543
rect 32631 11509 32640 11543
rect 32588 11500 32640 11509
rect 32772 11500 32824 11552
rect 36268 11645 36277 11679
rect 36277 11645 36311 11679
rect 36311 11645 36320 11679
rect 36268 11636 36320 11645
rect 36636 11679 36688 11688
rect 36636 11645 36645 11679
rect 36645 11645 36679 11679
rect 36679 11645 36688 11679
rect 36636 11636 36688 11645
rect 37004 11636 37056 11688
rect 38200 11636 38252 11688
rect 38476 11636 38528 11688
rect 39672 11704 39724 11756
rect 40224 11747 40276 11756
rect 40224 11713 40233 11747
rect 40233 11713 40267 11747
rect 40267 11713 40276 11747
rect 40224 11704 40276 11713
rect 40408 11704 40460 11756
rect 41604 11772 41656 11824
rect 43720 11772 43772 11824
rect 44640 11840 44692 11892
rect 44732 11840 44784 11892
rect 46112 11840 46164 11892
rect 47584 11883 47636 11892
rect 47584 11849 47593 11883
rect 47593 11849 47627 11883
rect 47627 11849 47636 11883
rect 47584 11840 47636 11849
rect 47676 11840 47728 11892
rect 48136 11840 48188 11892
rect 48596 11840 48648 11892
rect 49608 11840 49660 11892
rect 44824 11772 44876 11824
rect 45100 11815 45152 11824
rect 45100 11781 45134 11815
rect 45134 11781 45152 11815
rect 45100 11772 45152 11781
rect 45560 11772 45612 11824
rect 38936 11636 38988 11688
rect 39396 11679 39448 11688
rect 39396 11645 39405 11679
rect 39405 11645 39439 11679
rect 39439 11645 39448 11679
rect 39396 11636 39448 11645
rect 39856 11636 39908 11688
rect 40592 11636 40644 11688
rect 40776 11636 40828 11688
rect 40960 11636 41012 11688
rect 43628 11636 43680 11688
rect 44180 11747 44232 11756
rect 44180 11713 44189 11747
rect 44189 11713 44223 11747
rect 44223 11713 44232 11747
rect 44180 11704 44232 11713
rect 44364 11704 44416 11756
rect 46112 11704 46164 11756
rect 46756 11747 46808 11756
rect 46756 11713 46765 11747
rect 46765 11713 46799 11747
rect 46799 11713 46808 11747
rect 46756 11704 46808 11713
rect 47216 11704 47268 11756
rect 47860 11772 47912 11824
rect 48228 11772 48280 11824
rect 49884 11840 49936 11892
rect 35440 11611 35492 11620
rect 35440 11577 35449 11611
rect 35449 11577 35483 11611
rect 35483 11577 35492 11611
rect 35440 11568 35492 11577
rect 36728 11568 36780 11620
rect 35992 11500 36044 11552
rect 36176 11500 36228 11552
rect 36912 11500 36964 11552
rect 37188 11568 37240 11620
rect 37372 11568 37424 11620
rect 37556 11568 37608 11620
rect 38292 11568 38344 11620
rect 38752 11568 38804 11620
rect 44088 11568 44140 11620
rect 39028 11500 39080 11552
rect 40316 11500 40368 11552
rect 40776 11500 40828 11552
rect 41144 11500 41196 11552
rect 44180 11500 44232 11552
rect 44456 11543 44508 11552
rect 44456 11509 44465 11543
rect 44465 11509 44499 11543
rect 44499 11509 44508 11543
rect 44456 11500 44508 11509
rect 49516 11636 49568 11688
rect 49976 11747 50028 11756
rect 49976 11713 49985 11747
rect 49985 11713 50019 11747
rect 50019 11713 50028 11747
rect 50344 11747 50396 11756
rect 49976 11704 50028 11713
rect 50344 11713 50353 11747
rect 50353 11713 50387 11747
rect 50387 11713 50396 11747
rect 50344 11704 50396 11713
rect 52092 11883 52144 11892
rect 51080 11772 51132 11824
rect 52092 11849 52101 11883
rect 52101 11849 52135 11883
rect 52135 11849 52144 11883
rect 52092 11840 52144 11849
rect 52736 11883 52788 11892
rect 52736 11849 52745 11883
rect 52745 11849 52779 11883
rect 52779 11849 52788 11883
rect 52736 11840 52788 11849
rect 53196 11840 53248 11892
rect 53380 11840 53432 11892
rect 54668 11840 54720 11892
rect 54760 11883 54812 11892
rect 54760 11849 54769 11883
rect 54769 11849 54803 11883
rect 54803 11849 54812 11883
rect 54760 11840 54812 11849
rect 56508 11840 56560 11892
rect 51356 11704 51408 11756
rect 52000 11704 52052 11756
rect 52828 11704 52880 11756
rect 53748 11747 53800 11756
rect 53748 11713 53757 11747
rect 53757 11713 53791 11747
rect 53791 11713 53800 11747
rect 53748 11704 53800 11713
rect 53932 11747 53984 11756
rect 53932 11713 53941 11747
rect 53941 11713 53975 11747
rect 53975 11713 53984 11747
rect 53932 11704 53984 11713
rect 54208 11772 54260 11824
rect 56968 11815 57020 11824
rect 54116 11704 54168 11756
rect 56968 11781 56977 11815
rect 56977 11781 57011 11815
rect 57011 11781 57020 11815
rect 56968 11772 57020 11781
rect 57060 11772 57112 11824
rect 57520 11772 57572 11824
rect 58900 11815 58952 11824
rect 55220 11747 55272 11756
rect 46112 11568 46164 11620
rect 49884 11568 49936 11620
rect 54760 11636 54812 11688
rect 55220 11713 55229 11747
rect 55229 11713 55263 11747
rect 55263 11713 55272 11747
rect 55220 11704 55272 11713
rect 55128 11636 55180 11688
rect 55772 11704 55824 11756
rect 57152 11747 57204 11756
rect 57152 11713 57161 11747
rect 57161 11713 57195 11747
rect 57195 11713 57204 11747
rect 57152 11704 57204 11713
rect 57888 11747 57940 11756
rect 56508 11636 56560 11688
rect 57888 11713 57897 11747
rect 57897 11713 57931 11747
rect 57931 11713 57940 11747
rect 57888 11704 57940 11713
rect 58348 11704 58400 11756
rect 58900 11781 58909 11815
rect 58909 11781 58943 11815
rect 58943 11781 58952 11815
rect 58900 11772 58952 11781
rect 59176 11772 59228 11824
rect 60556 11840 60608 11892
rect 61108 11840 61160 11892
rect 61200 11840 61252 11892
rect 59084 11747 59136 11756
rect 59084 11713 59087 11747
rect 59087 11713 59136 11747
rect 58532 11636 58584 11688
rect 59084 11704 59136 11713
rect 59360 11704 59412 11756
rect 60004 11747 60056 11756
rect 60004 11713 60013 11747
rect 60013 11713 60047 11747
rect 60047 11713 60056 11747
rect 60004 11704 60056 11713
rect 62948 11772 63000 11824
rect 63592 11772 63644 11824
rect 60832 11679 60884 11688
rect 60832 11645 60841 11679
rect 60841 11645 60875 11679
rect 60875 11645 60884 11679
rect 60832 11636 60884 11645
rect 63408 11704 63460 11756
rect 62120 11636 62172 11688
rect 63592 11679 63644 11688
rect 63592 11645 63601 11679
rect 63601 11645 63635 11679
rect 63635 11645 63644 11679
rect 63592 11636 63644 11645
rect 64788 11840 64840 11892
rect 64880 11840 64932 11892
rect 66812 11840 66864 11892
rect 67180 11840 67232 11892
rect 67272 11840 67324 11892
rect 67548 11840 67600 11892
rect 69112 11840 69164 11892
rect 69204 11840 69256 11892
rect 69848 11840 69900 11892
rect 70032 11840 70084 11892
rect 71320 11840 71372 11892
rect 72332 11840 72384 11892
rect 65156 11772 65208 11824
rect 64052 11747 64104 11756
rect 64052 11713 64061 11747
rect 64061 11713 64095 11747
rect 64095 11713 64104 11747
rect 64052 11704 64104 11713
rect 64696 11747 64748 11756
rect 64696 11713 64705 11747
rect 64705 11713 64739 11747
rect 64739 11713 64748 11747
rect 64696 11704 64748 11713
rect 66996 11772 67048 11824
rect 66168 11747 66220 11756
rect 66168 11713 66177 11747
rect 66177 11713 66211 11747
rect 66211 11713 66220 11747
rect 66168 11704 66220 11713
rect 66260 11704 66312 11756
rect 68836 11772 68888 11824
rect 70860 11815 70912 11824
rect 70860 11781 70869 11815
rect 70869 11781 70903 11815
rect 70903 11781 70912 11815
rect 70860 11772 70912 11781
rect 67364 11704 67416 11756
rect 67548 11636 67600 11688
rect 68928 11747 68980 11756
rect 68928 11713 68937 11747
rect 68937 11713 68971 11747
rect 68971 11713 68980 11747
rect 68928 11704 68980 11713
rect 69112 11747 69164 11756
rect 69112 11713 69121 11747
rect 69121 11713 69155 11747
rect 69155 11713 69164 11747
rect 69112 11704 69164 11713
rect 69204 11747 69256 11756
rect 69204 11713 69213 11747
rect 69213 11713 69247 11747
rect 69247 11713 69256 11747
rect 69204 11704 69256 11713
rect 71504 11704 71556 11756
rect 88248 11747 88300 11756
rect 50252 11568 50304 11620
rect 45744 11500 45796 11552
rect 45836 11500 45888 11552
rect 47584 11500 47636 11552
rect 51080 11500 51132 11552
rect 51264 11500 51316 11552
rect 51356 11500 51408 11552
rect 52920 11500 52972 11552
rect 53104 11500 53156 11552
rect 54116 11500 54168 11552
rect 54852 11500 54904 11552
rect 56600 11500 56652 11552
rect 57152 11568 57204 11620
rect 58072 11568 58124 11620
rect 60556 11568 60608 11620
rect 61936 11568 61988 11620
rect 67180 11568 67232 11620
rect 67272 11568 67324 11620
rect 58900 11500 58952 11552
rect 59176 11543 59228 11552
rect 59176 11509 59185 11543
rect 59185 11509 59219 11543
rect 59219 11509 59228 11543
rect 59176 11500 59228 11509
rect 59268 11500 59320 11552
rect 61200 11500 61252 11552
rect 61476 11500 61528 11552
rect 62304 11500 62356 11552
rect 63224 11500 63276 11552
rect 64696 11500 64748 11552
rect 67088 11500 67140 11552
rect 71412 11636 71464 11688
rect 88248 11713 88257 11747
rect 88257 11713 88291 11747
rect 88291 11713 88300 11747
rect 88248 11704 88300 11713
rect 88064 11611 88116 11620
rect 88064 11577 88073 11611
rect 88073 11577 88107 11611
rect 88107 11577 88116 11611
rect 88064 11568 88116 11577
rect 70400 11500 70452 11552
rect 11924 11398 11976 11450
rect 11988 11398 12040 11450
rect 12052 11398 12104 11450
rect 12116 11398 12168 11450
rect 12180 11398 12232 11450
rect 33872 11398 33924 11450
rect 33936 11398 33988 11450
rect 34000 11398 34052 11450
rect 34064 11398 34116 11450
rect 34128 11398 34180 11450
rect 55820 11398 55872 11450
rect 55884 11398 55936 11450
rect 55948 11398 56000 11450
rect 56012 11398 56064 11450
rect 56076 11398 56128 11450
rect 77768 11398 77820 11450
rect 77832 11398 77884 11450
rect 77896 11398 77948 11450
rect 77960 11398 78012 11450
rect 78024 11398 78076 11450
rect 4804 11296 4856 11348
rect 14464 11296 14516 11348
rect 14740 11296 14792 11348
rect 24492 11339 24544 11348
rect 24492 11305 24501 11339
rect 24501 11305 24535 11339
rect 24535 11305 24544 11339
rect 24492 11296 24544 11305
rect 24860 11339 24912 11348
rect 24860 11305 24869 11339
rect 24869 11305 24903 11339
rect 24903 11305 24912 11339
rect 24860 11296 24912 11305
rect 27620 11339 27672 11348
rect 27620 11305 27629 11339
rect 27629 11305 27663 11339
rect 27663 11305 27672 11339
rect 27620 11296 27672 11305
rect 34244 11339 34296 11348
rect 25320 11271 25372 11280
rect 25320 11237 25329 11271
rect 25329 11237 25363 11271
rect 25363 11237 25372 11271
rect 25320 11228 25372 11237
rect 26884 11228 26936 11280
rect 18788 11160 18840 11212
rect 23480 11160 23532 11212
rect 23572 11160 23624 11212
rect 29552 11228 29604 11280
rect 31024 11228 31076 11280
rect 34244 11305 34253 11339
rect 34253 11305 34287 11339
rect 34287 11305 34296 11339
rect 34244 11296 34296 11305
rect 35716 11296 35768 11348
rect 35808 11296 35860 11348
rect 38568 11296 38620 11348
rect 38752 11339 38804 11348
rect 38752 11305 38761 11339
rect 38761 11305 38795 11339
rect 38795 11305 38804 11339
rect 38752 11296 38804 11305
rect 38844 11296 38896 11348
rect 39856 11339 39908 11348
rect 39856 11305 39865 11339
rect 39865 11305 39899 11339
rect 39899 11305 39908 11339
rect 39856 11296 39908 11305
rect 40132 11296 40184 11348
rect 41144 11296 41196 11348
rect 41236 11296 41288 11348
rect 39028 11228 39080 11280
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 15844 11092 15896 11144
rect 24216 11092 24268 11144
rect 24308 11024 24360 11076
rect 24584 11092 24636 11144
rect 25780 11135 25832 11144
rect 25780 11101 25789 11135
rect 25789 11101 25823 11135
rect 25823 11101 25832 11135
rect 25780 11092 25832 11101
rect 27160 11092 27212 11144
rect 29460 11160 29512 11212
rect 34980 11160 35032 11212
rect 1400 10999 1452 11008
rect 1400 10965 1409 10999
rect 1409 10965 1443 10999
rect 1443 10965 1452 10999
rect 1400 10956 1452 10965
rect 25044 11024 25096 11076
rect 26240 11024 26292 11076
rect 29184 11092 29236 11144
rect 29552 11135 29604 11144
rect 29552 11101 29561 11135
rect 29561 11101 29595 11135
rect 29595 11101 29604 11135
rect 29552 11092 29604 11101
rect 30748 11092 30800 11144
rect 31760 11135 31812 11144
rect 31760 11101 31769 11135
rect 31769 11101 31803 11135
rect 31803 11101 31812 11135
rect 31760 11092 31812 11101
rect 32496 11092 32548 11144
rect 35716 11092 35768 11144
rect 36544 11160 36596 11212
rect 37740 11160 37792 11212
rect 38200 11203 38252 11212
rect 38200 11169 38210 11203
rect 38210 11169 38244 11203
rect 38244 11169 38252 11203
rect 38200 11160 38252 11169
rect 38476 11160 38528 11212
rect 38844 11160 38896 11212
rect 41696 11271 41748 11280
rect 41696 11237 41705 11271
rect 41705 11237 41739 11271
rect 41739 11237 41748 11271
rect 41696 11228 41748 11237
rect 41880 11228 41932 11280
rect 44732 11296 44784 11348
rect 45100 11296 45152 11348
rect 44088 11228 44140 11280
rect 46112 11228 46164 11280
rect 46388 11296 46440 11348
rect 51172 11296 51224 11348
rect 51356 11296 51408 11348
rect 55128 11296 55180 11348
rect 55588 11296 55640 11348
rect 47584 11271 47636 11280
rect 41144 11160 41196 11212
rect 41328 11203 41380 11212
rect 41328 11169 41337 11203
rect 41337 11169 41371 11203
rect 41371 11169 41380 11203
rect 41328 11160 41380 11169
rect 42248 11160 42300 11212
rect 43076 11160 43128 11212
rect 47584 11237 47593 11271
rect 47593 11237 47627 11271
rect 47627 11237 47636 11271
rect 47584 11228 47636 11237
rect 35992 11135 36044 11144
rect 35992 11101 36001 11135
rect 36001 11101 36035 11135
rect 36035 11101 36044 11135
rect 35992 11092 36044 11101
rect 36084 11135 36136 11144
rect 36084 11101 36093 11135
rect 36093 11101 36127 11135
rect 36127 11101 36136 11135
rect 36084 11092 36136 11101
rect 36452 11092 36504 11144
rect 37096 11092 37148 11144
rect 38108 11135 38160 11144
rect 38108 11101 38117 11135
rect 38117 11101 38151 11135
rect 38151 11101 38160 11135
rect 38108 11092 38160 11101
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38936 11135 38988 11144
rect 38292 11092 38344 11101
rect 38936 11101 38945 11135
rect 38945 11101 38979 11135
rect 38979 11101 38988 11135
rect 38936 11092 38988 11101
rect 39028 11135 39080 11144
rect 39028 11101 39037 11135
rect 39037 11101 39071 11135
rect 39071 11101 39080 11135
rect 39028 11092 39080 11101
rect 39212 11135 39264 11144
rect 39212 11101 39221 11135
rect 39221 11101 39255 11135
rect 39255 11101 39264 11135
rect 40040 11135 40092 11144
rect 39212 11092 39264 11101
rect 40040 11101 40049 11135
rect 40049 11101 40083 11135
rect 40083 11101 40092 11135
rect 40040 11092 40092 11101
rect 40224 11092 40276 11144
rect 40868 11092 40920 11144
rect 41788 11092 41840 11144
rect 41972 11135 42024 11144
rect 41972 11101 41981 11135
rect 41981 11101 42015 11135
rect 42015 11101 42024 11135
rect 41972 11092 42024 11101
rect 42340 11092 42392 11144
rect 44272 11135 44324 11144
rect 44272 11101 44281 11135
rect 44281 11101 44315 11135
rect 44315 11101 44324 11135
rect 44272 11092 44324 11101
rect 44364 11135 44416 11144
rect 44364 11101 44373 11135
rect 44373 11101 44407 11135
rect 44407 11101 44416 11135
rect 44364 11092 44416 11101
rect 45560 11092 45612 11144
rect 46020 11135 46072 11144
rect 46020 11101 46029 11135
rect 46029 11101 46063 11135
rect 46063 11101 46072 11135
rect 46020 11092 46072 11101
rect 46204 11092 46256 11144
rect 46664 11135 46716 11144
rect 46664 11101 46673 11135
rect 46673 11101 46707 11135
rect 46707 11101 46716 11135
rect 46664 11092 46716 11101
rect 46756 11092 46808 11144
rect 47216 11092 47268 11144
rect 49240 11160 49292 11212
rect 49976 11228 50028 11280
rect 53932 11228 53984 11280
rect 49424 11135 49476 11144
rect 49424 11101 49433 11135
rect 49433 11101 49467 11135
rect 49467 11101 49476 11135
rect 49424 11092 49476 11101
rect 49792 11092 49844 11144
rect 25872 10956 25924 11008
rect 27160 10999 27212 11008
rect 27160 10965 27169 10999
rect 27169 10965 27203 10999
rect 27203 10965 27212 10999
rect 27160 10956 27212 10965
rect 27344 10956 27396 11008
rect 33140 11067 33192 11076
rect 33140 11033 33174 11067
rect 33174 11033 33192 11067
rect 33140 11024 33192 11033
rect 33232 11024 33284 11076
rect 37556 11024 37608 11076
rect 30012 10956 30064 11008
rect 32772 10956 32824 11008
rect 35072 10999 35124 11008
rect 35072 10965 35081 10999
rect 35081 10965 35115 10999
rect 35115 10965 35124 10999
rect 35072 10956 35124 10965
rect 35164 10956 35216 11008
rect 37740 10956 37792 11008
rect 38568 11024 38620 11076
rect 41328 11024 41380 11076
rect 41880 11067 41932 11076
rect 41880 11033 41889 11067
rect 41889 11033 41923 11067
rect 41923 11033 41932 11067
rect 41880 11024 41932 11033
rect 44640 11024 44692 11076
rect 49976 11024 50028 11076
rect 50160 11160 50212 11212
rect 50344 11160 50396 11212
rect 52276 11160 52328 11212
rect 57796 11228 57848 11280
rect 60004 11296 60056 11348
rect 60740 11296 60792 11348
rect 61936 11296 61988 11348
rect 62580 11296 62632 11348
rect 62672 11296 62724 11348
rect 67732 11296 67784 11348
rect 69296 11296 69348 11348
rect 73804 11296 73856 11348
rect 62212 11228 62264 11280
rect 55496 11160 55548 11212
rect 50528 11135 50580 11144
rect 50528 11101 50537 11135
rect 50537 11101 50571 11135
rect 50571 11101 50580 11135
rect 50528 11092 50580 11101
rect 50620 11135 50672 11144
rect 50620 11101 50629 11135
rect 50629 11101 50663 11135
rect 50663 11101 50672 11135
rect 50620 11092 50672 11101
rect 53104 11135 53156 11144
rect 53104 11101 53113 11135
rect 53113 11101 53147 11135
rect 53147 11101 53156 11135
rect 53104 11092 53156 11101
rect 55220 11092 55272 11144
rect 56048 11092 56100 11144
rect 56232 11092 56284 11144
rect 58440 11092 58492 11144
rect 59452 11092 59504 11144
rect 52736 11024 52788 11076
rect 52828 11024 52880 11076
rect 54576 11024 54628 11076
rect 54760 11024 54812 11076
rect 56692 11024 56744 11076
rect 57060 11024 57112 11076
rect 58072 11024 58124 11076
rect 58900 11024 58952 11076
rect 60556 11160 60608 11212
rect 60648 11135 60700 11144
rect 60648 11101 60657 11135
rect 60657 11101 60691 11135
rect 60691 11101 60700 11135
rect 60648 11092 60700 11101
rect 59636 11024 59688 11076
rect 61384 11135 61436 11144
rect 61384 11101 61393 11135
rect 61393 11101 61427 11135
rect 61427 11101 61436 11135
rect 61384 11092 61436 11101
rect 63040 11160 63092 11212
rect 65156 11160 65208 11212
rect 61200 11024 61252 11076
rect 62488 11092 62540 11144
rect 62856 11092 62908 11144
rect 40132 10956 40184 11008
rect 40316 10956 40368 11008
rect 41052 10956 41104 11008
rect 41144 10956 41196 11008
rect 61844 10956 61896 11008
rect 61936 10956 61988 11008
rect 63316 11024 63368 11076
rect 64052 11092 64104 11144
rect 64236 11135 64288 11144
rect 64236 11101 64245 11135
rect 64245 11101 64279 11135
rect 64279 11101 64288 11135
rect 64236 11092 64288 11101
rect 64328 11092 64380 11144
rect 64512 11092 64564 11144
rect 67456 11228 67508 11280
rect 67548 11228 67600 11280
rect 69112 11228 69164 11280
rect 69388 11228 69440 11280
rect 73988 11228 74040 11280
rect 67088 11160 67140 11212
rect 67824 11203 67876 11212
rect 67272 11135 67324 11144
rect 67272 11101 67281 11135
rect 67281 11101 67315 11135
rect 67315 11101 67324 11135
rect 67272 11092 67324 11101
rect 67824 11169 67833 11203
rect 67833 11169 67867 11203
rect 67867 11169 67876 11203
rect 67824 11160 67876 11169
rect 62764 10956 62816 11008
rect 67640 11024 67692 11076
rect 69112 11024 69164 11076
rect 87512 11160 87564 11212
rect 87420 11135 87472 11144
rect 87420 11101 87429 11135
rect 87429 11101 87463 11135
rect 87463 11101 87472 11135
rect 87420 11092 87472 11101
rect 67456 10956 67508 11008
rect 87696 10956 87748 11008
rect 22898 10854 22950 10906
rect 22962 10854 23014 10906
rect 23026 10854 23078 10906
rect 23090 10854 23142 10906
rect 23154 10854 23206 10906
rect 44846 10854 44898 10906
rect 44910 10854 44962 10906
rect 44974 10854 45026 10906
rect 45038 10854 45090 10906
rect 45102 10854 45154 10906
rect 66794 10854 66846 10906
rect 66858 10854 66910 10906
rect 66922 10854 66974 10906
rect 66986 10854 67038 10906
rect 67050 10854 67102 10906
rect 20904 10752 20956 10804
rect 26148 10795 26200 10804
rect 26148 10761 26157 10795
rect 26157 10761 26191 10795
rect 26191 10761 26200 10795
rect 26148 10752 26200 10761
rect 29736 10752 29788 10804
rect 30748 10752 30800 10804
rect 31484 10752 31536 10804
rect 33140 10752 33192 10804
rect 33600 10752 33652 10804
rect 33876 10752 33928 10804
rect 35164 10752 35216 10804
rect 37004 10752 37056 10804
rect 37556 10752 37608 10804
rect 38476 10752 38528 10804
rect 40224 10752 40276 10804
rect 87696 10795 87748 10804
rect 27160 10684 27212 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 23388 10548 23440 10600
rect 27068 10616 27120 10668
rect 29000 10659 29052 10668
rect 25872 10548 25924 10600
rect 24492 10480 24544 10532
rect 26424 10480 26476 10532
rect 29000 10625 29009 10659
rect 29009 10625 29043 10659
rect 29043 10625 29052 10659
rect 29000 10616 29052 10625
rect 29828 10684 29880 10736
rect 30288 10684 30340 10736
rect 32496 10684 32548 10736
rect 33784 10684 33836 10736
rect 29276 10616 29328 10668
rect 33508 10616 33560 10668
rect 35072 10684 35124 10736
rect 34244 10659 34296 10668
rect 34244 10625 34253 10659
rect 34253 10625 34287 10659
rect 34287 10625 34296 10659
rect 34244 10616 34296 10625
rect 36268 10616 36320 10668
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 38200 10684 38252 10736
rect 39120 10684 39172 10736
rect 51356 10684 51408 10736
rect 54300 10684 54352 10736
rect 56324 10684 56376 10736
rect 56508 10684 56560 10736
rect 58532 10684 58584 10736
rect 59820 10727 59872 10736
rect 29552 10548 29604 10600
rect 37372 10616 37424 10668
rect 37648 10616 37700 10668
rect 38568 10616 38620 10668
rect 37096 10548 37148 10600
rect 37556 10591 37608 10600
rect 37556 10557 37565 10591
rect 37565 10557 37599 10591
rect 37599 10557 37608 10591
rect 37556 10548 37608 10557
rect 38384 10591 38436 10600
rect 38384 10557 38393 10591
rect 38393 10557 38427 10591
rect 38427 10557 38436 10591
rect 38384 10548 38436 10557
rect 39396 10616 39448 10668
rect 39488 10616 39540 10668
rect 40316 10659 40368 10668
rect 40316 10625 40325 10659
rect 40325 10625 40359 10659
rect 40359 10625 40368 10659
rect 40316 10616 40368 10625
rect 40776 10659 40828 10668
rect 40776 10625 40785 10659
rect 40785 10625 40819 10659
rect 40819 10625 40828 10659
rect 40776 10616 40828 10625
rect 41420 10616 41472 10668
rect 39304 10591 39356 10600
rect 39304 10557 39313 10591
rect 39313 10557 39347 10591
rect 39347 10557 39356 10591
rect 39304 10548 39356 10557
rect 42616 10548 42668 10600
rect 43076 10616 43128 10668
rect 1400 10455 1452 10464
rect 1400 10421 1409 10455
rect 1409 10421 1443 10455
rect 1443 10421 1452 10455
rect 1400 10412 1452 10421
rect 25228 10412 25280 10464
rect 28080 10455 28132 10464
rect 28080 10421 28089 10455
rect 28089 10421 28123 10455
rect 28123 10421 28132 10455
rect 28080 10412 28132 10421
rect 30104 10412 30156 10464
rect 31116 10455 31168 10464
rect 31116 10421 31125 10455
rect 31125 10421 31159 10455
rect 31159 10421 31168 10455
rect 31116 10412 31168 10421
rect 32312 10412 32364 10464
rect 33876 10412 33928 10464
rect 34336 10455 34388 10464
rect 34336 10421 34345 10455
rect 34345 10421 34379 10455
rect 34379 10421 34388 10455
rect 34336 10412 34388 10421
rect 38752 10412 38804 10464
rect 38936 10412 38988 10464
rect 39764 10412 39816 10464
rect 41052 10480 41104 10532
rect 42892 10523 42944 10532
rect 42892 10489 42901 10523
rect 42901 10489 42935 10523
rect 42935 10489 42944 10523
rect 42892 10480 42944 10489
rect 42984 10480 43036 10532
rect 45284 10616 45336 10668
rect 43996 10591 44048 10600
rect 43996 10557 44005 10591
rect 44005 10557 44039 10591
rect 44039 10557 44048 10591
rect 43996 10548 44048 10557
rect 44640 10480 44692 10532
rect 45192 10548 45244 10600
rect 46296 10616 46348 10668
rect 45744 10591 45796 10600
rect 45744 10557 45753 10591
rect 45753 10557 45787 10591
rect 45787 10557 45796 10591
rect 45744 10548 45796 10557
rect 47124 10616 47176 10668
rect 48688 10659 48740 10668
rect 48688 10625 48697 10659
rect 48697 10625 48731 10659
rect 48731 10625 48740 10659
rect 48688 10616 48740 10625
rect 50528 10616 50580 10668
rect 50896 10616 50948 10668
rect 53104 10616 53156 10668
rect 54484 10616 54536 10668
rect 56600 10616 56652 10668
rect 57428 10659 57480 10668
rect 52092 10548 52144 10600
rect 45652 10480 45704 10532
rect 42432 10412 42484 10464
rect 43444 10412 43496 10464
rect 43536 10455 43588 10464
rect 43536 10421 43545 10455
rect 43545 10421 43579 10455
rect 43579 10421 43588 10455
rect 44456 10455 44508 10464
rect 43536 10412 43588 10421
rect 44456 10421 44465 10455
rect 44465 10421 44499 10455
rect 44499 10421 44508 10455
rect 44456 10412 44508 10421
rect 45560 10412 45612 10464
rect 46756 10412 46808 10464
rect 47216 10412 47268 10464
rect 52552 10480 52604 10532
rect 52736 10523 52788 10532
rect 52736 10489 52745 10523
rect 52745 10489 52779 10523
rect 52779 10489 52788 10523
rect 52736 10480 52788 10489
rect 48044 10412 48096 10464
rect 49976 10412 50028 10464
rect 53104 10412 53156 10464
rect 53288 10455 53340 10464
rect 53288 10421 53297 10455
rect 53297 10421 53331 10455
rect 53331 10421 53340 10455
rect 53288 10412 53340 10421
rect 53748 10548 53800 10600
rect 55680 10548 55732 10600
rect 57428 10625 57437 10659
rect 57437 10625 57471 10659
rect 57471 10625 57480 10659
rect 57428 10616 57480 10625
rect 58716 10616 58768 10668
rect 58900 10659 58952 10668
rect 58900 10625 58909 10659
rect 58909 10625 58943 10659
rect 58943 10625 58952 10659
rect 58900 10616 58952 10625
rect 59084 10616 59136 10668
rect 59820 10693 59829 10727
rect 59829 10693 59863 10727
rect 59863 10693 59872 10727
rect 59820 10684 59872 10693
rect 60648 10684 60700 10736
rect 60832 10684 60884 10736
rect 63684 10684 63736 10736
rect 87696 10761 87705 10795
rect 87705 10761 87739 10795
rect 87739 10761 87748 10795
rect 87696 10752 87748 10761
rect 60188 10616 60240 10668
rect 60740 10616 60792 10668
rect 62212 10616 62264 10668
rect 63224 10659 63276 10668
rect 63224 10625 63233 10659
rect 63233 10625 63267 10659
rect 63267 10625 63276 10659
rect 63224 10616 63276 10625
rect 63408 10659 63460 10668
rect 63408 10625 63417 10659
rect 63417 10625 63451 10659
rect 63451 10625 63460 10659
rect 63408 10616 63460 10625
rect 55404 10480 55456 10532
rect 63040 10548 63092 10600
rect 65616 10616 65668 10668
rect 87052 10684 87104 10736
rect 66536 10616 66588 10668
rect 67548 10616 67600 10668
rect 58072 10480 58124 10532
rect 59176 10480 59228 10532
rect 61936 10480 61988 10532
rect 62120 10523 62172 10532
rect 62120 10489 62129 10523
rect 62129 10489 62163 10523
rect 62163 10489 62172 10523
rect 62120 10480 62172 10489
rect 64788 10480 64840 10532
rect 55496 10412 55548 10464
rect 55680 10412 55732 10464
rect 56600 10412 56652 10464
rect 57796 10412 57848 10464
rect 58440 10455 58492 10464
rect 58440 10421 58449 10455
rect 58449 10421 58483 10455
rect 58483 10421 58492 10455
rect 58440 10412 58492 10421
rect 58900 10412 58952 10464
rect 64880 10412 64932 10464
rect 65156 10455 65208 10464
rect 65156 10421 65165 10455
rect 65165 10421 65199 10455
rect 65199 10421 65208 10455
rect 65156 10412 65208 10421
rect 88064 10455 88116 10464
rect 88064 10421 88073 10455
rect 88073 10421 88107 10455
rect 88107 10421 88116 10455
rect 88064 10412 88116 10421
rect 11924 10310 11976 10362
rect 11988 10310 12040 10362
rect 12052 10310 12104 10362
rect 12116 10310 12168 10362
rect 12180 10310 12232 10362
rect 33872 10310 33924 10362
rect 33936 10310 33988 10362
rect 34000 10310 34052 10362
rect 34064 10310 34116 10362
rect 34128 10310 34180 10362
rect 55820 10310 55872 10362
rect 55884 10310 55936 10362
rect 55948 10310 56000 10362
rect 56012 10310 56064 10362
rect 56076 10310 56128 10362
rect 77768 10310 77820 10362
rect 77832 10310 77884 10362
rect 77896 10310 77948 10362
rect 77960 10310 78012 10362
rect 78024 10310 78076 10362
rect 25044 10251 25096 10260
rect 25044 10217 25053 10251
rect 25053 10217 25087 10251
rect 25087 10217 25096 10251
rect 25044 10208 25096 10217
rect 29276 10208 29328 10260
rect 32496 10208 32548 10260
rect 33508 10208 33560 10260
rect 34244 10208 34296 10260
rect 34336 10208 34388 10260
rect 33784 10072 33836 10124
rect 35164 10140 35216 10192
rect 38108 10208 38160 10260
rect 38844 10208 38896 10260
rect 39212 10208 39264 10260
rect 40316 10208 40368 10260
rect 42248 10208 42300 10260
rect 42892 10208 42944 10260
rect 44456 10208 44508 10260
rect 47124 10208 47176 10260
rect 41972 10140 42024 10192
rect 21548 10004 21600 10056
rect 25228 10047 25280 10056
rect 25228 10013 25237 10047
rect 25237 10013 25271 10047
rect 25271 10013 25280 10047
rect 25228 10004 25280 10013
rect 29092 10047 29144 10056
rect 29092 10013 29101 10047
rect 29101 10013 29135 10047
rect 29135 10013 29144 10047
rect 29092 10004 29144 10013
rect 29552 10047 29604 10056
rect 29552 10013 29561 10047
rect 29561 10013 29595 10047
rect 29595 10013 29604 10047
rect 29552 10004 29604 10013
rect 31760 10004 31812 10056
rect 33232 10004 33284 10056
rect 34520 10004 34572 10056
rect 34888 10047 34940 10056
rect 34888 10013 34897 10047
rect 34897 10013 34931 10047
rect 34931 10013 34940 10047
rect 34888 10004 34940 10013
rect 28080 9936 28132 9988
rect 39304 10072 39356 10124
rect 35992 10047 36044 10056
rect 35992 10013 36001 10047
rect 36001 10013 36035 10047
rect 36035 10013 36044 10047
rect 35992 10004 36044 10013
rect 37556 10004 37608 10056
rect 40040 10047 40092 10056
rect 40040 10013 40049 10047
rect 40049 10013 40083 10047
rect 40083 10013 40092 10047
rect 40040 10004 40092 10013
rect 40132 10004 40184 10056
rect 1400 9911 1452 9920
rect 1400 9877 1409 9911
rect 1409 9877 1443 9911
rect 1443 9877 1452 9911
rect 1400 9868 1452 9877
rect 29000 9868 29052 9920
rect 34612 9868 34664 9920
rect 35808 9911 35860 9920
rect 35808 9877 35817 9911
rect 35817 9877 35851 9911
rect 35851 9877 35860 9911
rect 35808 9868 35860 9877
rect 38660 9936 38712 9988
rect 42800 10004 42852 10056
rect 45284 10140 45336 10192
rect 46664 10183 46716 10192
rect 46664 10149 46673 10183
rect 46673 10149 46707 10183
rect 46707 10149 46716 10183
rect 49700 10208 49752 10260
rect 51908 10208 51960 10260
rect 55496 10208 55548 10260
rect 46664 10140 46716 10149
rect 38108 9868 38160 9920
rect 38200 9868 38252 9920
rect 38844 9868 38896 9920
rect 41696 9936 41748 9988
rect 39304 9868 39356 9920
rect 42708 9936 42760 9988
rect 45376 10004 45428 10056
rect 49792 10140 49844 10192
rect 53104 10140 53156 10192
rect 55220 10140 55272 10192
rect 57428 10208 57480 10260
rect 60740 10208 60792 10260
rect 64604 10208 64656 10260
rect 65616 10208 65668 10260
rect 45560 9979 45612 9988
rect 45560 9945 45594 9979
rect 45594 9945 45612 9979
rect 45560 9936 45612 9945
rect 45652 9936 45704 9988
rect 46756 9936 46808 9988
rect 49976 10072 50028 10124
rect 53748 10115 53800 10124
rect 48964 10047 49016 10056
rect 48964 10013 48973 10047
rect 48973 10013 49007 10047
rect 49007 10013 49016 10047
rect 48964 10004 49016 10013
rect 42984 9868 43036 9920
rect 43444 9868 43496 9920
rect 47216 9911 47268 9920
rect 47216 9877 47241 9911
rect 47241 9877 47268 9911
rect 47216 9868 47268 9877
rect 47492 9868 47544 9920
rect 50068 10004 50120 10056
rect 53748 10081 53757 10115
rect 53757 10081 53791 10115
rect 53791 10081 53800 10115
rect 53748 10072 53800 10081
rect 53840 10072 53892 10124
rect 55036 10072 55088 10124
rect 55312 10115 55364 10124
rect 55312 10081 55321 10115
rect 55321 10081 55355 10115
rect 55355 10081 55364 10115
rect 55312 10072 55364 10081
rect 61936 10140 61988 10192
rect 86592 10208 86644 10260
rect 50988 10004 51040 10056
rect 51356 10004 51408 10056
rect 52184 10004 52236 10056
rect 53104 10004 53156 10056
rect 57796 10047 57848 10056
rect 49608 9936 49660 9988
rect 49700 9868 49752 9920
rect 50528 9911 50580 9920
rect 50528 9877 50537 9911
rect 50537 9877 50571 9911
rect 50571 9877 50580 9911
rect 50528 9868 50580 9877
rect 54392 9868 54444 9920
rect 54576 9911 54628 9920
rect 54576 9877 54585 9911
rect 54585 9877 54619 9911
rect 54619 9877 54628 9911
rect 54576 9868 54628 9877
rect 55404 9936 55456 9988
rect 57796 10013 57805 10047
rect 57805 10013 57839 10047
rect 57839 10013 57848 10047
rect 57796 10004 57848 10013
rect 56232 9868 56284 9920
rect 57244 9868 57296 9920
rect 58164 9936 58216 9988
rect 59176 10004 59228 10056
rect 58624 9868 58676 9920
rect 59820 9911 59872 9920
rect 59820 9877 59829 9911
rect 59829 9877 59863 9911
rect 59863 9877 59872 9911
rect 59820 9868 59872 9877
rect 64696 10072 64748 10124
rect 60832 10047 60884 10056
rect 60832 10013 60841 10047
rect 60841 10013 60875 10047
rect 60875 10013 60884 10047
rect 60832 10004 60884 10013
rect 62304 10004 62356 10056
rect 64236 10004 64288 10056
rect 64788 10004 64840 10056
rect 69020 9936 69072 9988
rect 60924 9911 60976 9920
rect 60924 9877 60933 9911
rect 60933 9877 60967 9911
rect 60967 9877 60976 9911
rect 60924 9868 60976 9877
rect 22898 9766 22950 9818
rect 22962 9766 23014 9818
rect 23026 9766 23078 9818
rect 23090 9766 23142 9818
rect 23154 9766 23206 9818
rect 44846 9766 44898 9818
rect 44910 9766 44962 9818
rect 44974 9766 45026 9818
rect 45038 9766 45090 9818
rect 45102 9766 45154 9818
rect 66794 9766 66846 9818
rect 66858 9766 66910 9818
rect 66922 9766 66974 9818
rect 66986 9766 67038 9818
rect 67050 9766 67102 9818
rect 29092 9664 29144 9716
rect 30288 9664 30340 9716
rect 32588 9664 32640 9716
rect 34520 9664 34572 9716
rect 36268 9664 36320 9716
rect 37648 9707 37700 9716
rect 37648 9673 37657 9707
rect 37657 9673 37691 9707
rect 37691 9673 37700 9707
rect 37648 9664 37700 9673
rect 38384 9664 38436 9716
rect 49424 9664 49476 9716
rect 33508 9639 33560 9648
rect 33508 9605 33517 9639
rect 33517 9605 33551 9639
rect 33551 9605 33560 9639
rect 33508 9596 33560 9605
rect 15384 9528 15436 9580
rect 31116 9528 31168 9580
rect 34612 9596 34664 9648
rect 35164 9571 35216 9580
rect 35164 9537 35173 9571
rect 35173 9537 35207 9571
rect 35207 9537 35216 9571
rect 35164 9528 35216 9537
rect 35808 9596 35860 9648
rect 38292 9596 38344 9648
rect 35716 9528 35768 9580
rect 30196 9503 30248 9512
rect 30196 9469 30205 9503
rect 30205 9469 30239 9503
rect 30239 9469 30248 9503
rect 30196 9460 30248 9469
rect 30288 9503 30340 9512
rect 30288 9469 30297 9503
rect 30297 9469 30331 9503
rect 30331 9469 30340 9503
rect 30288 9460 30340 9469
rect 23572 9392 23624 9444
rect 33784 9503 33836 9512
rect 33784 9469 33793 9503
rect 33793 9469 33827 9503
rect 33827 9469 33836 9503
rect 33784 9460 33836 9469
rect 37556 9528 37608 9580
rect 38016 9528 38068 9580
rect 47400 9596 47452 9648
rect 38844 9571 38896 9580
rect 38844 9537 38878 9571
rect 38878 9537 38896 9571
rect 40316 9571 40368 9580
rect 38844 9528 38896 9537
rect 40316 9537 40325 9571
rect 40325 9537 40359 9571
rect 40359 9537 40368 9571
rect 40316 9528 40368 9537
rect 40408 9528 40460 9580
rect 42892 9528 42944 9580
rect 44088 9528 44140 9580
rect 45836 9528 45888 9580
rect 49700 9664 49752 9716
rect 49792 9664 49844 9716
rect 50804 9664 50856 9716
rect 50988 9707 51040 9716
rect 50988 9673 50997 9707
rect 50997 9673 51031 9707
rect 51031 9673 51040 9707
rect 50988 9664 51040 9673
rect 54300 9664 54352 9716
rect 54484 9707 54536 9716
rect 54484 9673 54493 9707
rect 54493 9673 54527 9707
rect 54527 9673 54536 9707
rect 54484 9664 54536 9673
rect 54576 9664 54628 9716
rect 50160 9596 50212 9648
rect 50528 9596 50580 9648
rect 51172 9596 51224 9648
rect 53748 9596 53800 9648
rect 55036 9596 55088 9648
rect 55680 9664 55732 9716
rect 59268 9664 59320 9716
rect 60832 9707 60884 9716
rect 60832 9673 60841 9707
rect 60841 9673 60875 9707
rect 60875 9673 60884 9707
rect 60832 9664 60884 9673
rect 64696 9664 64748 9716
rect 42984 9503 43036 9512
rect 34888 9392 34940 9444
rect 42984 9469 42993 9503
rect 42993 9469 43027 9503
rect 43027 9469 43036 9503
rect 42984 9460 43036 9469
rect 45560 9460 45612 9512
rect 52736 9571 52788 9580
rect 52736 9537 52745 9571
rect 52745 9537 52779 9571
rect 52779 9537 52788 9571
rect 52736 9528 52788 9537
rect 53288 9528 53340 9580
rect 59820 9596 59872 9648
rect 64236 9639 64288 9648
rect 64236 9605 64245 9639
rect 64245 9605 64279 9639
rect 64279 9605 64288 9639
rect 64236 9596 64288 9605
rect 57244 9571 57296 9580
rect 43996 9392 44048 9444
rect 38568 9324 38620 9376
rect 39304 9324 39356 9376
rect 40224 9324 40276 9376
rect 41696 9367 41748 9376
rect 41696 9333 41705 9367
rect 41705 9333 41739 9367
rect 41739 9333 41748 9367
rect 41696 9324 41748 9333
rect 47492 9392 47544 9444
rect 46388 9324 46440 9376
rect 48596 9324 48648 9376
rect 52644 9324 52696 9376
rect 57244 9537 57253 9571
rect 57253 9537 57287 9571
rect 57287 9537 57296 9571
rect 57244 9528 57296 9537
rect 59452 9571 59504 9580
rect 59452 9537 59461 9571
rect 59461 9537 59495 9571
rect 59495 9537 59504 9571
rect 59452 9528 59504 9537
rect 68192 9528 68244 9580
rect 53104 9324 53156 9376
rect 63408 9460 63460 9512
rect 57060 9435 57112 9444
rect 57060 9401 57069 9435
rect 57069 9401 57103 9435
rect 57103 9401 57112 9435
rect 57060 9392 57112 9401
rect 67548 9460 67600 9512
rect 63408 9324 63460 9376
rect 65156 9324 65208 9376
rect 68284 9324 68336 9376
rect 11924 9222 11976 9274
rect 11988 9222 12040 9274
rect 12052 9222 12104 9274
rect 12116 9222 12168 9274
rect 12180 9222 12232 9274
rect 33872 9222 33924 9274
rect 33936 9222 33988 9274
rect 34000 9222 34052 9274
rect 34064 9222 34116 9274
rect 34128 9222 34180 9274
rect 55820 9222 55872 9274
rect 55884 9222 55936 9274
rect 55948 9222 56000 9274
rect 56012 9222 56064 9274
rect 56076 9222 56128 9274
rect 77768 9222 77820 9274
rect 77832 9222 77884 9274
rect 77896 9222 77948 9274
rect 77960 9222 78012 9274
rect 78024 9222 78076 9274
rect 35992 9120 36044 9172
rect 37372 9163 37424 9172
rect 37372 9129 37381 9163
rect 37381 9129 37415 9163
rect 37415 9129 37424 9163
rect 37372 9120 37424 9129
rect 38844 9120 38896 9172
rect 40868 9120 40920 9172
rect 41328 9120 41380 9172
rect 44088 9163 44140 9172
rect 33784 8984 33836 9036
rect 37740 9052 37792 9104
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 36268 8916 36320 8968
rect 37556 8959 37608 8968
rect 37556 8925 37565 8959
rect 37565 8925 37599 8959
rect 37599 8925 37608 8959
rect 37556 8916 37608 8925
rect 37648 8916 37700 8968
rect 40132 8984 40184 9036
rect 40316 8984 40368 9036
rect 42708 9027 42760 9036
rect 42708 8993 42717 9027
rect 42717 8993 42751 9027
rect 42751 8993 42760 9027
rect 42708 8984 42760 8993
rect 44088 9129 44097 9163
rect 44097 9129 44131 9163
rect 44131 9129 44140 9163
rect 44088 9120 44140 9129
rect 45836 9163 45888 9172
rect 45836 9129 45845 9163
rect 45845 9129 45879 9163
rect 45879 9129 45888 9163
rect 45836 9120 45888 9129
rect 48136 9163 48188 9172
rect 48136 9129 48145 9163
rect 48145 9129 48179 9163
rect 48179 9129 48188 9163
rect 48136 9120 48188 9129
rect 48412 9120 48464 9172
rect 55404 9120 55456 9172
rect 68192 9163 68244 9172
rect 68192 9129 68201 9163
rect 68201 9129 68235 9163
rect 68235 9129 68244 9163
rect 68192 9120 68244 9129
rect 31116 8848 31168 8900
rect 38752 8916 38804 8968
rect 42800 8916 42852 8968
rect 46112 8916 46164 8968
rect 46388 8959 46440 8968
rect 46388 8925 46397 8959
rect 46397 8925 46431 8959
rect 46431 8925 46440 8959
rect 46388 8916 46440 8925
rect 48412 8916 48464 8968
rect 48596 8984 48648 9036
rect 52736 9027 52788 9036
rect 52736 8993 52745 9027
rect 52745 8993 52779 9027
rect 52779 8993 52788 9027
rect 52736 8984 52788 8993
rect 48964 8916 49016 8968
rect 50160 8959 50212 8968
rect 50160 8925 50169 8959
rect 50169 8925 50203 8959
rect 50203 8925 50212 8959
rect 50160 8916 50212 8925
rect 50252 8916 50304 8968
rect 52368 8959 52420 8968
rect 52368 8925 52377 8959
rect 52377 8925 52411 8959
rect 52411 8925 52420 8959
rect 52368 8916 52420 8925
rect 55220 8916 55272 8968
rect 23388 8780 23440 8832
rect 36728 8823 36780 8832
rect 36728 8789 36737 8823
rect 36737 8789 36771 8823
rect 36771 8789 36780 8823
rect 36728 8780 36780 8789
rect 46480 8848 46532 8900
rect 46940 8848 46992 8900
rect 50068 8780 50120 8832
rect 50804 8780 50856 8832
rect 60924 9052 60976 9104
rect 67548 8984 67600 9036
rect 68284 8916 68336 8968
rect 87420 8959 87472 8968
rect 87420 8925 87429 8959
rect 87429 8925 87463 8959
rect 87463 8925 87472 8959
rect 87420 8916 87472 8925
rect 86408 8848 86460 8900
rect 53104 8780 53156 8832
rect 70768 8780 70820 8832
rect 22898 8678 22950 8730
rect 22962 8678 23014 8730
rect 23026 8678 23078 8730
rect 23090 8678 23142 8730
rect 23154 8678 23206 8730
rect 44846 8678 44898 8730
rect 44910 8678 44962 8730
rect 44974 8678 45026 8730
rect 45038 8678 45090 8730
rect 45102 8678 45154 8730
rect 66794 8678 66846 8730
rect 66858 8678 66910 8730
rect 66922 8678 66974 8730
rect 66986 8678 67038 8730
rect 67050 8678 67102 8730
rect 40408 8576 40460 8628
rect 42800 8619 42852 8628
rect 42800 8585 42809 8619
rect 42809 8585 42843 8619
rect 42843 8585 42852 8619
rect 42800 8576 42852 8585
rect 44088 8576 44140 8628
rect 46112 8619 46164 8628
rect 46112 8585 46121 8619
rect 46121 8585 46155 8619
rect 46155 8585 46164 8619
rect 46112 8576 46164 8585
rect 47492 8576 47544 8628
rect 48412 8576 48464 8628
rect 39028 8508 39080 8560
rect 50068 8576 50120 8628
rect 50252 8619 50304 8628
rect 50252 8585 50261 8619
rect 50261 8585 50295 8619
rect 50295 8585 50304 8619
rect 50252 8576 50304 8585
rect 52368 8576 52420 8628
rect 53104 8619 53156 8628
rect 53104 8585 53113 8619
rect 53113 8585 53147 8619
rect 53147 8585 53156 8619
rect 53104 8576 53156 8585
rect 27436 8440 27488 8492
rect 38200 8483 38252 8492
rect 38200 8449 38209 8483
rect 38209 8449 38243 8483
rect 38243 8449 38252 8483
rect 38200 8440 38252 8449
rect 41328 8440 41380 8492
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 33692 8372 33744 8424
rect 41420 8415 41472 8424
rect 41420 8381 41429 8415
rect 41429 8381 41463 8415
rect 41463 8381 41472 8415
rect 41420 8372 41472 8381
rect 42064 8372 42116 8424
rect 43536 8440 43588 8492
rect 45744 8372 45796 8424
rect 48596 8440 48648 8492
rect 67548 8508 67600 8560
rect 49608 8415 49660 8424
rect 39304 8304 39356 8356
rect 49608 8381 49617 8415
rect 49617 8381 49651 8415
rect 49651 8381 49660 8415
rect 49608 8372 49660 8381
rect 55588 8440 55640 8492
rect 88248 8483 88300 8492
rect 88248 8449 88257 8483
rect 88257 8449 88291 8483
rect 88291 8449 88300 8483
rect 88248 8440 88300 8449
rect 50804 8304 50856 8356
rect 82820 8304 82872 8356
rect 41880 8236 41932 8288
rect 11924 8134 11976 8186
rect 11988 8134 12040 8186
rect 12052 8134 12104 8186
rect 12116 8134 12168 8186
rect 12180 8134 12232 8186
rect 33872 8134 33924 8186
rect 33936 8134 33988 8186
rect 34000 8134 34052 8186
rect 34064 8134 34116 8186
rect 34128 8134 34180 8186
rect 55820 8134 55872 8186
rect 55884 8134 55936 8186
rect 55948 8134 56000 8186
rect 56012 8134 56064 8186
rect 56076 8134 56128 8186
rect 77768 8134 77820 8186
rect 77832 8134 77884 8186
rect 77896 8134 77948 8186
rect 77960 8134 78012 8186
rect 78024 8134 78076 8186
rect 46480 8075 46532 8084
rect 46480 8041 46489 8075
rect 46489 8041 46523 8075
rect 46523 8041 46532 8075
rect 46480 8032 46532 8041
rect 41880 7871 41932 7880
rect 41880 7837 41889 7871
rect 41889 7837 41923 7871
rect 41923 7837 41932 7871
rect 41880 7828 41932 7837
rect 48136 7828 48188 7880
rect 64328 7828 64380 7880
rect 20812 7760 20864 7812
rect 58440 7760 58492 7812
rect 1676 7692 1728 7744
rect 34428 7692 34480 7744
rect 41972 7692 42024 7744
rect 88064 7735 88116 7744
rect 88064 7701 88073 7735
rect 88073 7701 88107 7735
rect 88107 7701 88116 7735
rect 88064 7692 88116 7701
rect 22898 7590 22950 7642
rect 22962 7590 23014 7642
rect 23026 7590 23078 7642
rect 23090 7590 23142 7642
rect 23154 7590 23206 7642
rect 44846 7590 44898 7642
rect 44910 7590 44962 7642
rect 44974 7590 45026 7642
rect 45038 7590 45090 7642
rect 45102 7590 45154 7642
rect 66794 7590 66846 7642
rect 66858 7590 66910 7642
rect 66922 7590 66974 7642
rect 66986 7590 67038 7642
rect 67050 7590 67102 7642
rect 40316 7531 40368 7540
rect 40316 7497 40325 7531
rect 40325 7497 40359 7531
rect 40359 7497 40368 7531
rect 40316 7488 40368 7497
rect 38660 7420 38712 7472
rect 18604 7352 18656 7404
rect 88064 7395 88116 7404
rect 88064 7361 88073 7395
rect 88073 7361 88107 7395
rect 88107 7361 88116 7395
rect 88064 7352 88116 7361
rect 36728 7216 36780 7268
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 11924 7046 11976 7098
rect 11988 7046 12040 7098
rect 12052 7046 12104 7098
rect 12116 7046 12168 7098
rect 12180 7046 12232 7098
rect 33872 7046 33924 7098
rect 33936 7046 33988 7098
rect 34000 7046 34052 7098
rect 34064 7046 34116 7098
rect 34128 7046 34180 7098
rect 55820 7046 55872 7098
rect 55884 7046 55936 7098
rect 55948 7046 56000 7098
rect 56012 7046 56064 7098
rect 56076 7046 56128 7098
rect 77768 7046 77820 7098
rect 77832 7046 77884 7098
rect 77896 7046 77948 7098
rect 77960 7046 78012 7098
rect 78024 7046 78076 7098
rect 49884 6808 49936 6860
rect 53196 6808 53248 6860
rect 26424 6783 26476 6792
rect 26424 6749 26433 6783
rect 26433 6749 26467 6783
rect 26467 6749 26476 6783
rect 26424 6740 26476 6749
rect 31392 6672 31444 6724
rect 39120 6740 39172 6792
rect 56968 6740 57020 6792
rect 39948 6672 40000 6724
rect 20720 6604 20772 6656
rect 35256 6604 35308 6656
rect 56048 6604 56100 6656
rect 22898 6502 22950 6554
rect 22962 6502 23014 6554
rect 23026 6502 23078 6554
rect 23090 6502 23142 6554
rect 23154 6502 23206 6554
rect 44846 6502 44898 6554
rect 44910 6502 44962 6554
rect 44974 6502 45026 6554
rect 45038 6502 45090 6554
rect 45102 6502 45154 6554
rect 66794 6502 66846 6554
rect 66858 6502 66910 6554
rect 66922 6502 66974 6554
rect 66986 6502 67038 6554
rect 67050 6502 67102 6554
rect 48504 6400 48556 6452
rect 57336 6400 57388 6452
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 55312 6264 55364 6316
rect 56048 6307 56100 6316
rect 56048 6273 56057 6307
rect 56057 6273 56091 6307
rect 56091 6273 56100 6307
rect 56048 6264 56100 6273
rect 87420 6239 87472 6248
rect 87420 6205 87429 6239
rect 87429 6205 87463 6239
rect 87463 6205 87472 6239
rect 87420 6196 87472 6205
rect 87696 6239 87748 6248
rect 87696 6205 87705 6239
rect 87705 6205 87739 6239
rect 87739 6205 87748 6239
rect 87696 6196 87748 6205
rect 31576 6128 31628 6180
rect 34796 6128 34848 6180
rect 63960 6128 64012 6180
rect 11924 5958 11976 6010
rect 11988 5958 12040 6010
rect 12052 5958 12104 6010
rect 12116 5958 12168 6010
rect 12180 5958 12232 6010
rect 33872 5958 33924 6010
rect 33936 5958 33988 6010
rect 34000 5958 34052 6010
rect 34064 5958 34116 6010
rect 34128 5958 34180 6010
rect 55820 5958 55872 6010
rect 55884 5958 55936 6010
rect 55948 5958 56000 6010
rect 56012 5958 56064 6010
rect 56076 5958 56128 6010
rect 77768 5958 77820 6010
rect 77832 5958 77884 6010
rect 77896 5958 77948 6010
rect 77960 5958 78012 6010
rect 78024 5958 78076 6010
rect 56968 5899 57020 5908
rect 20996 5720 21048 5772
rect 1400 5559 1452 5568
rect 1400 5525 1409 5559
rect 1409 5525 1443 5559
rect 1443 5525 1452 5559
rect 1400 5516 1452 5525
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3700 5652 3752 5704
rect 25136 5695 25188 5704
rect 25136 5661 25145 5695
rect 25145 5661 25179 5695
rect 25179 5661 25188 5695
rect 25136 5652 25188 5661
rect 25780 5652 25832 5704
rect 26148 5584 26200 5636
rect 26424 5516 26476 5568
rect 56968 5865 56977 5899
rect 56977 5865 57011 5899
rect 57011 5865 57020 5899
rect 56968 5856 57020 5865
rect 57704 5720 57756 5772
rect 57336 5695 57388 5704
rect 57336 5661 57345 5695
rect 57345 5661 57379 5695
rect 57379 5661 57388 5695
rect 57336 5652 57388 5661
rect 87972 5695 88024 5704
rect 87972 5661 87981 5695
rect 87981 5661 88015 5695
rect 88015 5661 88024 5695
rect 87972 5652 88024 5661
rect 87696 5584 87748 5636
rect 22898 5414 22950 5466
rect 22962 5414 23014 5466
rect 23026 5414 23078 5466
rect 23090 5414 23142 5466
rect 23154 5414 23206 5466
rect 44846 5414 44898 5466
rect 44910 5414 44962 5466
rect 44974 5414 45026 5466
rect 45038 5414 45090 5466
rect 45102 5414 45154 5466
rect 66794 5414 66846 5466
rect 66858 5414 66910 5466
rect 66922 5414 66974 5466
rect 66986 5414 67038 5466
rect 67050 5414 67102 5466
rect 25136 5312 25188 5364
rect 26424 5244 26476 5296
rect 23664 5176 23716 5228
rect 17224 5108 17276 5160
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 29368 5312 29420 5364
rect 29460 5312 29512 5364
rect 30656 5244 30708 5296
rect 44548 5176 44600 5228
rect 26700 4972 26752 5024
rect 70676 4972 70728 5024
rect 71228 4972 71280 5024
rect 88064 5015 88116 5024
rect 88064 4981 88073 5015
rect 88073 4981 88107 5015
rect 88107 4981 88116 5015
rect 88064 4972 88116 4981
rect 11924 4870 11976 4922
rect 11988 4870 12040 4922
rect 12052 4870 12104 4922
rect 12116 4870 12168 4922
rect 12180 4870 12232 4922
rect 33872 4870 33924 4922
rect 33936 4870 33988 4922
rect 34000 4870 34052 4922
rect 34064 4870 34116 4922
rect 34128 4870 34180 4922
rect 55820 4870 55872 4922
rect 55884 4870 55936 4922
rect 55948 4870 56000 4922
rect 56012 4870 56064 4922
rect 56076 4870 56128 4922
rect 77768 4870 77820 4922
rect 77832 4870 77884 4922
rect 77896 4870 77948 4922
rect 77960 4870 78012 4922
rect 78024 4870 78076 4922
rect 31852 4768 31904 4820
rect 41236 4768 41288 4820
rect 50712 4768 50764 4820
rect 51448 4768 51500 4820
rect 63224 4768 63276 4820
rect 83832 4768 83884 4820
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 24768 4632 24820 4684
rect 37924 4700 37976 4752
rect 29368 4632 29420 4684
rect 26148 4607 26200 4616
rect 26148 4573 26157 4607
rect 26157 4573 26191 4607
rect 26191 4573 26200 4607
rect 26148 4564 26200 4573
rect 57336 4564 57388 4616
rect 71136 4564 71188 4616
rect 17224 4496 17276 4548
rect 17960 4428 18012 4480
rect 32956 4496 33008 4548
rect 33600 4539 33652 4548
rect 33600 4505 33609 4539
rect 33609 4505 33643 4539
rect 33643 4505 33652 4539
rect 33600 4496 33652 4505
rect 59452 4496 59504 4548
rect 22652 4428 22704 4480
rect 27528 4471 27580 4480
rect 27528 4437 27537 4471
rect 27537 4437 27571 4471
rect 27571 4437 27580 4471
rect 27528 4428 27580 4437
rect 27712 4428 27764 4480
rect 28908 4428 28960 4480
rect 38844 4428 38896 4480
rect 46296 4428 46348 4480
rect 49240 4428 49292 4480
rect 53104 4428 53156 4480
rect 55680 4471 55732 4480
rect 55680 4437 55689 4471
rect 55689 4437 55723 4471
rect 55723 4437 55732 4471
rect 55680 4428 55732 4437
rect 88064 4471 88116 4480
rect 88064 4437 88073 4471
rect 88073 4437 88107 4471
rect 88107 4437 88116 4471
rect 88064 4428 88116 4437
rect 22898 4326 22950 4378
rect 22962 4326 23014 4378
rect 23026 4326 23078 4378
rect 23090 4326 23142 4378
rect 23154 4326 23206 4378
rect 44846 4326 44898 4378
rect 44910 4326 44962 4378
rect 44974 4326 45026 4378
rect 45038 4326 45090 4378
rect 45102 4326 45154 4378
rect 66794 4326 66846 4378
rect 66858 4326 66910 4378
rect 66922 4326 66974 4378
rect 66986 4326 67038 4378
rect 67050 4326 67102 4378
rect 27528 4224 27580 4276
rect 49424 4267 49476 4276
rect 30656 4156 30708 4208
rect 31208 4156 31260 4208
rect 33600 4156 33652 4208
rect 49424 4233 49433 4267
rect 49433 4233 49467 4267
rect 49467 4233 49476 4267
rect 49424 4224 49476 4233
rect 53104 4224 53156 4276
rect 49240 4156 49292 4208
rect 51448 4156 51500 4208
rect 2780 3952 2832 4004
rect 2964 3884 3016 3936
rect 25412 4088 25464 4140
rect 44364 4088 44416 4140
rect 49976 4088 50028 4140
rect 19156 4020 19208 4072
rect 45376 4020 45428 4072
rect 7104 3952 7156 4004
rect 29000 3952 29052 4004
rect 29184 3952 29236 4004
rect 36544 3952 36596 4004
rect 38108 3952 38160 4004
rect 43444 3952 43496 4004
rect 51448 4020 51500 4072
rect 51816 4156 51868 4208
rect 59452 4156 59504 4208
rect 70676 4156 70728 4208
rect 54024 4088 54076 4140
rect 51908 4020 51960 4072
rect 63592 4088 63644 4140
rect 64052 4088 64104 4140
rect 71136 4063 71188 4072
rect 46480 3952 46532 4004
rect 71136 4029 71145 4063
rect 71145 4029 71179 4063
rect 71179 4029 71188 4063
rect 71136 4020 71188 4029
rect 86868 4088 86920 4140
rect 87696 4131 87748 4140
rect 87696 4097 87705 4131
rect 87705 4097 87739 4131
rect 87739 4097 87748 4131
rect 87696 4088 87748 4097
rect 87880 4088 87932 4140
rect 63868 3952 63920 4004
rect 72608 4020 72660 4072
rect 46296 3884 46348 3936
rect 49700 3884 49752 3936
rect 51632 3884 51684 3936
rect 59636 3927 59688 3936
rect 59636 3893 59645 3927
rect 59645 3893 59679 3927
rect 59679 3893 59688 3927
rect 59636 3884 59688 3893
rect 71596 3884 71648 3936
rect 81532 3952 81584 4004
rect 88248 3952 88300 4004
rect 86868 3884 86920 3936
rect 87880 3884 87932 3936
rect 88064 3927 88116 3936
rect 88064 3893 88073 3927
rect 88073 3893 88107 3927
rect 88107 3893 88116 3927
rect 88064 3884 88116 3893
rect 11924 3782 11976 3834
rect 11988 3782 12040 3834
rect 12052 3782 12104 3834
rect 12116 3782 12168 3834
rect 12180 3782 12232 3834
rect 33872 3782 33924 3834
rect 33936 3782 33988 3834
rect 34000 3782 34052 3834
rect 34064 3782 34116 3834
rect 34128 3782 34180 3834
rect 55820 3782 55872 3834
rect 55884 3782 55936 3834
rect 55948 3782 56000 3834
rect 56012 3782 56064 3834
rect 56076 3782 56128 3834
rect 77768 3782 77820 3834
rect 77832 3782 77884 3834
rect 77896 3782 77948 3834
rect 77960 3782 78012 3834
rect 78024 3782 78076 3834
rect 17224 3680 17276 3732
rect 27896 3680 27948 3732
rect 29184 3680 29236 3732
rect 30840 3723 30892 3732
rect 30840 3689 30849 3723
rect 30849 3689 30883 3723
rect 30883 3689 30892 3723
rect 30840 3680 30892 3689
rect 31392 3680 31444 3732
rect 31484 3680 31536 3732
rect 34704 3680 34756 3732
rect 34888 3680 34940 3732
rect 42616 3680 42668 3732
rect 42708 3680 42760 3732
rect 46296 3680 46348 3732
rect 47860 3680 47912 3732
rect 664 3612 716 3664
rect 9956 3612 10008 3664
rect 11704 3544 11756 3596
rect 22744 3612 22796 3664
rect 41880 3612 41932 3664
rect 3516 3476 3568 3528
rect 9312 3476 9364 3528
rect 18236 3476 18288 3528
rect 24400 3519 24452 3528
rect 24400 3485 24409 3519
rect 24409 3485 24443 3519
rect 24443 3485 24452 3519
rect 24400 3476 24452 3485
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 24952 3476 25004 3528
rect 26700 3519 26752 3528
rect 26700 3485 26709 3519
rect 26709 3485 26743 3519
rect 26743 3485 26752 3519
rect 26700 3476 26752 3485
rect 4988 3408 5040 3460
rect 1400 3383 1452 3392
rect 1400 3349 1409 3383
rect 1409 3349 1443 3383
rect 1443 3349 1452 3383
rect 1400 3340 1452 3349
rect 1492 3340 1544 3392
rect 13820 3408 13872 3460
rect 20720 3408 20772 3460
rect 21180 3340 21232 3392
rect 24768 3383 24820 3392
rect 24768 3349 24777 3383
rect 24777 3349 24811 3383
rect 24811 3349 24820 3383
rect 24768 3340 24820 3349
rect 25780 3340 25832 3392
rect 26608 3340 26660 3392
rect 28540 3476 28592 3528
rect 30748 3476 30800 3528
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 31392 3519 31444 3528
rect 31392 3485 31401 3519
rect 31401 3485 31435 3519
rect 31435 3485 31444 3519
rect 31392 3476 31444 3485
rect 33048 3519 33100 3528
rect 33048 3485 33057 3519
rect 33057 3485 33091 3519
rect 33091 3485 33100 3519
rect 33048 3476 33100 3485
rect 33508 3544 33560 3596
rect 35532 3544 35584 3596
rect 38108 3544 38160 3596
rect 39304 3544 39356 3596
rect 41420 3544 41472 3596
rect 42708 3544 42760 3596
rect 45376 3544 45428 3596
rect 47492 3544 47544 3596
rect 49608 3680 49660 3732
rect 49700 3680 49752 3732
rect 48228 3612 48280 3664
rect 51356 3612 51408 3664
rect 64144 3680 64196 3732
rect 87788 3680 87840 3732
rect 87880 3680 87932 3732
rect 89536 3680 89588 3732
rect 76748 3612 76800 3664
rect 86684 3612 86736 3664
rect 87604 3612 87656 3664
rect 48136 3544 48188 3596
rect 27712 3340 27764 3392
rect 27896 3340 27948 3392
rect 30012 3408 30064 3460
rect 30288 3408 30340 3460
rect 31300 3408 31352 3460
rect 33968 3408 34020 3460
rect 36544 3476 36596 3528
rect 43444 3476 43496 3528
rect 46020 3476 46072 3528
rect 48872 3476 48924 3528
rect 48964 3476 49016 3528
rect 37280 3408 37332 3460
rect 41236 3408 41288 3460
rect 48688 3408 48740 3460
rect 28724 3340 28776 3392
rect 31484 3340 31536 3392
rect 31668 3340 31720 3392
rect 32588 3340 32640 3392
rect 33048 3340 33100 3392
rect 39396 3340 39448 3392
rect 41880 3340 41932 3392
rect 45192 3340 45244 3392
rect 47124 3383 47176 3392
rect 47124 3349 47133 3383
rect 47133 3349 47167 3383
rect 47167 3349 47176 3383
rect 47124 3340 47176 3349
rect 47492 3383 47544 3392
rect 47492 3349 47501 3383
rect 47501 3349 47535 3383
rect 47535 3349 47544 3383
rect 47492 3340 47544 3349
rect 49240 3340 49292 3392
rect 49700 3544 49752 3596
rect 50160 3544 50212 3596
rect 52552 3544 52604 3596
rect 58348 3544 58400 3596
rect 58624 3544 58676 3596
rect 73528 3544 73580 3596
rect 50252 3476 50304 3528
rect 50528 3519 50580 3528
rect 50528 3485 50537 3519
rect 50537 3485 50571 3519
rect 50571 3485 50580 3519
rect 50528 3476 50580 3485
rect 51356 3476 51408 3528
rect 62396 3476 62448 3528
rect 70216 3476 70268 3528
rect 75184 3476 75236 3528
rect 86592 3519 86644 3528
rect 86592 3485 86601 3519
rect 86601 3485 86635 3519
rect 86635 3485 86644 3519
rect 86592 3476 86644 3485
rect 88156 3476 88208 3528
rect 49516 3408 49568 3460
rect 51448 3408 51500 3460
rect 52920 3383 52972 3392
rect 52920 3349 52929 3383
rect 52929 3349 52963 3383
rect 52963 3349 52972 3383
rect 53196 3408 53248 3460
rect 52920 3340 52972 3349
rect 22898 3238 22950 3290
rect 22962 3238 23014 3290
rect 23026 3238 23078 3290
rect 23090 3238 23142 3290
rect 23154 3238 23206 3290
rect 44846 3238 44898 3290
rect 44910 3238 44962 3290
rect 44974 3238 45026 3290
rect 45038 3238 45090 3290
rect 45102 3238 45154 3290
rect 66794 3238 66846 3290
rect 66858 3238 66910 3290
rect 66922 3238 66974 3290
rect 66986 3238 67038 3290
rect 67050 3238 67102 3290
rect 1676 3136 1728 3188
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 20 3000 72 3052
rect 16580 3136 16632 3188
rect 4528 3068 4580 3120
rect 9312 3068 9364 3120
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 4804 3043 4856 3052
rect 3700 3000 3752 3009
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 7104 3043 7156 3052
rect 7104 3009 7113 3043
rect 7113 3009 7147 3043
rect 7147 3009 7156 3043
rect 7104 3000 7156 3009
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 4528 2864 4580 2916
rect 9956 2864 10008 2916
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 16764 3000 16816 3052
rect 24216 3136 24268 3188
rect 46020 3136 46072 3188
rect 26148 3068 26200 3120
rect 17224 2864 17276 2916
rect 1952 2796 2004 2848
rect 4896 2796 4948 2848
rect 5540 2839 5592 2848
rect 5540 2805 5549 2839
rect 5549 2805 5583 2839
rect 5583 2805 5592 2839
rect 5540 2796 5592 2805
rect 6460 2796 6512 2848
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 10232 2796 10284 2848
rect 13544 2796 13596 2848
rect 17960 2864 18012 2916
rect 22744 3000 22796 3052
rect 24768 3000 24820 3052
rect 25412 3043 25464 3052
rect 25412 3009 25421 3043
rect 25421 3009 25455 3043
rect 25455 3009 25464 3043
rect 25412 3000 25464 3009
rect 25964 3043 26016 3052
rect 25964 3009 25973 3043
rect 25973 3009 26007 3043
rect 26007 3009 26016 3043
rect 25964 3000 26016 3009
rect 26332 3043 26384 3052
rect 26332 3009 26341 3043
rect 26341 3009 26375 3043
rect 26375 3009 26384 3043
rect 26332 3000 26384 3009
rect 27712 3000 27764 3052
rect 31760 3068 31812 3120
rect 33968 3111 34020 3120
rect 24216 2932 24268 2984
rect 26240 2932 26292 2984
rect 24400 2864 24452 2916
rect 17408 2796 17460 2848
rect 19984 2796 20036 2848
rect 22836 2839 22888 2848
rect 22836 2805 22845 2839
rect 22845 2805 22879 2839
rect 22879 2805 22888 2839
rect 22836 2796 22888 2805
rect 25136 2796 25188 2848
rect 25412 2796 25464 2848
rect 29184 2907 29236 2916
rect 29184 2873 29193 2907
rect 29193 2873 29227 2907
rect 29227 2873 29236 2907
rect 31668 3043 31720 3052
rect 31668 3009 31677 3043
rect 31677 3009 31711 3043
rect 31711 3009 31720 3043
rect 31668 3000 31720 3009
rect 33968 3077 33977 3111
rect 33977 3077 34011 3111
rect 34011 3077 34020 3111
rect 33968 3068 34020 3077
rect 34704 3068 34756 3120
rect 39120 3068 39172 3120
rect 32588 3043 32640 3052
rect 32588 3009 32597 3043
rect 32597 3009 32631 3043
rect 32631 3009 32640 3043
rect 32588 3000 32640 3009
rect 34888 3000 34940 3052
rect 38936 3000 38988 3052
rect 39304 3043 39356 3052
rect 39304 3009 39313 3043
rect 39313 3009 39347 3043
rect 39347 3009 39356 3043
rect 39304 3000 39356 3009
rect 40224 3043 40276 3052
rect 40224 3009 40233 3043
rect 40233 3009 40267 3043
rect 40267 3009 40276 3043
rect 40224 3000 40276 3009
rect 41604 3068 41656 3120
rect 43260 3068 43312 3120
rect 43904 3000 43956 3052
rect 47124 3043 47176 3052
rect 47124 3009 47133 3043
rect 47133 3009 47167 3043
rect 47167 3009 47176 3043
rect 47124 3000 47176 3009
rect 29184 2864 29236 2873
rect 33508 2864 33560 2916
rect 39396 2932 39448 2984
rect 46296 2932 46348 2984
rect 46388 2932 46440 2984
rect 50344 3136 50396 3188
rect 52000 3179 52052 3188
rect 49424 3068 49476 3120
rect 52000 3145 52009 3179
rect 52009 3145 52043 3179
rect 52043 3145 52052 3179
rect 52000 3136 52052 3145
rect 52184 3136 52236 3188
rect 59636 3136 59688 3188
rect 49608 3043 49660 3052
rect 49608 3009 49617 3043
rect 49617 3009 49651 3043
rect 49651 3009 49660 3043
rect 49608 3000 49660 3009
rect 50252 3000 50304 3052
rect 51632 3043 51684 3052
rect 51632 3009 51641 3043
rect 51641 3009 51675 3043
rect 51675 3009 51684 3043
rect 51632 3000 51684 3009
rect 41604 2864 41656 2916
rect 43444 2864 43496 2916
rect 29460 2796 29512 2848
rect 30380 2839 30432 2848
rect 30380 2805 30389 2839
rect 30389 2805 30423 2839
rect 30423 2805 30432 2839
rect 30380 2796 30432 2805
rect 31484 2839 31536 2848
rect 31484 2805 31493 2839
rect 31493 2805 31527 2839
rect 31527 2805 31536 2839
rect 31484 2796 31536 2805
rect 35716 2796 35768 2848
rect 37464 2796 37516 2848
rect 39764 2796 39816 2848
rect 39948 2796 40000 2848
rect 42800 2796 42852 2848
rect 43260 2796 43312 2848
rect 47492 2796 47544 2848
rect 51448 2907 51500 2916
rect 51448 2873 51457 2907
rect 51457 2873 51491 2907
rect 51491 2873 51500 2907
rect 51448 2864 51500 2873
rect 51724 2932 51776 2984
rect 53656 3000 53708 3052
rect 55680 3000 55732 3052
rect 58624 3043 58676 3052
rect 51908 2864 51960 2916
rect 52184 2864 52236 2916
rect 54944 2932 54996 2984
rect 58624 3009 58633 3043
rect 58633 3009 58667 3043
rect 58667 3009 58676 3043
rect 58624 3000 58676 3009
rect 63500 3136 63552 3188
rect 63132 3000 63184 3052
rect 75184 3136 75236 3188
rect 76748 3111 76800 3120
rect 71596 3043 71648 3052
rect 54392 2796 54444 2848
rect 56600 2796 56652 2848
rect 58348 2796 58400 2848
rect 59176 2796 59228 2848
rect 62488 2796 62540 2848
rect 64420 2932 64472 2984
rect 71596 3009 71605 3043
rect 71605 3009 71639 3043
rect 71639 3009 71648 3043
rect 71596 3000 71648 3009
rect 76748 3077 76757 3111
rect 76757 3077 76791 3111
rect 76791 3077 76800 3111
rect 76748 3068 76800 3077
rect 77116 3111 77168 3120
rect 77116 3077 77125 3111
rect 77125 3077 77159 3111
rect 77159 3077 77168 3111
rect 77116 3068 77168 3077
rect 79692 3068 79744 3120
rect 76748 2932 76800 2984
rect 81532 3043 81584 3052
rect 81532 3009 81541 3043
rect 81541 3009 81575 3043
rect 81575 3009 81584 3043
rect 81532 3000 81584 3009
rect 87696 3136 87748 3188
rect 87788 3136 87840 3188
rect 88340 3179 88392 3188
rect 88340 3145 88349 3179
rect 88349 3145 88383 3179
rect 88383 3145 88392 3179
rect 88340 3136 88392 3145
rect 85028 2932 85080 2984
rect 85120 2932 85172 2984
rect 86868 2932 86920 2984
rect 85488 2864 85540 2916
rect 67456 2796 67508 2848
rect 68376 2796 68428 2848
rect 71504 2796 71556 2848
rect 79968 2796 80020 2848
rect 81808 2796 81860 2848
rect 86960 2796 87012 2848
rect 11924 2694 11976 2746
rect 11988 2694 12040 2746
rect 12052 2694 12104 2746
rect 12116 2694 12168 2746
rect 12180 2694 12232 2746
rect 33872 2694 33924 2746
rect 33936 2694 33988 2746
rect 34000 2694 34052 2746
rect 34064 2694 34116 2746
rect 34128 2694 34180 2746
rect 55820 2694 55872 2746
rect 55884 2694 55936 2746
rect 55948 2694 56000 2746
rect 56012 2694 56064 2746
rect 56076 2694 56128 2746
rect 77768 2694 77820 2746
rect 77832 2694 77884 2746
rect 77896 2694 77948 2746
rect 77960 2694 78012 2746
rect 78024 2694 78076 2746
rect 4160 2524 4212 2576
rect 21180 2524 21232 2576
rect 23296 2524 23348 2576
rect 26424 2524 26476 2576
rect 26516 2524 26568 2576
rect 27252 2524 27304 2576
rect 27528 2524 27580 2576
rect 2872 2388 2924 2440
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5540 2388 5592 2440
rect 5816 2388 5868 2440
rect 7748 2388 7800 2440
rect 10232 2456 10284 2508
rect 15844 2456 15896 2508
rect 18696 2456 18748 2508
rect 9772 2388 9824 2440
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10508 2431 10560 2440
rect 10508 2397 10517 2431
rect 10517 2397 10551 2431
rect 10551 2397 10560 2431
rect 10508 2388 10560 2397
rect 1308 2320 1360 2372
rect 2688 2320 2740 2372
rect 3884 2320 3936 2372
rect 11612 2363 11664 2372
rect 11612 2329 11621 2363
rect 11621 2329 11655 2363
rect 11655 2329 11664 2363
rect 11612 2320 11664 2329
rect 12256 2388 12308 2440
rect 12900 2388 12952 2440
rect 14188 2388 14240 2440
rect 14372 2431 14424 2440
rect 14372 2397 14381 2431
rect 14381 2397 14415 2431
rect 14415 2397 14424 2431
rect 14372 2388 14424 2397
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16120 2388 16172 2440
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 18052 2388 18104 2440
rect 20168 2456 20220 2508
rect 20812 2431 20864 2440
rect 15384 2320 15436 2372
rect 20812 2397 20821 2431
rect 20821 2397 20855 2431
rect 20855 2397 20864 2431
rect 20812 2388 20864 2397
rect 22836 2456 22888 2508
rect 21916 2388 21968 2440
rect 23940 2431 23992 2440
rect 23940 2397 23949 2431
rect 23949 2397 23983 2431
rect 23983 2397 23992 2431
rect 23940 2388 23992 2397
rect 24216 2431 24268 2440
rect 24216 2397 24225 2431
rect 24225 2397 24259 2431
rect 24259 2397 24268 2431
rect 24216 2388 24268 2397
rect 24768 2431 24820 2440
rect 24768 2397 24777 2431
rect 24777 2397 24811 2431
rect 24811 2397 24820 2431
rect 24768 2388 24820 2397
rect 25412 2431 25464 2440
rect 25412 2397 25421 2431
rect 25421 2397 25455 2431
rect 25455 2397 25464 2431
rect 25412 2388 25464 2397
rect 26516 2431 26568 2440
rect 26516 2397 26525 2431
rect 26525 2397 26559 2431
rect 26559 2397 26568 2431
rect 26516 2388 26568 2397
rect 27620 2456 27672 2508
rect 27804 2592 27856 2644
rect 29920 2592 29972 2644
rect 30380 2592 30432 2644
rect 31116 2592 31168 2644
rect 45468 2592 45520 2644
rect 46296 2592 46348 2644
rect 49976 2592 50028 2644
rect 50252 2592 50304 2644
rect 53288 2592 53340 2644
rect 55588 2592 55640 2644
rect 59268 2592 59320 2644
rect 61292 2635 61344 2644
rect 61292 2601 61301 2635
rect 61301 2601 61335 2635
rect 61335 2601 61344 2635
rect 61292 2592 61344 2601
rect 63684 2592 63736 2644
rect 69020 2635 69072 2644
rect 31668 2524 31720 2576
rect 31852 2524 31904 2576
rect 27896 2388 27948 2440
rect 31576 2456 31628 2508
rect 34888 2524 34940 2576
rect 38752 2524 38804 2576
rect 38936 2524 38988 2576
rect 29920 2431 29972 2440
rect 29920 2397 29929 2431
rect 29929 2397 29963 2431
rect 29963 2397 29972 2431
rect 29920 2388 29972 2397
rect 26148 2320 26200 2372
rect 2596 2295 2648 2304
rect 2596 2261 2605 2295
rect 2605 2261 2639 2295
rect 2639 2261 2648 2295
rect 2596 2252 2648 2261
rect 3240 2252 3292 2304
rect 4252 2295 4304 2304
rect 4252 2261 4261 2295
rect 4261 2261 4295 2295
rect 4295 2261 4304 2295
rect 4252 2252 4304 2261
rect 5172 2252 5224 2304
rect 8208 2252 8260 2304
rect 8392 2252 8444 2304
rect 9036 2252 9088 2304
rect 9680 2252 9732 2304
rect 10324 2295 10376 2304
rect 10324 2261 10333 2295
rect 10333 2261 10367 2295
rect 10367 2261 10376 2295
rect 10324 2252 10376 2261
rect 10968 2252 11020 2304
rect 12348 2295 12400 2304
rect 12348 2261 12357 2295
rect 12357 2261 12391 2295
rect 12391 2261 12400 2295
rect 12348 2252 12400 2261
rect 15476 2252 15528 2304
rect 19340 2252 19392 2304
rect 20628 2295 20680 2304
rect 20628 2261 20637 2295
rect 20637 2261 20671 2295
rect 20671 2261 20680 2295
rect 20628 2252 20680 2261
rect 21272 2252 21324 2304
rect 22192 2295 22244 2304
rect 22192 2261 22201 2295
rect 22201 2261 22235 2295
rect 22235 2261 22244 2295
rect 22192 2252 22244 2261
rect 23848 2252 23900 2304
rect 24032 2252 24084 2304
rect 24400 2252 24452 2304
rect 24492 2252 24544 2304
rect 26976 2320 27028 2372
rect 27804 2320 27856 2372
rect 29000 2320 29052 2372
rect 31484 2388 31536 2440
rect 32864 2388 32916 2440
rect 34796 2388 34848 2440
rect 35348 2388 35400 2440
rect 35440 2388 35492 2440
rect 36360 2456 36412 2508
rect 36820 2431 36872 2440
rect 36820 2397 36829 2431
rect 36829 2397 36863 2431
rect 36863 2397 36872 2431
rect 36820 2388 36872 2397
rect 37648 2431 37700 2440
rect 37648 2397 37657 2431
rect 37657 2397 37691 2431
rect 37691 2397 37700 2431
rect 37648 2388 37700 2397
rect 39764 2456 39816 2508
rect 38752 2388 38804 2440
rect 39304 2388 39356 2440
rect 40500 2456 40552 2508
rect 43720 2524 43772 2576
rect 45284 2524 45336 2576
rect 41972 2431 42024 2440
rect 41972 2397 41981 2431
rect 41981 2397 42015 2431
rect 42015 2397 42024 2431
rect 41972 2388 42024 2397
rect 42800 2431 42852 2440
rect 42800 2397 42809 2431
rect 42809 2397 42843 2431
rect 42843 2397 42852 2431
rect 42800 2388 42852 2397
rect 43444 2431 43496 2440
rect 43444 2397 43453 2431
rect 43453 2397 43487 2431
rect 43487 2397 43496 2431
rect 43444 2388 43496 2397
rect 27068 2252 27120 2304
rect 28264 2295 28316 2304
rect 28264 2261 28273 2295
rect 28273 2261 28307 2295
rect 28307 2261 28316 2295
rect 28264 2252 28316 2261
rect 29184 2252 29236 2304
rect 29644 2252 29696 2304
rect 31116 2320 31168 2372
rect 31300 2320 31352 2372
rect 32680 2320 32732 2372
rect 32220 2252 32272 2304
rect 34060 2252 34112 2304
rect 34152 2252 34204 2304
rect 36084 2295 36136 2304
rect 36084 2261 36093 2295
rect 36093 2261 36127 2295
rect 36127 2261 36136 2295
rect 36084 2252 36136 2261
rect 36728 2252 36780 2304
rect 37372 2252 37424 2304
rect 39120 2320 39172 2372
rect 41696 2320 41748 2372
rect 46848 2456 46900 2508
rect 50712 2499 50764 2508
rect 44456 2388 44508 2440
rect 45192 2388 45244 2440
rect 46388 2388 46440 2440
rect 46756 2388 46808 2440
rect 47032 2388 47084 2440
rect 48228 2388 48280 2440
rect 48412 2388 48464 2440
rect 49608 2388 49660 2440
rect 50712 2465 50721 2499
rect 50721 2465 50755 2499
rect 50755 2465 50764 2499
rect 50712 2456 50764 2465
rect 50988 2456 51040 2508
rect 54392 2431 54444 2440
rect 54392 2397 54401 2431
rect 54401 2397 54435 2431
rect 54435 2397 54444 2431
rect 54392 2388 54444 2397
rect 54760 2388 54812 2440
rect 56600 2431 56652 2440
rect 47860 2320 47912 2372
rect 38660 2252 38712 2304
rect 38752 2295 38804 2304
rect 38752 2261 38761 2295
rect 38761 2261 38795 2295
rect 38795 2261 38804 2295
rect 38752 2252 38804 2261
rect 40592 2252 40644 2304
rect 41880 2252 41932 2304
rect 42524 2252 42576 2304
rect 43168 2252 43220 2304
rect 43812 2295 43864 2304
rect 43812 2261 43821 2295
rect 43821 2261 43855 2295
rect 43855 2261 43864 2295
rect 43812 2252 43864 2261
rect 45560 2252 45612 2304
rect 48044 2252 48096 2304
rect 48228 2252 48280 2304
rect 48780 2252 48832 2304
rect 50344 2252 50396 2304
rect 50620 2295 50672 2304
rect 50620 2261 50629 2295
rect 50629 2261 50663 2295
rect 50663 2261 50672 2295
rect 50896 2320 50948 2372
rect 52828 2320 52880 2372
rect 55404 2320 55456 2372
rect 56600 2397 56609 2431
rect 56609 2397 56643 2431
rect 56643 2397 56652 2431
rect 56600 2388 56652 2397
rect 57152 2431 57204 2440
rect 57152 2397 57161 2431
rect 57161 2397 57195 2431
rect 57195 2397 57204 2431
rect 57152 2388 57204 2397
rect 57980 2388 58032 2440
rect 58348 2388 58400 2440
rect 59176 2431 59228 2440
rect 59176 2397 59185 2431
rect 59185 2397 59219 2431
rect 59219 2397 59228 2431
rect 59176 2388 59228 2397
rect 59268 2388 59320 2440
rect 59912 2388 59964 2440
rect 61200 2388 61252 2440
rect 62212 2456 62264 2508
rect 63132 2388 63184 2440
rect 63500 2431 63552 2440
rect 63500 2397 63509 2431
rect 63509 2397 63543 2431
rect 63543 2397 63552 2431
rect 63500 2388 63552 2397
rect 64972 2456 65024 2508
rect 66260 2388 66312 2440
rect 66444 2388 66496 2440
rect 67456 2431 67508 2440
rect 67456 2397 67465 2431
rect 67465 2397 67499 2431
rect 67499 2397 67508 2431
rect 67456 2388 67508 2397
rect 68376 2431 68428 2440
rect 68376 2397 68385 2431
rect 68385 2397 68419 2431
rect 68419 2397 68428 2431
rect 68376 2388 68428 2397
rect 69020 2601 69029 2635
rect 69029 2601 69063 2635
rect 69063 2601 69072 2635
rect 69020 2592 69072 2601
rect 70768 2635 70820 2644
rect 70768 2601 70777 2635
rect 70777 2601 70811 2635
rect 70811 2601 70820 2635
rect 70768 2592 70820 2601
rect 71412 2592 71464 2644
rect 71596 2592 71648 2644
rect 68928 2524 68980 2576
rect 68836 2388 68888 2440
rect 68928 2388 68980 2440
rect 70216 2388 70268 2440
rect 70860 2320 70912 2372
rect 72148 2388 72200 2440
rect 73528 2431 73580 2440
rect 73528 2397 73537 2431
rect 73537 2397 73571 2431
rect 73571 2397 73580 2431
rect 73528 2388 73580 2397
rect 74080 2388 74132 2440
rect 74724 2320 74776 2372
rect 78588 2524 78640 2576
rect 79232 2524 79284 2576
rect 80796 2567 80848 2576
rect 80796 2533 80805 2567
rect 80805 2533 80839 2567
rect 80839 2533 80848 2567
rect 80796 2524 80848 2533
rect 81164 2524 81216 2576
rect 76748 2431 76800 2440
rect 76748 2397 76757 2431
rect 76757 2397 76791 2431
rect 76791 2397 76800 2431
rect 76748 2388 76800 2397
rect 77024 2388 77076 2440
rect 79508 2431 79560 2440
rect 79508 2397 79517 2431
rect 79517 2397 79551 2431
rect 79551 2397 79560 2431
rect 79508 2388 79560 2397
rect 79968 2388 80020 2440
rect 77944 2320 77996 2372
rect 50620 2252 50672 2261
rect 50988 2252 51040 2304
rect 51448 2295 51500 2304
rect 51448 2261 51457 2295
rect 51457 2261 51491 2295
rect 51491 2261 51500 2295
rect 51448 2252 51500 2261
rect 53196 2295 53248 2304
rect 53196 2261 53205 2295
rect 53205 2261 53239 2295
rect 53239 2261 53248 2295
rect 53196 2252 53248 2261
rect 54116 2252 54168 2304
rect 56048 2252 56100 2304
rect 56692 2252 56744 2304
rect 57336 2252 57388 2304
rect 57980 2252 58032 2304
rect 58624 2252 58676 2304
rect 61844 2252 61896 2304
rect 65064 2252 65116 2304
rect 65708 2252 65760 2304
rect 66720 2295 66772 2304
rect 66720 2261 66729 2295
rect 66729 2261 66763 2295
rect 66763 2261 66772 2295
rect 66720 2252 66772 2261
rect 67180 2252 67232 2304
rect 67640 2252 67692 2304
rect 69572 2252 69624 2304
rect 72424 2295 72476 2304
rect 72424 2261 72433 2295
rect 72433 2261 72467 2295
rect 72467 2261 72476 2295
rect 72424 2252 72476 2261
rect 72792 2252 72844 2304
rect 75368 2252 75420 2304
rect 76656 2252 76708 2304
rect 77024 2295 77076 2304
rect 77024 2261 77033 2295
rect 77033 2261 77067 2295
rect 77067 2261 77076 2295
rect 77024 2252 77076 2261
rect 77300 2252 77352 2304
rect 79692 2320 79744 2372
rect 80520 2388 80572 2440
rect 83832 2431 83884 2440
rect 83832 2397 83841 2431
rect 83841 2397 83875 2431
rect 83875 2397 83884 2431
rect 83832 2388 83884 2397
rect 82452 2320 82504 2372
rect 85028 2388 85080 2440
rect 86316 2524 86368 2576
rect 85488 2456 85540 2508
rect 88892 2320 88944 2372
rect 80060 2252 80112 2304
rect 81440 2295 81492 2304
rect 81440 2261 81449 2295
rect 81449 2261 81483 2295
rect 81483 2261 81492 2295
rect 81440 2252 81492 2261
rect 82728 2295 82780 2304
rect 82728 2261 82737 2295
rect 82737 2261 82771 2295
rect 82771 2261 82780 2295
rect 82728 2252 82780 2261
rect 83096 2252 83148 2304
rect 84200 2295 84252 2304
rect 84200 2261 84209 2295
rect 84209 2261 84243 2295
rect 84243 2261 84252 2295
rect 84200 2252 84252 2261
rect 84384 2252 84436 2304
rect 85304 2295 85356 2304
rect 85304 2261 85313 2295
rect 85313 2261 85347 2295
rect 85347 2261 85356 2295
rect 85304 2252 85356 2261
rect 85672 2252 85724 2304
rect 87052 2252 87104 2304
rect 87972 2295 88024 2304
rect 87972 2261 87981 2295
rect 87981 2261 88015 2295
rect 88015 2261 88024 2295
rect 87972 2252 88024 2261
rect 22898 2150 22950 2202
rect 22962 2150 23014 2202
rect 23026 2150 23078 2202
rect 23090 2150 23142 2202
rect 23154 2150 23206 2202
rect 44846 2150 44898 2202
rect 44910 2150 44962 2202
rect 44974 2150 45026 2202
rect 45038 2150 45090 2202
rect 45102 2150 45154 2202
rect 66794 2150 66846 2202
rect 66858 2150 66910 2202
rect 66922 2150 66974 2202
rect 66986 2150 67038 2202
rect 67050 2150 67102 2202
rect 24768 2048 24820 2100
rect 28816 2048 28868 2100
rect 28908 2048 28960 2100
rect 62028 2048 62080 2100
rect 64696 2048 64748 2100
rect 82728 2048 82780 2100
rect 15752 1980 15804 2032
rect 45560 1980 45612 2032
rect 45652 1980 45704 2032
rect 48780 1980 48832 2032
rect 48872 1980 48924 2032
rect 50436 1980 50488 2032
rect 50620 1980 50672 2032
rect 51632 1980 51684 2032
rect 52920 1980 52972 2032
rect 81440 1980 81492 2032
rect 8208 1912 8260 1964
rect 22192 1912 22244 1964
rect 28908 1912 28960 1964
rect 2872 1776 2924 1828
rect 27804 1844 27856 1896
rect 10508 1708 10560 1760
rect 24216 1708 24268 1760
rect 24400 1776 24452 1828
rect 26332 1776 26384 1828
rect 26516 1776 26568 1828
rect 26608 1708 26660 1760
rect 26976 1776 27028 1828
rect 27712 1776 27764 1828
rect 59360 1912 59412 1964
rect 63408 1912 63460 1964
rect 66720 1912 66772 1964
rect 31668 1844 31720 1896
rect 53196 1844 53248 1896
rect 58992 1844 59044 1896
rect 62304 1844 62356 1896
rect 64144 1844 64196 1896
rect 76748 1844 76800 1896
rect 31392 1776 31444 1828
rect 84200 1776 84252 1828
rect 28632 1708 28684 1760
rect 87972 1708 88024 1760
rect 12348 1640 12400 1692
rect 45560 1640 45612 1692
rect 45836 1640 45888 1692
rect 79508 1640 79560 1692
rect 16948 1572 17000 1624
rect 45376 1572 45428 1624
rect 47124 1572 47176 1624
rect 85304 1572 85356 1624
rect 4252 1504 4304 1556
rect 26056 1504 26108 1556
rect 26148 1504 26200 1556
rect 30196 1504 30248 1556
rect 30288 1504 30340 1556
rect 31760 1504 31812 1556
rect 31852 1504 31904 1556
rect 72424 1504 72476 1556
rect 22008 1436 22060 1488
rect 51448 1436 51500 1488
rect 14372 1368 14424 1420
rect 23572 1368 23624 1420
rect 23940 1368 23992 1420
rect 30288 1368 30340 1420
rect 26056 1300 26108 1352
rect 29092 1300 29144 1352
rect 25872 1232 25924 1284
rect 45560 1368 45612 1420
rect 45744 1368 45796 1420
rect 45376 1300 45428 1352
rect 38660 1232 38712 1284
rect 39120 1232 39172 1284
rect 39212 1232 39264 1284
rect 47124 1368 47176 1420
rect 46756 1300 46808 1352
rect 50804 1368 50856 1420
rect 62212 1436 62264 1488
rect 62304 1436 62356 1488
rect 71596 1436 71648 1488
rect 49424 1300 49476 1352
rect 51632 1368 51684 1420
rect 63500 1368 63552 1420
rect 64052 1368 64104 1420
rect 77024 1436 77076 1488
rect 27620 1164 27672 1216
rect 28356 1164 28408 1216
<< metal2 >>
rect 18 29200 74 30000
rect 662 29200 718 30000
rect 1306 29200 1362 30000
rect 2594 29322 2650 30000
rect 2594 29294 2728 29322
rect 2594 29200 2650 29294
rect 32 27130 60 29200
rect 20 27124 72 27130
rect 20 27066 72 27072
rect 676 25770 704 29200
rect 1320 27470 1348 29200
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 1490 27976 1546 27985
rect 1490 27911 1546 27920
rect 1308 27464 1360 27470
rect 1308 27406 1360 27412
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 25945 1440 26318
rect 1504 26042 1532 27911
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1688 26625 1716 27270
rect 1780 27062 1808 28591
rect 2700 27606 2728 29294
rect 2778 29200 2834 29209
rect 3238 29200 3294 30000
rect 3882 29322 3938 30000
rect 4526 29322 4582 30000
rect 5170 29322 5226 30000
rect 3882 29294 4016 29322
rect 3882 29200 3938 29294
rect 2778 29135 2834 29144
rect 2688 27600 2740 27606
rect 2688 27542 2740 27548
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 1768 27056 1820 27062
rect 1768 26998 1820 27004
rect 2044 26852 2096 26858
rect 2044 26794 2096 26800
rect 1674 26616 1730 26625
rect 1674 26551 1730 26560
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1492 26036 1544 26042
rect 1492 25978 1544 25984
rect 1398 25936 1454 25945
rect 1398 25871 1454 25880
rect 664 25764 716 25770
rect 664 25706 716 25712
rect 1400 25288 1452 25294
rect 1398 25256 1400 25265
rect 1452 25256 1454 25265
rect 1398 25191 1454 25200
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1412 24585 1440 24686
rect 1398 24576 1454 24585
rect 1398 24511 1454 24520
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1780 23225 1808 23666
rect 1766 23216 1822 23225
rect 1766 23151 1822 23160
rect 1584 22568 1636 22574
rect 1582 22536 1584 22545
rect 1636 22536 1638 22545
rect 1582 22471 1638 22480
rect 1400 21888 1452 21894
rect 1398 21856 1400 21865
rect 1452 21856 1454 21865
rect 1398 21791 1454 21800
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21185 1440 21490
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1398 21176 1454 21185
rect 1596 21146 1624 21286
rect 1398 21111 1454 21120
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1400 20800 1452 20806
rect 1400 20742 1452 20748
rect 1412 20505 1440 20742
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 1400 19848 1452 19854
rect 1398 19816 1400 19825
rect 1676 19848 1728 19854
rect 1452 19816 1454 19825
rect 1676 19790 1728 19796
rect 1398 19751 1454 19760
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 1412 18465 1440 18566
rect 1398 18456 1454 18465
rect 1398 18391 1454 18400
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 17785 1440 18022
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1400 16448 1452 16454
rect 1398 16416 1400 16425
rect 1452 16416 1454 16425
rect 1398 16351 1454 16360
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 15065 1624 15302
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1582 15056 1638 15065
rect 1582 14991 1638 15000
rect 1584 14408 1636 14414
rect 1582 14376 1584 14385
rect 1636 14376 1638 14385
rect 1582 14311 1638 14320
rect 1400 13728 1452 13734
rect 1398 13696 1400 13705
rect 1452 13696 1454 13705
rect 1398 13631 1454 13640
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 13025 1624 13262
rect 1582 13016 1638 13025
rect 1582 12951 1638 12960
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 12345 1440 12718
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1688 12102 1716 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1780 19145 1808 19314
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1872 18358 1900 26318
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1860 18352 1912 18358
rect 1860 18294 1912 18300
rect 1964 17882 1992 20742
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 2056 17746 2084 26794
rect 2240 26586 2268 27406
rect 2228 26580 2280 26586
rect 2228 26522 2280 26528
rect 2792 26042 2820 29135
rect 3252 27470 3280 29200
rect 3148 27464 3200 27470
rect 3148 27406 3200 27412
rect 3240 27464 3292 27470
rect 3240 27406 3292 27412
rect 3054 27296 3110 27305
rect 3054 27231 3110 27240
rect 3068 27130 3096 27231
rect 3056 27124 3108 27130
rect 3056 27066 3108 27072
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2780 26036 2832 26042
rect 2780 25978 2832 25984
rect 2596 25900 2648 25906
rect 2596 25842 2648 25848
rect 2688 25900 2740 25906
rect 2688 25842 2740 25848
rect 2608 21418 2636 25842
rect 2596 21412 2648 21418
rect 2596 21354 2648 21360
rect 2596 19236 2648 19242
rect 2596 19178 2648 19184
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1780 17105 1808 17138
rect 1766 17096 1822 17105
rect 1766 17031 1822 17040
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 2608 11694 2636 19178
rect 2700 17678 2728 25842
rect 2884 17814 2912 26930
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 2872 17808 2924 17814
rect 2872 17750 2924 17756
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2976 16250 3004 16526
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2596 11688 2648 11694
rect 1398 11656 1454 11665
rect 2596 11630 2648 11636
rect 1398 11591 1400 11600
rect 1452 11591 1454 11600
rect 1400 11562 1452 11568
rect 1400 11008 1452 11014
rect 1398 10976 1400 10985
rect 1452 10976 1454 10985
rect 1398 10911 1454 10920
rect 1582 10704 1638 10713
rect 1582 10639 1584 10648
rect 1636 10639 1638 10648
rect 1584 10610 1636 10616
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 10305 1440 10406
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 9625 1440 9862
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1584 8968 1636 8974
rect 1582 8936 1584 8945
rect 1636 8936 1638 8945
rect 1582 8871 1638 8880
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 6905 1440 7142
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 1400 5568 1452 5574
rect 1398 5536 1400 5545
rect 1452 5536 1454 5545
rect 1398 5471 1454 5480
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1596 4185 1624 4558
rect 1582 4176 1638 4185
rect 1582 4111 1638 4120
rect 664 3664 716 3670
rect 664 3606 716 3612
rect 20 3052 72 3058
rect 20 2994 72 3000
rect 32 800 60 2994
rect 676 800 704 3606
rect 1398 3496 1454 3505
rect 1398 3431 1454 3440
rect 1412 3398 1440 3431
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1504 2825 1532 3334
rect 1688 3194 1716 7686
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1780 6225 1808 6258
rect 1766 6216 1822 6225
rect 1766 6151 1822 6160
rect 3068 5710 3096 26318
rect 3160 25702 3188 27406
rect 3988 27130 4016 29294
rect 4526 29294 4752 29322
rect 4526 29200 4582 29294
rect 4724 27470 4752 29294
rect 5170 29294 5304 29322
rect 5170 29200 5226 29294
rect 5276 27606 5304 29294
rect 5814 29200 5870 30000
rect 6458 29322 6514 30000
rect 7102 29322 7158 30000
rect 6458 29294 6776 29322
rect 6458 29200 6514 29294
rect 5264 27600 5316 27606
rect 5264 27542 5316 27548
rect 5828 27538 5856 29200
rect 5816 27532 5868 27538
rect 5816 27474 5868 27480
rect 4712 27464 4764 27470
rect 4712 27406 4764 27412
rect 6644 27464 6696 27470
rect 6644 27406 6696 27412
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4804 27328 4856 27334
rect 4804 27270 4856 27276
rect 3976 27124 4028 27130
rect 3976 27066 4028 27072
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 3792 26240 3844 26246
rect 3792 26182 3844 26188
rect 3804 25906 3832 26182
rect 3792 25900 3844 25906
rect 3792 25842 3844 25848
rect 3148 25696 3200 25702
rect 3148 25638 3200 25644
rect 3988 21690 4016 26318
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3988 12782 4016 21490
rect 4080 17610 4108 27270
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4172 19174 4200 26930
rect 4816 22982 4844 27270
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1952 2848 2004 2854
rect 1490 2816 1546 2825
rect 1952 2790 2004 2796
rect 1490 2751 1546 2760
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 800 1348 2314
rect 1964 800 1992 2790
rect 2686 2408 2742 2417
rect 2686 2343 2688 2352
rect 2740 2343 2742 2352
rect 2688 2314 2740 2320
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 800 2636 2246
rect 2792 1465 2820 3946
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2884 1834 2912 2382
rect 2976 2145 3004 3878
rect 3344 2446 3372 12718
rect 4816 11354 4844 21422
rect 6656 14550 6684 27406
rect 6748 27062 6776 29294
rect 7102 29294 7328 29322
rect 7102 29200 7158 29294
rect 7300 27130 7328 29294
rect 7746 29200 7802 30000
rect 8390 29322 8446 30000
rect 9034 29322 9090 30000
rect 10322 29322 10378 30000
rect 8390 29294 8524 29322
rect 8390 29200 8446 29294
rect 7760 27606 7788 29200
rect 8496 27606 8524 29294
rect 9034 29294 9168 29322
rect 9034 29200 9090 29294
rect 9140 27606 9168 29294
rect 10322 29294 10456 29322
rect 10322 29200 10378 29294
rect 7748 27600 7800 27606
rect 7748 27542 7800 27548
rect 8484 27600 8536 27606
rect 8484 27542 8536 27548
rect 9128 27600 9180 27606
rect 9128 27542 9180 27548
rect 9220 27600 9272 27606
rect 9220 27542 9272 27548
rect 9232 27470 9260 27542
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9692 27334 9720 27406
rect 9680 27328 9732 27334
rect 9680 27270 9732 27276
rect 7288 27124 7340 27130
rect 7288 27066 7340 27072
rect 6736 27056 6788 27062
rect 6736 26998 6788 27004
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 6920 26852 6972 26858
rect 6920 26794 6972 26800
rect 6932 22778 6960 26794
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 7484 18154 7512 26930
rect 9692 26858 9720 27270
rect 10428 27130 10456 29294
rect 10966 29200 11022 30000
rect 11610 29200 11666 30000
rect 12254 29322 12310 30000
rect 12898 29322 12954 30000
rect 12254 29294 12388 29322
rect 12254 29200 12310 29294
rect 10508 27464 10560 27470
rect 10508 27406 10560 27412
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10520 27062 10548 27406
rect 10980 27402 11008 29200
rect 11624 27538 11652 29200
rect 11924 27772 12232 27781
rect 11924 27770 11930 27772
rect 11986 27770 12010 27772
rect 12066 27770 12090 27772
rect 12146 27770 12170 27772
rect 12226 27770 12232 27772
rect 11986 27718 11988 27770
rect 12168 27718 12170 27770
rect 11924 27716 11930 27718
rect 11986 27716 12010 27718
rect 12066 27716 12090 27718
rect 12146 27716 12170 27718
rect 12226 27716 12232 27718
rect 11924 27707 12232 27716
rect 12164 27600 12216 27606
rect 12164 27542 12216 27548
rect 11612 27532 11664 27538
rect 11612 27474 11664 27480
rect 12176 27402 12204 27542
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 10968 27396 11020 27402
rect 10968 27338 11020 27344
rect 12164 27396 12216 27402
rect 12164 27338 12216 27344
rect 10508 27056 10560 27062
rect 10508 26998 10560 27004
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 9680 26852 9732 26858
rect 9680 26794 9732 26800
rect 10612 24138 10640 26930
rect 11924 26684 12232 26693
rect 11924 26682 11930 26684
rect 11986 26682 12010 26684
rect 12066 26682 12090 26684
rect 12146 26682 12170 26684
rect 12226 26682 12232 26684
rect 11986 26630 11988 26682
rect 12168 26630 12170 26682
rect 11924 26628 11930 26630
rect 11986 26628 12010 26630
rect 12066 26628 12090 26630
rect 12146 26628 12170 26630
rect 12226 26628 12232 26630
rect 11924 26619 12232 26628
rect 11924 25596 12232 25605
rect 11924 25594 11930 25596
rect 11986 25594 12010 25596
rect 12066 25594 12090 25596
rect 12146 25594 12170 25596
rect 12226 25594 12232 25596
rect 11986 25542 11988 25594
rect 12168 25542 12170 25594
rect 11924 25540 11930 25542
rect 11986 25540 12010 25542
rect 12066 25540 12090 25542
rect 12146 25540 12170 25542
rect 12226 25540 12232 25542
rect 11924 25531 12232 25540
rect 11924 24508 12232 24517
rect 11924 24506 11930 24508
rect 11986 24506 12010 24508
rect 12066 24506 12090 24508
rect 12146 24506 12170 24508
rect 12226 24506 12232 24508
rect 11986 24454 11988 24506
rect 12168 24454 12170 24506
rect 11924 24452 11930 24454
rect 11986 24452 12010 24454
rect 12066 24452 12090 24454
rect 12146 24452 12170 24454
rect 12226 24452 12232 24454
rect 11924 24443 12232 24452
rect 10600 24132 10652 24138
rect 10600 24074 10652 24080
rect 11924 23420 12232 23429
rect 11924 23418 11930 23420
rect 11986 23418 12010 23420
rect 12066 23418 12090 23420
rect 12146 23418 12170 23420
rect 12226 23418 12232 23420
rect 11986 23366 11988 23418
rect 12168 23366 12170 23418
rect 11924 23364 11930 23366
rect 11986 23364 12010 23366
rect 12066 23364 12090 23366
rect 12146 23364 12170 23366
rect 12226 23364 12232 23366
rect 11924 23355 12232 23364
rect 11924 22332 12232 22341
rect 11924 22330 11930 22332
rect 11986 22330 12010 22332
rect 12066 22330 12090 22332
rect 12146 22330 12170 22332
rect 12226 22330 12232 22332
rect 11986 22278 11988 22330
rect 12168 22278 12170 22330
rect 11924 22276 11930 22278
rect 11986 22276 12010 22278
rect 12066 22276 12090 22278
rect 12146 22276 12170 22278
rect 12226 22276 12232 22278
rect 11924 22267 12232 22276
rect 11924 21244 12232 21253
rect 11924 21242 11930 21244
rect 11986 21242 12010 21244
rect 12066 21242 12090 21244
rect 12146 21242 12170 21244
rect 12226 21242 12232 21244
rect 11986 21190 11988 21242
rect 12168 21190 12170 21242
rect 11924 21188 11930 21190
rect 11986 21188 12010 21190
rect 12066 21188 12090 21190
rect 12146 21188 12170 21190
rect 12226 21188 12232 21190
rect 11924 21179 12232 21188
rect 11924 20156 12232 20165
rect 11924 20154 11930 20156
rect 11986 20154 12010 20156
rect 12066 20154 12090 20156
rect 12146 20154 12170 20156
rect 12226 20154 12232 20156
rect 11986 20102 11988 20154
rect 12168 20102 12170 20154
rect 11924 20100 11930 20102
rect 11986 20100 12010 20102
rect 12066 20100 12090 20102
rect 12146 20100 12170 20102
rect 12226 20100 12232 20102
rect 11924 20091 12232 20100
rect 11924 19068 12232 19077
rect 11924 19066 11930 19068
rect 11986 19066 12010 19068
rect 12066 19066 12090 19068
rect 12146 19066 12170 19068
rect 12226 19066 12232 19068
rect 11986 19014 11988 19066
rect 12168 19014 12170 19066
rect 11924 19012 11930 19014
rect 11986 19012 12010 19014
rect 12066 19012 12090 19014
rect 12146 19012 12170 19014
rect 12226 19012 12232 19014
rect 11924 19003 12232 19012
rect 12268 18329 12296 27406
rect 12360 26994 12388 29294
rect 12820 29294 12954 29322
rect 12820 27470 12848 29294
rect 12898 29200 12954 29294
rect 13542 29322 13598 30000
rect 14186 29322 14242 30000
rect 14830 29322 14886 30000
rect 15474 29322 15530 30000
rect 16118 29322 16174 30000
rect 16762 29322 16818 30000
rect 13542 29294 13676 29322
rect 13542 29200 13598 29294
rect 12808 27464 12860 27470
rect 12808 27406 12860 27412
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12544 26586 12572 26726
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 13096 25770 13124 27406
rect 13648 27130 13676 29294
rect 14186 29294 14320 29322
rect 14186 29200 14242 29294
rect 14292 27606 14320 29294
rect 14830 29294 14964 29322
rect 14830 29200 14886 29294
rect 14936 27606 14964 29294
rect 15474 29294 15608 29322
rect 15474 29200 15530 29294
rect 15580 27606 15608 29294
rect 16118 29294 16528 29322
rect 16118 29200 16174 29294
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 14924 27600 14976 27606
rect 14924 27542 14976 27548
rect 15568 27600 15620 27606
rect 15568 27542 15620 27548
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 15108 27464 15160 27470
rect 15108 27406 15160 27412
rect 15752 27464 15804 27470
rect 16500 27452 16528 29294
rect 16762 29294 17080 29322
rect 16762 29200 16818 29294
rect 16580 27464 16632 27470
rect 16500 27424 16580 27452
rect 15752 27406 15804 27412
rect 16580 27406 16632 27412
rect 13636 27124 13688 27130
rect 13636 27066 13688 27072
rect 13544 27056 13596 27062
rect 13544 26998 13596 27004
rect 13556 26314 13584 26998
rect 14476 26518 14504 27406
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14464 26512 14516 26518
rect 14464 26454 14516 26460
rect 13544 26308 13596 26314
rect 13544 26250 13596 26256
rect 13084 25764 13136 25770
rect 13084 25706 13136 25712
rect 12254 18320 12310 18329
rect 12254 18255 12310 18264
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 7472 18148 7524 18154
rect 7472 18090 7524 18096
rect 11924 17980 12232 17989
rect 11924 17978 11930 17980
rect 11986 17978 12010 17980
rect 12066 17978 12090 17980
rect 12146 17978 12170 17980
rect 12226 17978 12232 17980
rect 11986 17926 11988 17978
rect 12168 17926 12170 17978
rect 11924 17924 11930 17926
rect 11986 17924 12010 17926
rect 12066 17924 12090 17926
rect 12146 17924 12170 17926
rect 12226 17924 12232 17926
rect 11924 17915 12232 17924
rect 11924 16892 12232 16901
rect 11924 16890 11930 16892
rect 11986 16890 12010 16892
rect 12066 16890 12090 16892
rect 12146 16890 12170 16892
rect 12226 16890 12232 16892
rect 11986 16838 11988 16890
rect 12168 16838 12170 16890
rect 11924 16836 11930 16838
rect 11986 16836 12010 16838
rect 12066 16836 12090 16838
rect 12146 16836 12170 16838
rect 12226 16836 12232 16838
rect 11924 16827 12232 16836
rect 11924 15804 12232 15813
rect 11924 15802 11930 15804
rect 11986 15802 12010 15804
rect 12066 15802 12090 15804
rect 12146 15802 12170 15804
rect 12226 15802 12232 15804
rect 11986 15750 11988 15802
rect 12168 15750 12170 15802
rect 11924 15748 11930 15750
rect 11986 15748 12010 15750
rect 12066 15748 12090 15750
rect 12146 15748 12170 15750
rect 12226 15748 12232 15750
rect 11924 15739 12232 15748
rect 12360 15366 12388 18226
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12544 17762 12572 17818
rect 12440 17740 12492 17746
rect 12544 17734 12664 17762
rect 12440 17682 12492 17688
rect 12452 17338 12480 17682
rect 12636 17678 12664 17734
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12544 17490 12572 17614
rect 12716 17536 12768 17542
rect 12544 17484 12716 17490
rect 12544 17478 12768 17484
rect 12544 17462 12756 17478
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3528 3194 3556 3470
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3712 3058 3740 5646
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 4540 2922 4568 3062
rect 4816 3058 4844 11290
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 5000 3058 5028 3402
rect 7116 3058 7144 3946
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9324 3126 9352 3470
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9968 3058 9996 3606
rect 11716 3602 11744 15098
rect 12728 15094 12756 16050
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 11924 14716 12232 14725
rect 11924 14714 11930 14716
rect 11986 14714 12010 14716
rect 12066 14714 12090 14716
rect 12146 14714 12170 14716
rect 12226 14714 12232 14716
rect 11986 14662 11988 14714
rect 12168 14662 12170 14714
rect 11924 14660 11930 14662
rect 11986 14660 12010 14662
rect 12066 14660 12090 14662
rect 12146 14660 12170 14662
rect 12226 14660 12232 14662
rect 11924 14651 12232 14660
rect 11924 13628 12232 13637
rect 11924 13626 11930 13628
rect 11986 13626 12010 13628
rect 12066 13626 12090 13628
rect 12146 13626 12170 13628
rect 12226 13626 12232 13628
rect 11986 13574 11988 13626
rect 12168 13574 12170 13626
rect 11924 13572 11930 13574
rect 11986 13572 12010 13574
rect 12066 13572 12090 13574
rect 12146 13572 12170 13574
rect 12226 13572 12232 13574
rect 11924 13563 12232 13572
rect 11924 12540 12232 12549
rect 11924 12538 11930 12540
rect 11986 12538 12010 12540
rect 12066 12538 12090 12540
rect 12146 12538 12170 12540
rect 12226 12538 12232 12540
rect 11986 12486 11988 12538
rect 12168 12486 12170 12538
rect 11924 12484 11930 12486
rect 11986 12484 12010 12486
rect 12066 12484 12090 12486
rect 12146 12484 12170 12486
rect 12226 12484 12232 12486
rect 11924 12475 12232 12484
rect 11924 11452 12232 11461
rect 11924 11450 11930 11452
rect 11986 11450 12010 11452
rect 12066 11450 12090 11452
rect 12146 11450 12170 11452
rect 12226 11450 12232 11452
rect 11986 11398 11988 11450
rect 12168 11398 12170 11450
rect 11924 11396 11930 11398
rect 11986 11396 12010 11398
rect 12066 11396 12090 11398
rect 12146 11396 12170 11398
rect 12226 11396 12232 11398
rect 11924 11387 12232 11396
rect 14462 11384 14518 11393
rect 14752 11354 14780 26930
rect 15120 15473 15148 27406
rect 15764 27062 15792 27406
rect 15660 27056 15712 27062
rect 15660 26998 15712 27004
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15672 26858 15700 26998
rect 17052 26994 17080 29294
rect 18050 29200 18106 30000
rect 18694 29322 18750 30000
rect 18616 29294 18750 29322
rect 18064 27606 18092 29200
rect 18616 27606 18644 29294
rect 18694 29200 18750 29294
rect 19338 29322 19394 30000
rect 19338 29294 19656 29322
rect 19338 29200 19394 29294
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 18604 27600 18656 27606
rect 18604 27542 18656 27548
rect 19628 27470 19656 29294
rect 19982 29200 20038 30000
rect 20626 29200 20682 30000
rect 21270 29322 21326 30000
rect 21914 29322 21970 30000
rect 22558 29322 22614 30000
rect 23202 29322 23258 30000
rect 21270 29294 21404 29322
rect 21270 29200 21326 29294
rect 19996 27606 20024 29200
rect 20640 27606 20668 29200
rect 19984 27600 20036 27606
rect 19984 27542 20036 27548
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 21376 27470 21404 29294
rect 21914 29294 22048 29322
rect 21914 29200 21970 29294
rect 22020 27606 22048 29294
rect 22558 29294 22876 29322
rect 22558 29200 22614 29294
rect 22008 27600 22060 27606
rect 22008 27542 22060 27548
rect 22560 27600 22612 27606
rect 22560 27542 22612 27548
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20352 27464 20404 27470
rect 20352 27406 20404 27412
rect 21364 27464 21416 27470
rect 21364 27406 21416 27412
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 17132 27396 17184 27402
rect 17132 27338 17184 27344
rect 17040 26988 17092 26994
rect 17040 26930 17092 26936
rect 15660 26852 15712 26858
rect 15660 26794 15712 26800
rect 17144 26790 17172 27338
rect 18064 26994 18092 27406
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 16856 26784 16908 26790
rect 16856 26726 16908 26732
rect 17132 26784 17184 26790
rect 17132 26726 17184 26732
rect 16868 26382 16896 26726
rect 18248 26450 18276 27406
rect 18800 27130 18828 27406
rect 19800 27328 19852 27334
rect 19800 27270 19852 27276
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 16856 26376 16908 26382
rect 16856 26318 16908 26324
rect 19444 26246 19472 26930
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 17960 25220 18012 25226
rect 17960 25162 18012 25168
rect 17972 23730 18000 25162
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 15106 15464 15162 15473
rect 15106 15399 15162 15408
rect 16500 15162 16528 21966
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18248 13938 18276 14214
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18248 13734 18276 13874
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 14462 11319 14464 11328
rect 14516 11319 14518 11328
rect 14740 11348 14792 11354
rect 14464 11290 14516 11296
rect 14740 11290 14792 11296
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 11924 10364 12232 10373
rect 11924 10362 11930 10364
rect 11986 10362 12010 10364
rect 12066 10362 12090 10364
rect 12146 10362 12170 10364
rect 12226 10362 12232 10364
rect 11986 10310 11988 10362
rect 12168 10310 12170 10362
rect 11924 10308 11930 10310
rect 11986 10308 12010 10310
rect 12066 10308 12090 10310
rect 12146 10308 12170 10310
rect 12226 10308 12232 10310
rect 11924 10299 12232 10308
rect 15396 9586 15424 11086
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 11924 9276 12232 9285
rect 11924 9274 11930 9276
rect 11986 9274 12010 9276
rect 12066 9274 12090 9276
rect 12146 9274 12170 9276
rect 12226 9274 12232 9276
rect 11986 9222 11988 9274
rect 12168 9222 12170 9274
rect 11924 9220 11930 9222
rect 11986 9220 12010 9222
rect 12066 9220 12090 9222
rect 12146 9220 12170 9222
rect 12226 9220 12232 9222
rect 11924 9211 12232 9220
rect 11924 8188 12232 8197
rect 11924 8186 11930 8188
rect 11986 8186 12010 8188
rect 12066 8186 12090 8188
rect 12146 8186 12170 8188
rect 12226 8186 12232 8188
rect 11986 8134 11988 8186
rect 12168 8134 12170 8186
rect 11924 8132 11930 8134
rect 11986 8132 12010 8134
rect 12066 8132 12090 8134
rect 12146 8132 12170 8134
rect 12226 8132 12232 8134
rect 11924 8123 12232 8132
rect 11924 7100 12232 7109
rect 11924 7098 11930 7100
rect 11986 7098 12010 7100
rect 12066 7098 12090 7100
rect 12146 7098 12170 7100
rect 12226 7098 12232 7100
rect 11986 7046 11988 7098
rect 12168 7046 12170 7098
rect 11924 7044 11930 7046
rect 11986 7044 12010 7046
rect 12066 7044 12090 7046
rect 12146 7044 12170 7046
rect 12226 7044 12232 7046
rect 11924 7035 12232 7044
rect 11924 6012 12232 6021
rect 11924 6010 11930 6012
rect 11986 6010 12010 6012
rect 12066 6010 12090 6012
rect 12146 6010 12170 6012
rect 12226 6010 12232 6012
rect 11986 5958 11988 6010
rect 12168 5958 12170 6010
rect 11924 5956 11930 5958
rect 11986 5956 12010 5958
rect 12066 5956 12090 5958
rect 12146 5956 12170 5958
rect 12226 5956 12232 5958
rect 11924 5947 12232 5956
rect 11924 4924 12232 4933
rect 11924 4922 11930 4924
rect 11986 4922 12010 4924
rect 12066 4922 12090 4924
rect 12146 4922 12170 4924
rect 12226 4922 12232 4924
rect 11986 4870 11988 4922
rect 12168 4870 12170 4922
rect 11924 4868 11930 4870
rect 11986 4868 12010 4870
rect 12066 4868 12090 4870
rect 12146 4868 12170 4870
rect 12226 4868 12232 4870
rect 11924 4859 12232 4868
rect 11924 3836 12232 3845
rect 11924 3834 11930 3836
rect 11986 3834 12010 3836
rect 12066 3834 12090 3836
rect 12146 3834 12170 3836
rect 12226 3834 12232 3836
rect 11986 3782 11988 3834
rect 12168 3782 12170 3834
rect 11924 3780 11930 3782
rect 11986 3780 12010 3782
rect 12066 3780 12090 3782
rect 12146 3780 12170 3782
rect 12226 3780 12232 3782
rect 11924 3771 12232 3780
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 13832 3058 13860 3402
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3884 2372 3936 2378
rect 3884 2314 3936 2320
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 2962 2136 3018 2145
rect 2962 2071 3018 2080
rect 2872 1828 2924 1834
rect 2872 1770 2924 1776
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3252 800 3280 2246
rect 3896 800 3924 2314
rect 4066 912 4122 921
rect 4172 898 4200 2518
rect 4908 2446 4936 2790
rect 5552 2446 5580 2790
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 4264 1562 4292 2246
rect 4252 1556 4304 1562
rect 4252 1498 4304 1504
rect 4122 870 4200 898
rect 4066 847 4122 856
rect 5184 800 5212 2246
rect 5828 800 5856 2382
rect 6472 800 6500 2790
rect 9784 2446 9812 2790
rect 9968 2446 9996 2858
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 10244 2514 10272 2790
rect 11924 2748 12232 2757
rect 11924 2746 11930 2748
rect 11986 2746 12010 2748
rect 12066 2746 12090 2748
rect 12146 2746 12170 2748
rect 12226 2746 12232 2748
rect 11986 2694 11988 2746
rect 12168 2694 12170 2746
rect 11924 2692 11930 2694
rect 11986 2692 12010 2694
rect 12066 2692 12090 2694
rect 12146 2692 12170 2694
rect 12226 2692 12232 2694
rect 11924 2683 12232 2692
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 7760 800 7788 2382
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 8220 1970 8248 2246
rect 8208 1964 8260 1970
rect 8208 1906 8260 1912
rect 8404 800 8432 2246
rect 9048 800 9076 2246
rect 9692 800 9720 2246
rect 10336 800 10364 2246
rect 10520 1766 10548 2382
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10508 1760 10560 1766
rect 10508 1702 10560 1708
rect 10980 800 11008 2246
rect 11624 800 11652 2314
rect 12268 800 12296 2382
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12360 1698 12388 2246
rect 12348 1692 12400 1698
rect 12348 1634 12400 1640
rect 12912 800 12940 2382
rect 13556 800 13584 2790
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14200 800 14228 2382
rect 14384 1426 14412 2382
rect 15396 2378 15424 9522
rect 15856 2514 15884 11086
rect 16592 3194 16620 11766
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17236 4554 17264 5102
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 14372 1420 14424 1426
rect 14372 1362 14424 1368
rect 15488 800 15516 2246
rect 15764 2038 15792 2382
rect 15752 2032 15804 2038
rect 15752 1974 15804 1980
rect 16132 800 16160 2382
rect 16776 800 16804 2994
rect 17236 2922 17264 3674
rect 17972 2922 18000 4422
rect 18248 3534 18276 13262
rect 18800 11762 18828 14962
rect 18984 12374 19012 14962
rect 19076 13530 19104 14962
rect 19812 13938 19840 27270
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19892 21412 19944 21418
rect 19892 21354 19944 21360
rect 19904 15162 19932 21354
rect 19996 15348 20024 26930
rect 20076 26512 20128 26518
rect 20076 26454 20128 26460
rect 20088 16794 20116 26454
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20272 16250 20300 27406
rect 20364 27130 20392 27406
rect 20444 27396 20496 27402
rect 20444 27338 20496 27344
rect 20456 27130 20484 27338
rect 21272 27328 21324 27334
rect 21272 27270 21324 27276
rect 20352 27124 20404 27130
rect 20352 27066 20404 27072
rect 20444 27124 20496 27130
rect 20444 27066 20496 27072
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20456 26518 20484 26930
rect 21284 26858 21312 27270
rect 22204 26994 22232 27406
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 21272 26852 21324 26858
rect 21272 26794 21324 26800
rect 20444 26512 20496 26518
rect 20444 26454 20496 26460
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 19996 15320 20116 15348
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19076 12782 19104 13262
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 18984 11762 19012 12310
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18616 7410 18644 11494
rect 18800 11218 18828 11698
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18892 11393 18920 11562
rect 18878 11384 18934 11393
rect 18878 11319 18934 11328
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 19168 4078 19196 13670
rect 19536 12850 19564 13670
rect 19628 13394 19656 13806
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19720 12782 19748 13262
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19812 12646 19840 13874
rect 19890 13696 19946 13705
rect 19890 13631 19946 13640
rect 19904 13462 19932 13631
rect 20088 13569 20116 15320
rect 20364 14414 20392 26250
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20074 13560 20130 13569
rect 19984 13524 20036 13530
rect 20074 13495 20130 13504
rect 19984 13466 20036 13472
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 19996 13326 20024 13466
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19708 11756 19760 11762
rect 19904 11744 19932 12786
rect 19996 12617 20024 13262
rect 19982 12608 20038 12617
rect 19982 12543 20038 12552
rect 20088 12442 20116 13262
rect 20180 12850 20208 13398
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 19760 11716 19932 11744
rect 19708 11698 19760 11704
rect 20088 11694 20116 12378
rect 20180 12102 20208 12378
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20180 11558 20208 11766
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16960 1630 16988 2382
rect 16948 1624 17000 1630
rect 16948 1566 17000 1572
rect 17420 800 17448 2790
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 18064 800 18092 2382
rect 18708 800 18736 2450
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19352 800 19380 2246
rect 19996 800 20024 2790
rect 20272 2774 20300 14214
rect 20364 12850 20392 14350
rect 20456 14006 20484 26454
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20456 12782 20484 13194
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20548 12102 20576 16526
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20732 15162 20760 15370
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14278 20668 14894
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20824 13920 20852 18226
rect 21100 16794 21128 25638
rect 22020 20602 22048 26386
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 21822 16960 21878 16969
rect 21822 16895 21878 16904
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 21652 16590 21680 16730
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21376 16182 21404 16526
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20916 15162 20944 15506
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20732 13892 20852 13920
rect 20732 13326 20760 13892
rect 20812 13796 20864 13802
rect 20812 13738 20864 13744
rect 20824 13530 20852 13738
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12850 20760 13126
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20916 12714 20944 14282
rect 21100 13716 21128 15438
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21192 14618 21220 14758
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21192 13870 21220 14010
rect 21376 14006 21404 14758
rect 21652 14618 21680 16526
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21560 14006 21588 14214
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21548 14000 21600 14006
rect 21548 13942 21600 13948
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21744 13734 21772 14418
rect 21272 13728 21324 13734
rect 21100 13688 21220 13716
rect 21088 13320 21140 13326
rect 21192 13297 21220 13688
rect 21272 13670 21324 13676
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21088 13262 21140 13268
rect 21178 13288 21234 13297
rect 21100 12866 21128 13262
rect 21178 13223 21234 13232
rect 21008 12838 21128 12866
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20824 12306 20852 12582
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20732 11558 20760 12174
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20916 10810 20944 12650
rect 21008 12434 21036 12838
rect 21008 12406 21128 12434
rect 21100 12374 21128 12406
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21008 11694 21036 12174
rect 20996 11688 21048 11694
rect 21100 11665 21128 12174
rect 20996 11630 21048 11636
rect 21086 11656 21142 11665
rect 21086 11591 21142 11600
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20732 3466 20760 6598
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 20180 2746 20300 2774
rect 20180 2514 20208 2746
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 20824 2446 20852 7754
rect 21008 5778 21036 11494
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21192 3398 21220 13223
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 21284 2774 21312 13670
rect 21836 13530 21864 16895
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21928 15570 21956 16050
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21928 14385 21956 15506
rect 22020 15026 22048 18702
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22204 15706 22232 16050
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22204 15434 22232 15642
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22020 14929 22048 14962
rect 22006 14920 22062 14929
rect 22006 14855 22062 14864
rect 22112 14822 22140 15098
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22100 14408 22152 14414
rect 21914 14376 21970 14385
rect 22100 14350 22152 14356
rect 21914 14311 21970 14320
rect 22112 13977 22140 14350
rect 22098 13968 22154 13977
rect 22098 13903 22154 13912
rect 22204 13870 22232 14486
rect 22296 14414 22324 23462
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 22480 19378 22508 20470
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22374 17640 22430 17649
rect 22374 17575 22430 17584
rect 22388 17270 22416 17575
rect 22376 17264 22428 17270
rect 22376 17206 22428 17212
rect 22480 15162 22508 19314
rect 22572 16250 22600 27542
rect 22848 27470 22876 29294
rect 23124 29294 23258 29322
rect 23124 27538 23152 29294
rect 23202 29200 23258 29294
rect 23846 29322 23902 30000
rect 24490 29322 24546 30000
rect 25778 29322 25834 30000
rect 23846 29294 24164 29322
rect 23846 29200 23902 29294
rect 23112 27532 23164 27538
rect 23112 27474 23164 27480
rect 22836 27464 22888 27470
rect 22836 27406 22888 27412
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 22898 27228 23206 27237
rect 22898 27226 22904 27228
rect 22960 27226 22984 27228
rect 23040 27226 23064 27228
rect 23120 27226 23144 27228
rect 23200 27226 23206 27228
rect 22960 27174 22962 27226
rect 23142 27174 23144 27226
rect 22898 27172 22904 27174
rect 22960 27172 22984 27174
rect 23040 27172 23064 27174
rect 23120 27172 23144 27174
rect 23200 27172 23206 27174
rect 22898 27163 23206 27172
rect 23400 26761 23428 27406
rect 24136 26994 24164 29294
rect 24490 29294 24624 29322
rect 24490 29200 24546 29294
rect 24596 27606 24624 29294
rect 25778 29294 26004 29322
rect 25778 29200 25834 29294
rect 25872 27668 25924 27674
rect 25872 27610 25924 27616
rect 24584 27600 24636 27606
rect 24584 27542 24636 27548
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 25410 27432 25466 27441
rect 23940 26988 23992 26994
rect 24124 26988 24176 26994
rect 23992 26948 24072 26976
rect 23940 26930 23992 26936
rect 24044 26790 24072 26948
rect 24124 26930 24176 26936
rect 23940 26784 23992 26790
rect 23386 26752 23442 26761
rect 23940 26726 23992 26732
rect 24032 26784 24084 26790
rect 24032 26726 24084 26732
rect 23386 26687 23442 26696
rect 23952 26314 23980 26726
rect 23388 26308 23440 26314
rect 23388 26250 23440 26256
rect 23940 26308 23992 26314
rect 23940 26250 23992 26256
rect 22898 26140 23206 26149
rect 22898 26138 22904 26140
rect 22960 26138 22984 26140
rect 23040 26138 23064 26140
rect 23120 26138 23144 26140
rect 23200 26138 23206 26140
rect 22960 26086 22962 26138
rect 23142 26086 23144 26138
rect 22898 26084 22904 26086
rect 22960 26084 22984 26086
rect 23040 26084 23064 26086
rect 23120 26084 23144 26086
rect 23200 26084 23206 26086
rect 22898 26075 23206 26084
rect 22898 25052 23206 25061
rect 22898 25050 22904 25052
rect 22960 25050 22984 25052
rect 23040 25050 23064 25052
rect 23120 25050 23144 25052
rect 23200 25050 23206 25052
rect 22960 24998 22962 25050
rect 23142 24998 23144 25050
rect 22898 24996 22904 24998
rect 22960 24996 22984 24998
rect 23040 24996 23064 24998
rect 23120 24996 23144 24998
rect 23200 24996 23206 24998
rect 22898 24987 23206 24996
rect 22744 24676 22796 24682
rect 22744 24618 22796 24624
rect 22756 17338 22784 24618
rect 22898 23964 23206 23973
rect 22898 23962 22904 23964
rect 22960 23962 22984 23964
rect 23040 23962 23064 23964
rect 23120 23962 23144 23964
rect 23200 23962 23206 23964
rect 22960 23910 22962 23962
rect 23142 23910 23144 23962
rect 22898 23908 22904 23910
rect 22960 23908 22984 23910
rect 23040 23908 23064 23910
rect 23120 23908 23144 23910
rect 23200 23908 23206 23910
rect 22898 23899 23206 23908
rect 22898 22876 23206 22885
rect 22898 22874 22904 22876
rect 22960 22874 22984 22876
rect 23040 22874 23064 22876
rect 23120 22874 23144 22876
rect 23200 22874 23206 22876
rect 22960 22822 22962 22874
rect 23142 22822 23144 22874
rect 22898 22820 22904 22822
rect 22960 22820 22984 22822
rect 23040 22820 23064 22822
rect 23120 22820 23144 22822
rect 23200 22820 23206 22822
rect 22898 22811 23206 22820
rect 22898 21788 23206 21797
rect 22898 21786 22904 21788
rect 22960 21786 22984 21788
rect 23040 21786 23064 21788
rect 23120 21786 23144 21788
rect 23200 21786 23206 21788
rect 22960 21734 22962 21786
rect 23142 21734 23144 21786
rect 22898 21732 22904 21734
rect 22960 21732 22984 21734
rect 23040 21732 23064 21734
rect 23120 21732 23144 21734
rect 23200 21732 23206 21734
rect 22898 21723 23206 21732
rect 22898 20700 23206 20709
rect 22898 20698 22904 20700
rect 22960 20698 22984 20700
rect 23040 20698 23064 20700
rect 23120 20698 23144 20700
rect 23200 20698 23206 20700
rect 22960 20646 22962 20698
rect 23142 20646 23144 20698
rect 22898 20644 22904 20646
rect 22960 20644 22984 20646
rect 23040 20644 23064 20646
rect 23120 20644 23144 20646
rect 23200 20644 23206 20646
rect 22898 20635 23206 20644
rect 22898 19612 23206 19621
rect 22898 19610 22904 19612
rect 22960 19610 22984 19612
rect 23040 19610 23064 19612
rect 23120 19610 23144 19612
rect 23200 19610 23206 19612
rect 22960 19558 22962 19610
rect 23142 19558 23144 19610
rect 22898 19556 22904 19558
rect 22960 19556 22984 19558
rect 23040 19556 23064 19558
rect 23120 19556 23144 19558
rect 23200 19556 23206 19558
rect 22898 19547 23206 19556
rect 22898 18524 23206 18533
rect 22898 18522 22904 18524
rect 22960 18522 22984 18524
rect 23040 18522 23064 18524
rect 23120 18522 23144 18524
rect 23200 18522 23206 18524
rect 22960 18470 22962 18522
rect 23142 18470 23144 18522
rect 22898 18468 22904 18470
rect 22960 18468 22984 18470
rect 23040 18468 23064 18470
rect 23120 18468 23144 18470
rect 23200 18468 23206 18470
rect 22898 18459 23206 18468
rect 22898 17436 23206 17445
rect 22898 17434 22904 17436
rect 22960 17434 22984 17436
rect 23040 17434 23064 17436
rect 23120 17434 23144 17436
rect 23200 17434 23206 17436
rect 22960 17382 22962 17434
rect 23142 17382 23144 17434
rect 22898 17380 22904 17382
rect 22960 17380 22984 17382
rect 23040 17380 23064 17382
rect 23120 17380 23144 17382
rect 23200 17380 23206 17382
rect 22898 17371 23206 17380
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22898 16348 23206 16357
rect 22898 16346 22904 16348
rect 22960 16346 22984 16348
rect 23040 16346 23064 16348
rect 23120 16346 23144 16348
rect 23200 16346 23206 16348
rect 22960 16294 22962 16346
rect 23142 16294 23144 16346
rect 22898 16292 22904 16294
rect 22960 16292 22984 16294
rect 23040 16292 23064 16294
rect 23120 16292 23144 16294
rect 23200 16292 23206 16294
rect 22898 16283 23206 16292
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22296 13870 22324 14350
rect 22192 13864 22244 13870
rect 22098 13832 22154 13841
rect 22192 13806 22244 13812
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22098 13767 22100 13776
rect 22152 13767 22154 13776
rect 22100 13738 22152 13744
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 22388 13326 22416 14962
rect 22572 14550 22600 15302
rect 22560 14544 22612 14550
rect 22560 14486 22612 14492
rect 22572 14346 22600 14486
rect 22560 14340 22612 14346
rect 22560 14282 22612 14288
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22480 13818 22508 14214
rect 22480 13802 22600 13818
rect 22480 13796 22612 13802
rect 22480 13790 22560 13796
rect 22560 13738 22612 13744
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 22020 12918 22048 13262
rect 22480 13190 22508 13670
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22572 13326 22600 13466
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21376 11830 21404 12378
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21560 12102 21588 12174
rect 21548 12096 21600 12102
rect 21548 12038 21600 12044
rect 21364 11824 21416 11830
rect 21364 11766 21416 11772
rect 21560 11393 21588 12038
rect 21546 11384 21602 11393
rect 21546 11319 21602 11328
rect 21560 10062 21588 11319
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 21192 2746 21312 2774
rect 21192 2582 21220 2746
rect 21180 2576 21232 2582
rect 21180 2518 21232 2524
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 20640 800 20668 2246
rect 21284 800 21312 2246
rect 21928 800 21956 2382
rect 22020 1494 22048 12854
rect 22664 4486 22692 15438
rect 22756 15144 22784 16050
rect 23296 16040 23348 16046
rect 23296 15982 23348 15988
rect 22898 15260 23206 15269
rect 22898 15258 22904 15260
rect 22960 15258 22984 15260
rect 23040 15258 23064 15260
rect 23120 15258 23144 15260
rect 23200 15258 23206 15260
rect 22960 15206 22962 15258
rect 23142 15206 23144 15258
rect 22898 15204 22904 15206
rect 22960 15204 22984 15206
rect 23040 15204 23064 15206
rect 23120 15204 23144 15206
rect 23200 15204 23206 15206
rect 22898 15195 23206 15204
rect 22756 15116 22876 15144
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 22756 14618 22784 14962
rect 22744 14612 22796 14618
rect 22744 14554 22796 14560
rect 22848 14521 22876 15116
rect 23308 15026 23336 15982
rect 23400 15337 23428 26250
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23768 18290 23796 20402
rect 24596 18970 24624 27406
rect 25410 27367 25412 27376
rect 25464 27367 25466 27376
rect 25412 27338 25464 27344
rect 25884 27334 25912 27610
rect 25976 27470 26004 29294
rect 26422 29200 26478 30000
rect 27066 29322 27122 30000
rect 27710 29322 27766 30000
rect 27066 29294 27200 29322
rect 27066 29200 27122 29294
rect 26436 27606 26464 29200
rect 27172 27606 27200 29294
rect 27710 29294 27844 29322
rect 27710 29200 27766 29294
rect 27816 27606 27844 29294
rect 28354 29200 28410 30000
rect 28998 29322 29054 30000
rect 29642 29322 29698 30000
rect 28998 29294 29132 29322
rect 28998 29200 29054 29294
rect 26424 27600 26476 27606
rect 26424 27542 26476 27548
rect 27160 27600 27212 27606
rect 27160 27542 27212 27548
rect 27804 27600 27856 27606
rect 27804 27542 27856 27548
rect 28368 27470 28396 29200
rect 29104 27470 29132 29294
rect 29642 29294 29776 29322
rect 29642 29200 29698 29294
rect 29748 27606 29776 29294
rect 30286 29200 30342 30000
rect 30930 29322 30986 30000
rect 30852 29294 30986 29322
rect 29736 27600 29788 27606
rect 29736 27542 29788 27548
rect 29368 27532 29420 27538
rect 29368 27474 29420 27480
rect 25964 27464 26016 27470
rect 25964 27406 26016 27412
rect 26700 27464 26752 27470
rect 26700 27406 26752 27412
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 28356 27464 28408 27470
rect 28356 27406 28408 27412
rect 29092 27464 29144 27470
rect 29092 27406 29144 27412
rect 25872 27328 25924 27334
rect 25872 27270 25924 27276
rect 26056 27328 26108 27334
rect 26056 27270 26108 27276
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 25964 26376 26016 26382
rect 25964 26318 26016 26324
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 24768 20392 24820 20398
rect 24768 20334 24820 20340
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 24492 18828 24544 18834
rect 24492 18770 24544 18776
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23952 15434 23980 17138
rect 24216 17128 24268 17134
rect 24044 17088 24216 17116
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 23386 15328 23442 15337
rect 23386 15263 23442 15272
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23112 14816 23164 14822
rect 23110 14784 23112 14793
rect 23164 14784 23166 14793
rect 23110 14719 23166 14728
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 22834 14512 22890 14521
rect 22834 14447 22890 14456
rect 23308 14385 23336 14554
rect 23294 14376 23350 14385
rect 23294 14311 23350 14320
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22756 13938 22784 14214
rect 22898 14172 23206 14181
rect 22898 14170 22904 14172
rect 22960 14170 22984 14172
rect 23040 14170 23064 14172
rect 23120 14170 23144 14172
rect 23200 14170 23206 14172
rect 22960 14118 22962 14170
rect 23142 14118 23144 14170
rect 22898 14116 22904 14118
rect 22960 14116 22984 14118
rect 23040 14116 23064 14118
rect 23120 14116 23144 14118
rect 23200 14116 23206 14118
rect 22898 14107 23206 14116
rect 22834 13968 22890 13977
rect 22744 13932 22796 13938
rect 22834 13903 22836 13912
rect 22744 13874 22796 13880
rect 22888 13903 22890 13912
rect 22836 13874 22888 13880
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22756 12986 22784 13670
rect 23308 13530 23336 13806
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 22898 13084 23206 13093
rect 22898 13082 22904 13084
rect 22960 13082 22984 13084
rect 23040 13082 23064 13084
rect 23120 13082 23144 13084
rect 23200 13082 23206 13084
rect 22960 13030 22962 13082
rect 23142 13030 23144 13082
rect 22898 13028 22904 13030
rect 22960 13028 22984 13030
rect 23040 13028 23064 13030
rect 23120 13028 23144 13030
rect 23200 13028 23206 13030
rect 22898 13019 23206 13028
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 23400 12646 23428 15030
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23492 12782 23520 14010
rect 23572 13796 23624 13802
rect 23572 13738 23624 13744
rect 23584 13258 23612 13738
rect 23676 13734 23704 14010
rect 23860 13938 23888 14758
rect 23940 14340 23992 14346
rect 23940 14282 23992 14288
rect 23952 14249 23980 14282
rect 23938 14240 23994 14249
rect 23938 14175 23994 14184
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 24044 13818 24072 17088
rect 24216 17070 24268 17076
rect 24214 15736 24270 15745
rect 24214 15671 24270 15680
rect 24228 15026 24256 15671
rect 24308 15156 24360 15162
rect 24308 15098 24360 15104
rect 24320 15026 24348 15098
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24136 14657 24164 14894
rect 24122 14648 24178 14657
rect 24122 14583 24178 14592
rect 23952 13790 24072 13818
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23756 13728 23808 13734
rect 23756 13670 23808 13676
rect 23664 13388 23716 13394
rect 23768 13376 23796 13670
rect 23716 13348 23796 13376
rect 23664 13330 23716 13336
rect 23952 13258 23980 13790
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 23572 13252 23624 13258
rect 23572 13194 23624 13200
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 22898 11996 23206 12005
rect 22898 11994 22904 11996
rect 22960 11994 22984 11996
rect 23040 11994 23064 11996
rect 23120 11994 23144 11996
rect 23200 11994 23206 11996
rect 22960 11942 22962 11994
rect 23142 11942 23144 11994
rect 22898 11940 22904 11942
rect 22960 11940 22984 11942
rect 23040 11940 23064 11942
rect 23120 11940 23144 11942
rect 23200 11940 23206 11942
rect 22898 11931 23206 11940
rect 23492 11218 23520 12174
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23584 11218 23612 11834
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 22898 10908 23206 10917
rect 22898 10906 22904 10908
rect 22960 10906 22984 10908
rect 23040 10906 23064 10908
rect 23120 10906 23144 10908
rect 23200 10906 23206 10908
rect 22960 10854 22962 10906
rect 23142 10854 23144 10906
rect 22898 10852 22904 10854
rect 22960 10852 22984 10854
rect 23040 10852 23064 10854
rect 23120 10852 23144 10854
rect 23200 10852 23206 10854
rect 22898 10843 23206 10852
rect 23388 10600 23440 10606
rect 23388 10542 23440 10548
rect 22898 9820 23206 9829
rect 22898 9818 22904 9820
rect 22960 9818 22984 9820
rect 23040 9818 23064 9820
rect 23120 9818 23144 9820
rect 23200 9818 23206 9820
rect 22960 9766 22962 9818
rect 23142 9766 23144 9818
rect 22898 9764 22904 9766
rect 22960 9764 22984 9766
rect 23040 9764 23064 9766
rect 23120 9764 23144 9766
rect 23200 9764 23206 9766
rect 22898 9755 23206 9764
rect 23400 8838 23428 10542
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 22898 8732 23206 8741
rect 22898 8730 22904 8732
rect 22960 8730 22984 8732
rect 23040 8730 23064 8732
rect 23120 8730 23144 8732
rect 23200 8730 23206 8732
rect 22960 8678 22962 8730
rect 23142 8678 23144 8730
rect 22898 8676 22904 8678
rect 22960 8676 22984 8678
rect 23040 8676 23064 8678
rect 23120 8676 23144 8678
rect 23200 8676 23206 8678
rect 22898 8667 23206 8676
rect 22898 7644 23206 7653
rect 22898 7642 22904 7644
rect 22960 7642 22984 7644
rect 23040 7642 23064 7644
rect 23120 7642 23144 7644
rect 23200 7642 23206 7644
rect 22960 7590 22962 7642
rect 23142 7590 23144 7642
rect 22898 7588 22904 7590
rect 22960 7588 22984 7590
rect 23040 7588 23064 7590
rect 23120 7588 23144 7590
rect 23200 7588 23206 7590
rect 22898 7579 23206 7588
rect 22898 6556 23206 6565
rect 22898 6554 22904 6556
rect 22960 6554 22984 6556
rect 23040 6554 23064 6556
rect 23120 6554 23144 6556
rect 23200 6554 23206 6556
rect 22960 6502 22962 6554
rect 23142 6502 23144 6554
rect 22898 6500 22904 6502
rect 22960 6500 22984 6502
rect 23040 6500 23064 6502
rect 23120 6500 23144 6502
rect 23200 6500 23206 6502
rect 22898 6491 23206 6500
rect 22898 5468 23206 5477
rect 22898 5466 22904 5468
rect 22960 5466 22984 5468
rect 23040 5466 23064 5468
rect 23120 5466 23144 5468
rect 23200 5466 23206 5468
rect 22960 5414 22962 5466
rect 23142 5414 23144 5466
rect 22898 5412 22904 5414
rect 22960 5412 22984 5414
rect 23040 5412 23064 5414
rect 23120 5412 23144 5414
rect 23200 5412 23206 5414
rect 22898 5403 23206 5412
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22898 4380 23206 4389
rect 22898 4378 22904 4380
rect 22960 4378 22984 4380
rect 23040 4378 23064 4380
rect 23120 4378 23144 4380
rect 23200 4378 23206 4380
rect 22960 4326 22962 4378
rect 23142 4326 23144 4378
rect 22898 4324 22904 4326
rect 22960 4324 22984 4326
rect 23040 4324 23064 4326
rect 23120 4324 23144 4326
rect 23200 4324 23206 4326
rect 22898 4315 23206 4324
rect 22744 3664 22796 3670
rect 22744 3606 22796 3612
rect 22756 3058 22784 3606
rect 22898 3292 23206 3301
rect 22898 3290 22904 3292
rect 22960 3290 22984 3292
rect 23040 3290 23064 3292
rect 23120 3290 23144 3292
rect 23200 3290 23206 3292
rect 22960 3238 22962 3290
rect 23142 3238 23144 3290
rect 22898 3236 22904 3238
rect 22960 3236 22984 3238
rect 23040 3236 23064 3238
rect 23120 3236 23144 3238
rect 23200 3236 23206 3238
rect 22898 3227 23206 3236
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 22848 2514 22876 2790
rect 23296 2576 23348 2582
rect 23296 2518 23348 2524
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22204 1970 22232 2246
rect 22898 2204 23206 2213
rect 22898 2202 22904 2204
rect 22960 2202 22984 2204
rect 23040 2202 23064 2204
rect 23120 2202 23144 2204
rect 23200 2202 23206 2204
rect 22960 2150 22962 2202
rect 23142 2150 23144 2202
rect 22898 2148 22904 2150
rect 22960 2148 22984 2150
rect 23040 2148 23064 2150
rect 23120 2148 23144 2150
rect 23200 2148 23206 2150
rect 22898 2139 23206 2148
rect 22192 1964 22244 1970
rect 22192 1906 22244 1912
rect 22008 1488 22060 1494
rect 22008 1430 22060 1436
rect 23308 1170 23336 2518
rect 23584 1426 23612 9386
rect 23676 5234 23704 13194
rect 23938 13152 23994 13161
rect 23938 13087 23994 13096
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23768 11898 23796 12718
rect 23952 12714 23980 13087
rect 24044 12889 24072 13670
rect 24228 13326 24256 14962
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24320 14074 24348 14758
rect 24412 14414 24440 14894
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24412 14074 24440 14350
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 24504 13954 24532 18770
rect 24780 18766 24808 20334
rect 24952 19372 25004 19378
rect 24952 19314 25004 19320
rect 24964 18766 24992 19314
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24964 17678 24992 18022
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24676 17604 24728 17610
rect 24676 17546 24728 17552
rect 24584 17536 24636 17542
rect 24582 17504 24584 17513
rect 24636 17504 24638 17513
rect 24582 17439 24638 17448
rect 24688 17270 24716 17546
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24676 17128 24728 17134
rect 24674 17096 24676 17105
rect 24728 17096 24730 17105
rect 24964 17066 24992 17138
rect 24674 17031 24730 17040
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 25320 16448 25372 16454
rect 25320 16390 25372 16396
rect 25042 16280 25098 16289
rect 24584 16244 24636 16250
rect 25042 16215 25098 16224
rect 24584 16186 24636 16192
rect 24596 16046 24624 16186
rect 25056 16114 25084 16215
rect 25332 16182 25360 16390
rect 25320 16176 25372 16182
rect 25320 16118 25372 16124
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 24688 14346 24716 15030
rect 24780 14550 24808 16050
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24768 14544 24820 14550
rect 24768 14486 24820 14492
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24676 14340 24728 14346
rect 24676 14282 24728 14288
rect 24320 13926 24532 13954
rect 24676 13932 24728 13938
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24030 12880 24086 12889
rect 24030 12815 24086 12824
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 24136 2774 24164 13262
rect 24214 13016 24270 13025
rect 24214 12951 24270 12960
rect 24228 12714 24256 12951
rect 24216 12708 24268 12714
rect 24216 12650 24268 12656
rect 24320 11762 24348 13926
rect 24676 13874 24728 13880
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24492 13796 24544 13802
rect 24492 13738 24544 13744
rect 24504 12986 24532 13738
rect 24596 13394 24624 13806
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24412 12170 24440 12786
rect 24688 12481 24716 13874
rect 24780 13530 24808 14350
rect 24872 14278 24900 15098
rect 25056 15026 25084 16050
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25410 15872 25466 15881
rect 25240 15502 25268 15846
rect 25410 15807 25466 15816
rect 25424 15570 25452 15807
rect 25412 15564 25464 15570
rect 25412 15506 25464 15512
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25136 15360 25188 15366
rect 25136 15302 25188 15308
rect 25148 15026 25176 15302
rect 25516 15162 25544 26182
rect 25872 20528 25924 20534
rect 25872 20470 25924 20476
rect 25884 19446 25912 20470
rect 25872 19440 25924 19446
rect 25872 19382 25924 19388
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25596 16448 25648 16454
rect 25596 16390 25648 16396
rect 25608 16250 25636 16390
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25608 15162 25636 15642
rect 25700 15434 25728 16934
rect 25792 16658 25820 17682
rect 25884 16833 25912 19382
rect 25976 18426 26004 26318
rect 25964 18420 26016 18426
rect 25964 18362 26016 18368
rect 25870 16824 25926 16833
rect 25870 16759 25926 16768
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25792 16289 25820 16594
rect 25964 16584 26016 16590
rect 25964 16526 26016 16532
rect 25778 16280 25834 16289
rect 25778 16215 25834 16224
rect 25976 15706 26004 16526
rect 26068 16153 26096 27270
rect 26252 26994 26280 27270
rect 26240 26988 26292 26994
rect 26240 26930 26292 26936
rect 26516 26988 26568 26994
rect 26516 26930 26568 26936
rect 26424 26784 26476 26790
rect 26424 26726 26476 26732
rect 26436 26625 26464 26726
rect 26422 26616 26478 26625
rect 26422 26551 26478 26560
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26252 18222 26280 18906
rect 26240 18216 26292 18222
rect 26240 18158 26292 18164
rect 26240 18080 26292 18086
rect 26240 18022 26292 18028
rect 26252 17202 26280 18022
rect 26332 17536 26384 17542
rect 26330 17504 26332 17513
rect 26384 17504 26386 17513
rect 26330 17439 26386 17448
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 26252 16572 26280 16934
rect 26332 16584 26384 16590
rect 26252 16544 26332 16572
rect 26332 16526 26384 16532
rect 26148 16516 26200 16522
rect 26148 16458 26200 16464
rect 26160 16402 26188 16458
rect 26160 16374 26280 16402
rect 26146 16280 26202 16289
rect 26252 16250 26280 16374
rect 26146 16215 26202 16224
rect 26240 16244 26292 16250
rect 26054 16144 26110 16153
rect 26054 16079 26110 16088
rect 25964 15700 26016 15706
rect 25964 15642 26016 15648
rect 26160 15502 26188 16215
rect 26240 16186 26292 16192
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 25688 15428 25740 15434
rect 25688 15370 25740 15376
rect 26056 15360 26108 15366
rect 25976 15308 26056 15314
rect 25976 15302 26108 15308
rect 25976 15286 26096 15302
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25596 15156 25648 15162
rect 25596 15098 25648 15104
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 25594 14512 25650 14521
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24964 14074 24992 14486
rect 25594 14447 25650 14456
rect 25608 14414 25636 14447
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25870 14376 25926 14385
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25240 13938 25268 14214
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25792 13870 25820 14350
rect 25870 14311 25926 14320
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 24768 13524 24820 13530
rect 24768 13466 24820 13472
rect 25042 13424 25098 13433
rect 25700 13394 25728 13670
rect 25884 13462 25912 14311
rect 25872 13456 25924 13462
rect 25872 13398 25924 13404
rect 25042 13359 25098 13368
rect 25504 13388 25556 13394
rect 25056 13326 25084 13359
rect 25504 13330 25556 13336
rect 25688 13388 25740 13394
rect 25688 13330 25740 13336
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 25424 12986 25452 13262
rect 25516 12986 25544 13330
rect 25976 13308 26004 15286
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 26068 14278 26096 14554
rect 26160 14385 26188 15438
rect 26528 15026 26556 26930
rect 26712 26518 26740 27406
rect 27252 27396 27304 27402
rect 27252 27338 27304 27344
rect 27264 26518 27292 27338
rect 28080 27328 28132 27334
rect 28080 27270 28132 27276
rect 27528 26988 27580 26994
rect 27528 26930 27580 26936
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27436 26784 27488 26790
rect 27436 26726 27488 26732
rect 27342 26616 27398 26625
rect 27342 26551 27398 26560
rect 26700 26512 26752 26518
rect 26700 26454 26752 26460
rect 27252 26512 27304 26518
rect 27252 26454 27304 26460
rect 26700 26308 26752 26314
rect 26700 26250 26752 26256
rect 26712 26042 26740 26250
rect 26700 26036 26752 26042
rect 26700 25978 26752 25984
rect 26792 25832 26844 25838
rect 26792 25774 26844 25780
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26620 19334 26648 25638
rect 26620 19306 26740 19334
rect 26516 15020 26568 15026
rect 26516 14962 26568 14968
rect 26240 14952 26292 14958
rect 26240 14894 26292 14900
rect 26146 14376 26202 14385
rect 26146 14311 26202 14320
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 26252 13938 26280 14894
rect 26424 14816 26476 14822
rect 26424 14758 26476 14764
rect 26516 14816 26568 14822
rect 26516 14758 26568 14764
rect 26436 14074 26464 14758
rect 26528 14414 26556 14758
rect 26608 14544 26660 14550
rect 26608 14486 26660 14492
rect 26712 14498 26740 19306
rect 26804 14958 26832 25774
rect 27356 22094 27384 26551
rect 27448 26382 27476 26726
rect 27540 26489 27568 26930
rect 27526 26480 27582 26489
rect 27724 26450 27752 26930
rect 27802 26752 27858 26761
rect 27802 26687 27858 26696
rect 27526 26415 27582 26424
rect 27712 26444 27764 26450
rect 27712 26386 27764 26392
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 27724 22094 27752 26386
rect 27816 26382 27844 26687
rect 27804 26376 27856 26382
rect 27804 26318 27856 26324
rect 27356 22066 27568 22094
rect 27724 22066 27936 22094
rect 27068 18964 27120 18970
rect 27068 18906 27120 18912
rect 26976 18352 27028 18358
rect 26976 18294 27028 18300
rect 26988 17610 27016 18294
rect 26976 17604 27028 17610
rect 26976 17546 27028 17552
rect 26976 17128 27028 17134
rect 26976 17070 27028 17076
rect 26988 16289 27016 17070
rect 26974 16280 27030 16289
rect 26974 16215 27030 16224
rect 26884 16108 26936 16114
rect 26884 16050 26936 16056
rect 26792 14952 26844 14958
rect 26792 14894 26844 14900
rect 26896 14618 26924 16050
rect 26988 16046 27016 16215
rect 26976 16040 27028 16046
rect 26976 15982 27028 15988
rect 26976 15904 27028 15910
rect 26976 15846 27028 15852
rect 26988 15502 27016 15846
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 26516 14408 26568 14414
rect 26516 14350 26568 14356
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26516 14068 26568 14074
rect 26516 14010 26568 14016
rect 26240 13932 26292 13938
rect 26160 13892 26240 13920
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 25884 13280 26004 13308
rect 26068 13297 26096 13466
rect 26054 13288 26110 13297
rect 25228 12980 25280 12986
rect 25412 12980 25464 12986
rect 25280 12940 25360 12968
rect 25228 12922 25280 12928
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24674 12472 24730 12481
rect 24674 12407 24730 12416
rect 24400 12164 24452 12170
rect 24400 12106 24452 12112
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24228 11150 24256 11630
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24320 11257 24348 11494
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24306 11248 24362 11257
rect 24306 11183 24362 11192
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24306 11112 24362 11121
rect 24306 11047 24308 11056
rect 24360 11047 24362 11056
rect 24308 11018 24360 11024
rect 24504 10538 24532 11290
rect 24596 11150 24624 11698
rect 24872 11354 24900 12786
rect 25228 12640 25280 12646
rect 25228 12582 25280 12588
rect 25240 12442 25268 12582
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 25148 12345 25176 12378
rect 25134 12336 25190 12345
rect 24952 12300 25004 12306
rect 25134 12271 25190 12280
rect 24952 12242 25004 12248
rect 24964 12186 24992 12242
rect 25228 12232 25280 12238
rect 25226 12200 25228 12209
rect 25280 12200 25282 12209
rect 24964 12158 25084 12186
rect 25056 12102 25084 12158
rect 25226 12135 25282 12144
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 25044 12096 25096 12102
rect 25332 12073 25360 12940
rect 25412 12922 25464 12928
rect 25504 12980 25556 12986
rect 25504 12922 25556 12928
rect 25044 12038 25096 12044
rect 25318 12064 25374 12073
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24492 10532 24544 10538
rect 24492 10474 24544 10480
rect 24596 3534 24624 11086
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24780 4690 24808 5102
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 24964 3534 24992 12038
rect 25056 11937 25084 12038
rect 25318 11999 25374 12008
rect 25042 11928 25098 11937
rect 25042 11863 25098 11872
rect 25320 11824 25372 11830
rect 25320 11766 25372 11772
rect 25686 11792 25742 11801
rect 25332 11286 25360 11766
rect 25884 11762 25912 13280
rect 26054 13223 26110 13232
rect 26056 13184 26108 13190
rect 26056 13126 26108 13132
rect 26068 12753 26096 13126
rect 26160 13025 26188 13892
rect 26240 13874 26292 13880
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26240 13184 26292 13190
rect 26344 13161 26372 13874
rect 26436 13734 26464 14010
rect 26424 13728 26476 13734
rect 26424 13670 26476 13676
rect 26424 13388 26476 13394
rect 26424 13330 26476 13336
rect 26240 13126 26292 13132
rect 26330 13152 26386 13161
rect 26146 13016 26202 13025
rect 26146 12951 26202 12960
rect 26148 12912 26200 12918
rect 26252 12900 26280 13126
rect 26330 13087 26386 13096
rect 26436 12968 26464 13330
rect 26528 13326 26556 14010
rect 26620 14006 26648 14486
rect 26712 14470 26832 14498
rect 26700 14408 26752 14414
rect 26698 14376 26700 14385
rect 26752 14376 26754 14385
rect 26698 14311 26754 14320
rect 26608 14000 26660 14006
rect 26608 13942 26660 13948
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 26608 13796 26660 13802
rect 26608 13738 26660 13744
rect 26620 13326 26648 13738
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26516 12980 26568 12986
rect 26436 12940 26516 12968
rect 26516 12922 26568 12928
rect 26200 12872 26280 12900
rect 26514 12880 26570 12889
rect 26148 12854 26200 12860
rect 26514 12815 26516 12824
rect 26568 12815 26570 12824
rect 26516 12786 26568 12792
rect 26712 12782 26740 13874
rect 26804 13705 26832 14470
rect 26884 13932 26936 13938
rect 26884 13874 26936 13880
rect 26896 13802 26924 13874
rect 26884 13796 26936 13802
rect 26884 13738 26936 13744
rect 26790 13696 26846 13705
rect 26790 13631 26846 13640
rect 26700 12776 26752 12782
rect 26054 12744 26110 12753
rect 26700 12718 26752 12724
rect 26054 12679 26110 12688
rect 26330 12608 26386 12617
rect 26330 12543 26386 12552
rect 26056 12300 26108 12306
rect 26056 12242 26108 12248
rect 26068 11898 26096 12242
rect 26344 12238 26372 12543
rect 26804 12238 26832 13631
rect 26882 13560 26938 13569
rect 26882 13495 26938 13504
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 25686 11727 25742 11736
rect 25780 11756 25832 11762
rect 25700 11694 25728 11727
rect 25780 11698 25832 11704
rect 25872 11756 25924 11762
rect 25872 11698 25924 11704
rect 26056 11756 26108 11762
rect 26056 11698 26108 11704
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 25792 11558 25820 11698
rect 25596 11552 25648 11558
rect 25594 11520 25596 11529
rect 25780 11552 25832 11558
rect 25648 11520 25650 11529
rect 25780 11494 25832 11500
rect 25594 11455 25650 11464
rect 25884 11393 25912 11698
rect 25964 11688 26016 11694
rect 26068 11665 26096 11698
rect 25964 11630 26016 11636
rect 26054 11656 26110 11665
rect 25870 11384 25926 11393
rect 25870 11319 25926 11328
rect 25320 11280 25372 11286
rect 25320 11222 25372 11228
rect 25780 11144 25832 11150
rect 25976 11132 26004 11630
rect 26054 11591 26110 11600
rect 25832 11104 26004 11132
rect 25780 11086 25832 11092
rect 25044 11076 25096 11082
rect 25044 11018 25096 11024
rect 25056 10266 25084 11018
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 25240 10062 25268 10406
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25792 5710 25820 11086
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 25884 10606 25912 10950
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 25148 5370 25176 5646
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24228 2990 24256 3130
rect 24216 2984 24268 2990
rect 24216 2926 24268 2932
rect 24044 2746 24164 2774
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 23572 1420 23624 1426
rect 23572 1362 23624 1368
rect 23216 1142 23336 1170
rect 23216 800 23244 1142
rect 23860 800 23888 2246
rect 23952 1426 23980 2382
rect 24044 2310 24072 2746
rect 24228 2446 24256 2926
rect 24412 2922 24440 3470
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24780 3058 24808 3334
rect 25424 3058 25452 4082
rect 25780 3392 25832 3398
rect 25780 3334 25832 3340
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 24400 2916 24452 2922
rect 24400 2858 24452 2864
rect 25136 2848 25188 2854
rect 25136 2790 25188 2796
rect 25412 2848 25464 2854
rect 25412 2790 25464 2796
rect 24216 2440 24268 2446
rect 24216 2382 24268 2388
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 24032 2304 24084 2310
rect 24400 2304 24452 2310
rect 24032 2246 24084 2252
rect 24214 2272 24270 2281
rect 24400 2246 24452 2252
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24214 2207 24270 2216
rect 24228 1766 24256 2207
rect 24412 1834 24440 2246
rect 24400 1828 24452 1834
rect 24400 1770 24452 1776
rect 24216 1760 24268 1766
rect 24216 1702 24268 1708
rect 23940 1420 23992 1426
rect 23940 1362 23992 1368
rect 24504 800 24532 2246
rect 24780 2106 24808 2382
rect 24768 2100 24820 2106
rect 24768 2042 24820 2048
rect 25148 800 25176 2790
rect 25424 2446 25452 2790
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 25792 800 25820 3334
rect 25884 1290 25912 10542
rect 26068 9674 26096 11591
rect 26160 10810 26188 12174
rect 26422 12064 26478 12073
rect 26422 11999 26478 12008
rect 26436 11898 26464 11999
rect 26514 11928 26570 11937
rect 26424 11892 26476 11898
rect 26514 11863 26570 11872
rect 26792 11892 26844 11898
rect 26424 11834 26476 11840
rect 26528 11762 26556 11863
rect 26792 11834 26844 11840
rect 26332 11756 26384 11762
rect 26332 11698 26384 11704
rect 26516 11756 26568 11762
rect 26516 11698 26568 11704
rect 26344 11529 26372 11698
rect 26804 11626 26832 11834
rect 26792 11620 26844 11626
rect 26792 11562 26844 11568
rect 26330 11520 26386 11529
rect 26330 11455 26386 11464
rect 26238 11248 26294 11257
rect 26238 11183 26294 11192
rect 26252 11082 26280 11183
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26148 10804 26200 10810
rect 26148 10746 26200 10752
rect 26068 9646 26280 9674
rect 26148 5636 26200 5642
rect 26148 5578 26200 5584
rect 26160 4622 26188 5578
rect 26148 4616 26200 4622
rect 26148 4558 26200 4564
rect 26160 3126 26188 4558
rect 26148 3120 26200 3126
rect 25962 3088 26018 3097
rect 26148 3062 26200 3068
rect 25962 3023 25964 3032
rect 26016 3023 26018 3032
rect 25964 2994 26016 3000
rect 26252 2990 26280 9646
rect 26344 5114 26372 11455
rect 26896 11286 26924 13495
rect 26988 12617 27016 15438
rect 27080 14822 27108 18906
rect 27436 18284 27488 18290
rect 27436 18226 27488 18232
rect 27158 17776 27214 17785
rect 27344 17740 27396 17746
rect 27158 17711 27214 17720
rect 27172 17678 27200 17711
rect 27264 17700 27344 17728
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 27264 17134 27292 17700
rect 27344 17682 27396 17688
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27448 16454 27476 18226
rect 27436 16448 27488 16454
rect 27436 16390 27488 16396
rect 27342 16008 27398 16017
rect 27342 15943 27398 15952
rect 27356 15366 27384 15943
rect 27448 15745 27476 16390
rect 27434 15736 27490 15745
rect 27434 15671 27490 15680
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27342 15192 27398 15201
rect 27540 15162 27568 22066
rect 27804 19236 27856 19242
rect 27804 19178 27856 19184
rect 27816 18834 27844 19178
rect 27908 19174 27936 22066
rect 27988 19440 28040 19446
rect 27988 19382 28040 19388
rect 27896 19168 27948 19174
rect 27896 19110 27948 19116
rect 27804 18828 27856 18834
rect 27804 18770 27856 18776
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27724 18222 27752 18702
rect 27896 18624 27948 18630
rect 27896 18566 27948 18572
rect 27908 18222 27936 18566
rect 28000 18306 28028 19382
rect 28092 19242 28120 27270
rect 28184 26858 28212 27406
rect 28540 27328 28592 27334
rect 28540 27270 28592 27276
rect 28264 26920 28316 26926
rect 28264 26862 28316 26868
rect 28172 26852 28224 26858
rect 28172 26794 28224 26800
rect 28276 22094 28304 26862
rect 28184 22066 28304 22094
rect 28080 19236 28132 19242
rect 28080 19178 28132 19184
rect 28000 18290 28120 18306
rect 28000 18284 28132 18290
rect 28000 18278 28080 18284
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27896 18216 27948 18222
rect 27896 18158 27948 18164
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27632 17746 27660 18022
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27724 17626 27752 18158
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 27632 17598 27752 17626
rect 27632 15638 27660 17598
rect 27816 17270 27844 18022
rect 27804 17264 27856 17270
rect 27804 17206 27856 17212
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27724 16017 27752 16050
rect 27710 16008 27766 16017
rect 27710 15943 27766 15952
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27802 15872 27858 15881
rect 27620 15632 27672 15638
rect 27620 15574 27672 15580
rect 27342 15127 27344 15136
rect 27396 15127 27398 15136
rect 27528 15156 27580 15162
rect 27344 15098 27396 15104
rect 27528 15098 27580 15104
rect 27540 15042 27568 15098
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27356 15014 27568 15042
rect 27068 14816 27120 14822
rect 27068 14758 27120 14764
rect 27068 14612 27120 14618
rect 27068 14554 27120 14560
rect 27080 14521 27108 14554
rect 27066 14512 27122 14521
rect 27066 14447 27122 14456
rect 27264 14414 27292 14962
rect 27252 14408 27304 14414
rect 27252 14350 27304 14356
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 26974 12608 27030 12617
rect 26974 12543 27030 12552
rect 26884 11280 26936 11286
rect 26884 11222 26936 11228
rect 27080 10674 27108 14282
rect 27264 13938 27292 14350
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 27264 12102 27292 12582
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27252 12096 27304 12102
rect 27252 12038 27304 12044
rect 27172 11150 27200 12038
rect 27160 11144 27212 11150
rect 27160 11086 27212 11092
rect 27356 11014 27384 15014
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27448 14226 27476 14894
rect 27540 14822 27568 14894
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27540 14346 27568 14758
rect 27528 14340 27580 14346
rect 27528 14282 27580 14288
rect 27448 14198 27568 14226
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27160 11008 27212 11014
rect 27160 10950 27212 10956
rect 27344 11008 27396 11014
rect 27344 10950 27396 10956
rect 27172 10742 27200 10950
rect 27160 10736 27212 10742
rect 27160 10678 27212 10684
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 26424 10532 26476 10538
rect 26424 10474 26476 10480
rect 26436 6798 26464 10474
rect 27448 8498 27476 13806
rect 27540 13530 27568 14198
rect 27632 13802 27660 15574
rect 27724 15026 27752 15846
rect 27802 15807 27858 15816
rect 27816 15706 27844 15807
rect 27804 15700 27856 15706
rect 27804 15642 27856 15648
rect 27894 15600 27950 15609
rect 27894 15535 27896 15544
rect 27948 15535 27950 15544
rect 27896 15506 27948 15512
rect 28000 15178 28028 18278
rect 28080 18226 28132 18232
rect 28080 17536 28132 17542
rect 28080 17478 28132 17484
rect 28092 17202 28120 17478
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 28078 16824 28134 16833
rect 28078 16759 28134 16768
rect 28092 15366 28120 16759
rect 28184 16658 28212 22066
rect 28264 19168 28316 19174
rect 28264 19110 28316 19116
rect 28276 18630 28304 19110
rect 28264 18624 28316 18630
rect 28264 18566 28316 18572
rect 28276 16969 28304 18566
rect 28552 18426 28580 27270
rect 28724 26988 28776 26994
rect 28724 26930 28776 26936
rect 28540 18420 28592 18426
rect 28540 18362 28592 18368
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28368 17898 28396 18226
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 28368 17870 28580 17898
rect 28448 17808 28500 17814
rect 28448 17750 28500 17756
rect 28460 17649 28488 17750
rect 28552 17746 28580 17870
rect 28540 17740 28592 17746
rect 28540 17682 28592 17688
rect 28446 17640 28502 17649
rect 28356 17604 28408 17610
rect 28446 17575 28502 17584
rect 28356 17546 28408 17552
rect 28368 17338 28396 17546
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28356 17128 28408 17134
rect 28354 17096 28356 17105
rect 28408 17096 28410 17105
rect 28354 17031 28410 17040
rect 28540 16992 28592 16998
rect 28262 16960 28318 16969
rect 28262 16895 28318 16904
rect 28538 16960 28540 16969
rect 28592 16960 28594 16969
rect 28538 16895 28594 16904
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 28080 15360 28132 15366
rect 28080 15302 28132 15308
rect 27816 15150 28028 15178
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 27712 14340 27764 14346
rect 27712 14282 27764 14288
rect 27620 13796 27672 13802
rect 27620 13738 27672 13744
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27540 13326 27568 13466
rect 27528 13320 27580 13326
rect 27528 13262 27580 13268
rect 27620 12708 27672 12714
rect 27620 12650 27672 12656
rect 27632 12170 27660 12650
rect 27620 12164 27672 12170
rect 27620 12106 27672 12112
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27632 11354 27660 11630
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27724 9674 27752 14282
rect 27816 13977 27844 15150
rect 27988 14816 28040 14822
rect 27988 14758 28040 14764
rect 27896 14476 27948 14482
rect 27896 14418 27948 14424
rect 27908 14278 27936 14418
rect 27896 14272 27948 14278
rect 27896 14214 27948 14220
rect 27802 13968 27858 13977
rect 27802 13903 27858 13912
rect 27896 13456 27948 13462
rect 27894 13424 27896 13433
rect 27948 13424 27950 13433
rect 27894 13359 27950 13368
rect 27804 13184 27856 13190
rect 27804 13126 27856 13132
rect 27816 12442 27844 13126
rect 27804 12436 27856 12442
rect 28000 12434 28028 14758
rect 28184 14657 28212 16594
rect 28448 16584 28500 16590
rect 28448 16526 28500 16532
rect 28262 16280 28318 16289
rect 28262 16215 28318 16224
rect 28276 15502 28304 16215
rect 28264 15496 28316 15502
rect 28264 15438 28316 15444
rect 28170 14648 28226 14657
rect 28170 14583 28226 14592
rect 28184 14362 28212 14583
rect 28184 14334 28304 14362
rect 28080 14000 28132 14006
rect 28078 13968 28080 13977
rect 28132 13968 28134 13977
rect 28078 13903 28134 13912
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 27804 12378 27856 12384
rect 27908 12406 28028 12434
rect 27632 9646 27752 9674
rect 27436 8492 27488 8498
rect 27436 8434 27488 8440
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 26436 5574 26464 6734
rect 26424 5568 26476 5574
rect 26424 5510 26476 5516
rect 26436 5302 26464 5510
rect 26424 5296 26476 5302
rect 26424 5238 26476 5244
rect 26344 5086 26464 5114
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 26344 2553 26372 2994
rect 26436 2666 26464 5086
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 26712 3534 26740 4966
rect 27528 4480 27580 4486
rect 27528 4422 27580 4428
rect 27540 4282 27568 4422
rect 27528 4276 27580 4282
rect 27528 4218 27580 4224
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 26608 3392 26660 3398
rect 26608 3334 26660 3340
rect 26436 2638 26556 2666
rect 26528 2582 26556 2638
rect 26424 2576 26476 2582
rect 26330 2544 26386 2553
rect 26424 2518 26476 2524
rect 26516 2576 26568 2582
rect 26516 2518 26568 2524
rect 26330 2479 26386 2488
rect 26148 2372 26200 2378
rect 26148 2314 26200 2320
rect 26160 1562 26188 2314
rect 26330 1864 26386 1873
rect 26330 1799 26332 1808
rect 26384 1799 26386 1808
rect 26332 1770 26384 1776
rect 26056 1556 26108 1562
rect 26056 1498 26108 1504
rect 26148 1556 26200 1562
rect 26148 1498 26200 1504
rect 26068 1358 26096 1498
rect 26056 1352 26108 1358
rect 26056 1294 26108 1300
rect 25872 1284 25924 1290
rect 25872 1226 25924 1232
rect 26436 800 26464 2518
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 26528 1834 26556 2382
rect 26516 1828 26568 1834
rect 26516 1770 26568 1776
rect 26620 1766 26648 3334
rect 27252 2576 27304 2582
rect 27252 2518 27304 2524
rect 27528 2576 27580 2582
rect 27528 2518 27580 2524
rect 26976 2372 27028 2378
rect 26976 2314 27028 2320
rect 26988 1834 27016 2314
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 26976 1828 27028 1834
rect 26976 1770 27028 1776
rect 26608 1760 26660 1766
rect 26608 1702 26660 1708
rect 27080 800 27108 2246
rect 27264 1601 27292 2518
rect 27540 2394 27568 2518
rect 27632 2514 27660 9646
rect 27712 4480 27764 4486
rect 27712 4422 27764 4428
rect 27724 3398 27752 4422
rect 27908 3738 27936 12406
rect 27986 12336 28042 12345
rect 27986 12271 28042 12280
rect 28000 11830 28028 12271
rect 28092 12170 28120 13806
rect 28276 13530 28304 14334
rect 28264 13524 28316 13530
rect 28264 13466 28316 13472
rect 28460 13462 28488 16526
rect 28644 16522 28672 18158
rect 28736 16726 28764 26930
rect 28816 26920 28868 26926
rect 29380 26897 29408 27474
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 28816 26862 28868 26868
rect 29366 26888 29422 26897
rect 28724 16720 28776 16726
rect 28724 16662 28776 16668
rect 28632 16516 28684 16522
rect 28632 16458 28684 16464
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28552 14929 28580 14962
rect 28538 14920 28594 14929
rect 28538 14855 28594 14864
rect 28540 14816 28592 14822
rect 28538 14784 28540 14793
rect 28592 14784 28594 14793
rect 28538 14719 28594 14728
rect 28644 13734 28672 16458
rect 28828 14618 28856 26862
rect 29932 26858 29960 27406
rect 30300 26976 30328 29200
rect 30852 27538 30880 29294
rect 30930 29200 30986 29294
rect 31574 29322 31630 30000
rect 32862 29322 32918 30000
rect 31574 29294 31708 29322
rect 31574 29200 31630 29294
rect 31300 27668 31352 27674
rect 31300 27610 31352 27616
rect 30840 27532 30892 27538
rect 30840 27474 30892 27480
rect 31116 27464 31168 27470
rect 31116 27406 31168 27412
rect 31206 27432 31262 27441
rect 30380 26988 30432 26994
rect 30300 26948 30380 26976
rect 30380 26930 30432 26936
rect 30392 26858 30788 26874
rect 29366 26823 29422 26832
rect 29920 26852 29972 26858
rect 29920 26794 29972 26800
rect 30012 26852 30064 26858
rect 30012 26794 30064 26800
rect 30392 26852 30800 26858
rect 30392 26846 30748 26852
rect 29642 26616 29698 26625
rect 29642 26551 29698 26560
rect 29656 26382 29684 26551
rect 29184 26376 29236 26382
rect 29184 26318 29236 26324
rect 29460 26376 29512 26382
rect 29460 26318 29512 26324
rect 29644 26376 29696 26382
rect 29644 26318 29696 26324
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 29012 17785 29040 17818
rect 28998 17776 29054 17785
rect 28998 17711 29054 17720
rect 29196 16454 29224 26318
rect 29184 16448 29236 16454
rect 29184 16390 29236 16396
rect 29184 16040 29236 16046
rect 29182 16008 29184 16017
rect 29236 16008 29238 16017
rect 29092 15972 29144 15978
rect 29182 15943 29238 15952
rect 29092 15914 29144 15920
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 28906 15328 28962 15337
rect 28906 15263 28962 15272
rect 28920 15094 28948 15263
rect 28908 15088 28960 15094
rect 28908 15030 28960 15036
rect 29012 15026 29040 15506
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 28908 14952 28960 14958
rect 28908 14894 28960 14900
rect 28816 14612 28868 14618
rect 28816 14554 28868 14560
rect 28920 14414 28948 14894
rect 28908 14408 28960 14414
rect 28908 14350 28960 14356
rect 28816 14340 28868 14346
rect 28816 14282 28868 14288
rect 28828 14249 28856 14282
rect 28814 14240 28870 14249
rect 28814 14175 28870 14184
rect 29104 14074 29132 15914
rect 29184 15428 29236 15434
rect 29184 15370 29236 15376
rect 29196 15026 29224 15370
rect 29184 15020 29236 15026
rect 29184 14962 29236 14968
rect 29276 14408 29328 14414
rect 29276 14350 29328 14356
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29184 14000 29236 14006
rect 29184 13942 29236 13948
rect 28724 13796 28776 13802
rect 28724 13738 28776 13744
rect 28632 13728 28684 13734
rect 28632 13670 28684 13676
rect 28448 13456 28500 13462
rect 28448 13398 28500 13404
rect 28460 12782 28488 13398
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 28448 12776 28500 12782
rect 28448 12718 28500 12724
rect 28172 12708 28224 12714
rect 28172 12650 28224 12656
rect 28080 12164 28132 12170
rect 28080 12106 28132 12112
rect 27988 11824 28040 11830
rect 27988 11766 28040 11772
rect 28184 11694 28212 12650
rect 28354 12472 28410 12481
rect 28354 12407 28410 12416
rect 28264 12368 28316 12374
rect 28262 12336 28264 12345
rect 28316 12336 28318 12345
rect 28262 12271 28318 12280
rect 28368 12073 28396 12407
rect 28354 12064 28410 12073
rect 28354 11999 28410 12008
rect 28460 11898 28488 12718
rect 28552 12442 28580 12922
rect 28540 12436 28592 12442
rect 28540 12378 28592 12384
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28172 11688 28224 11694
rect 28172 11630 28224 11636
rect 28080 10464 28132 10470
rect 28080 10406 28132 10412
rect 28092 9994 28120 10406
rect 28080 9988 28132 9994
rect 28080 9930 28132 9936
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 2774 27752 2994
rect 27724 2746 27844 2774
rect 27816 2650 27844 2746
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 27620 2508 27672 2514
rect 27620 2450 27672 2456
rect 27908 2446 27936 3334
rect 28552 3097 28580 3470
rect 28538 3088 28594 3097
rect 28538 3023 28594 3032
rect 27896 2440 27948 2446
rect 27540 2366 27660 2394
rect 27896 2382 27948 2388
rect 27250 1592 27306 1601
rect 27250 1527 27306 1536
rect 27632 1222 27660 2366
rect 27804 2372 27856 2378
rect 27804 2314 27856 2320
rect 27816 1902 27844 2314
rect 28264 2304 28316 2310
rect 28262 2272 28264 2281
rect 28316 2272 28318 2281
rect 28262 2207 28318 2216
rect 27804 1896 27856 1902
rect 27804 1838 27856 1844
rect 27712 1828 27764 1834
rect 27712 1770 27764 1776
rect 27620 1216 27672 1222
rect 27620 1158 27672 1164
rect 27724 800 27752 1770
rect 28644 1766 28672 12174
rect 28736 3398 28764 13738
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 28908 12708 28960 12714
rect 28908 12650 28960 12656
rect 28816 12436 28868 12442
rect 28816 12378 28868 12384
rect 28828 12345 28856 12378
rect 28814 12336 28870 12345
rect 28814 12271 28870 12280
rect 28920 12186 28948 12650
rect 28828 12158 28948 12186
rect 28828 11801 28856 12158
rect 28908 12096 28960 12102
rect 28906 12064 28908 12073
rect 28960 12064 28962 12073
rect 28906 11999 28962 12008
rect 28814 11792 28870 11801
rect 29012 11762 29040 13466
rect 29196 13394 29224 13942
rect 29184 13388 29236 13394
rect 29184 13330 29236 13336
rect 29184 13252 29236 13258
rect 29184 13194 29236 13200
rect 29196 12986 29224 13194
rect 29184 12980 29236 12986
rect 29184 12922 29236 12928
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 29104 12238 29132 12582
rect 29092 12232 29144 12238
rect 29092 12174 29144 12180
rect 28814 11727 28870 11736
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29184 11552 29236 11558
rect 29184 11494 29236 11500
rect 29196 11150 29224 11494
rect 29184 11144 29236 11150
rect 28906 11112 28962 11121
rect 29184 11086 29236 11092
rect 28906 11047 28962 11056
rect 28920 4486 28948 11047
rect 29288 10996 29316 14350
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29196 10968 29316 10996
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 29012 9926 29040 10610
rect 29092 10056 29144 10062
rect 29092 9998 29144 10004
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 28908 4480 28960 4486
rect 28908 4422 28960 4428
rect 29012 4010 29040 9862
rect 29104 9722 29132 9998
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 29196 7562 29224 10968
rect 29276 10668 29328 10674
rect 29276 10610 29328 10616
rect 29288 10266 29316 10610
rect 29276 10260 29328 10266
rect 29276 10202 29328 10208
rect 29104 7534 29224 7562
rect 29000 4004 29052 4010
rect 29000 3946 29052 3952
rect 28724 3392 28776 3398
rect 28724 3334 28776 3340
rect 28736 2774 28764 3334
rect 28736 2746 28856 2774
rect 28828 2106 28856 2746
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 28816 2100 28868 2106
rect 28816 2042 28868 2048
rect 28908 2100 28960 2106
rect 28908 2042 28960 2048
rect 28920 1970 28948 2042
rect 28908 1964 28960 1970
rect 28908 1906 28960 1912
rect 28632 1760 28684 1766
rect 28632 1702 28684 1708
rect 28356 1216 28408 1222
rect 28356 1158 28408 1164
rect 28368 800 28396 1158
rect 29012 800 29040 2314
rect 29104 1358 29132 7534
rect 29380 5370 29408 14010
rect 29472 11218 29500 26318
rect 30024 26246 30052 26794
rect 30392 26382 30420 26846
rect 30748 26794 30800 26800
rect 30472 26784 30524 26790
rect 30472 26726 30524 26732
rect 30656 26784 30708 26790
rect 30656 26726 30708 26732
rect 30380 26376 30432 26382
rect 30380 26318 30432 26324
rect 30484 26246 30512 26726
rect 30668 26382 30696 26726
rect 30656 26376 30708 26382
rect 30656 26318 30708 26324
rect 31024 26376 31076 26382
rect 31024 26318 31076 26324
rect 30012 26240 30064 26246
rect 30012 26182 30064 26188
rect 30472 26240 30524 26246
rect 30472 26182 30524 26188
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 30012 17536 30064 17542
rect 30012 17478 30064 17484
rect 30840 17536 30892 17542
rect 30840 17478 30892 17484
rect 30024 17338 30052 17478
rect 30012 17332 30064 17338
rect 30012 17274 30064 17280
rect 30852 16590 30880 17478
rect 30840 16584 30892 16590
rect 30840 16526 30892 16532
rect 29736 16448 29788 16454
rect 29736 16390 29788 16396
rect 30656 16448 30708 16454
rect 30656 16390 30708 16396
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29564 12306 29592 15438
rect 29644 14408 29696 14414
rect 29644 14350 29696 14356
rect 29656 14074 29684 14350
rect 29644 14068 29696 14074
rect 29644 14010 29696 14016
rect 29642 13288 29698 13297
rect 29642 13223 29644 13232
rect 29696 13223 29698 13232
rect 29644 13194 29696 13200
rect 29552 12300 29604 12306
rect 29552 12242 29604 12248
rect 29550 12064 29606 12073
rect 29550 11999 29606 12008
rect 29564 11286 29592 11999
rect 29552 11280 29604 11286
rect 29552 11222 29604 11228
rect 29460 11212 29512 11218
rect 29460 11154 29512 11160
rect 29472 5370 29500 11154
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29564 10606 29592 11086
rect 29748 10985 29776 16390
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 30116 15026 30144 16050
rect 30196 15428 30248 15434
rect 30196 15370 30248 15376
rect 30104 15020 30156 15026
rect 30104 14962 30156 14968
rect 30012 14272 30064 14278
rect 30012 14214 30064 14220
rect 29828 13796 29880 13802
rect 29828 13738 29880 13744
rect 29840 13190 29868 13738
rect 29828 13184 29880 13190
rect 29828 13126 29880 13132
rect 30024 12646 30052 14214
rect 30116 13938 30144 14962
rect 30208 14414 30236 15370
rect 30286 14920 30342 14929
rect 30286 14855 30342 14864
rect 30196 14408 30248 14414
rect 30196 14350 30248 14356
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 30116 13326 30144 13874
rect 30300 13530 30328 14855
rect 30484 14482 30512 16118
rect 30562 15872 30618 15881
rect 30562 15807 30618 15816
rect 30576 15638 30604 15807
rect 30564 15632 30616 15638
rect 30564 15574 30616 15580
rect 30668 15434 30696 16390
rect 30760 16250 30788 16390
rect 30748 16244 30800 16250
rect 30748 16186 30800 16192
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 30656 15428 30708 15434
rect 30656 15370 30708 15376
rect 30852 14822 30880 16118
rect 30840 14816 30892 14822
rect 30840 14758 30892 14764
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 30748 14340 30800 14346
rect 30748 14282 30800 14288
rect 30760 13734 30788 14282
rect 30838 14240 30894 14249
rect 30838 14175 30894 14184
rect 30852 14006 30880 14175
rect 30840 14000 30892 14006
rect 30840 13942 30892 13948
rect 30472 13728 30524 13734
rect 30472 13670 30524 13676
rect 30748 13728 30800 13734
rect 30748 13670 30800 13676
rect 30484 13530 30512 13670
rect 30288 13524 30340 13530
rect 30288 13466 30340 13472
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30852 13326 30880 13942
rect 30944 13841 30972 20402
rect 30930 13832 30986 13841
rect 30930 13767 30986 13776
rect 30944 13394 30972 13767
rect 30932 13388 30984 13394
rect 30932 13330 30984 13336
rect 30104 13320 30156 13326
rect 30104 13262 30156 13268
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30012 12640 30064 12646
rect 30012 12582 30064 12588
rect 30024 12209 30052 12582
rect 30010 12200 30066 12209
rect 30010 12135 30066 12144
rect 29826 11928 29882 11937
rect 30116 11898 30144 13262
rect 30380 13252 30432 13258
rect 30380 13194 30432 13200
rect 30392 12850 30420 13194
rect 30656 13184 30708 13190
rect 30656 13126 30708 13132
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 29826 11863 29882 11872
rect 30012 11892 30064 11898
rect 29840 11830 29868 11863
rect 30012 11834 30064 11840
rect 30104 11892 30156 11898
rect 30104 11834 30156 11840
rect 29828 11824 29880 11830
rect 29828 11766 29880 11772
rect 29828 11688 29880 11694
rect 29828 11630 29880 11636
rect 29734 10976 29790 10985
rect 29734 10911 29790 10920
rect 29748 10810 29776 10911
rect 29736 10804 29788 10810
rect 29736 10746 29788 10752
rect 29840 10742 29868 11630
rect 30024 11014 30052 11834
rect 30012 11008 30064 11014
rect 30012 10950 30064 10956
rect 29828 10736 29880 10742
rect 29828 10678 29880 10684
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29564 10062 29592 10542
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29368 5364 29420 5370
rect 29368 5306 29420 5312
rect 29460 5364 29512 5370
rect 29460 5306 29512 5312
rect 29380 4690 29408 5306
rect 29368 4684 29420 4690
rect 29368 4626 29420 4632
rect 29184 4004 29236 4010
rect 29184 3946 29236 3952
rect 29196 3738 29224 3946
rect 29184 3732 29236 3738
rect 29184 3674 29236 3680
rect 29184 2916 29236 2922
rect 29184 2858 29236 2864
rect 29196 2310 29224 2858
rect 29472 2854 29500 5306
rect 30024 3466 30052 10950
rect 30288 10736 30340 10742
rect 30288 10678 30340 10684
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30116 9674 30144 10406
rect 30300 9722 30328 10678
rect 30288 9716 30340 9722
rect 30116 9646 30236 9674
rect 30288 9658 30340 9664
rect 30208 9518 30236 9646
rect 30300 9518 30328 9658
rect 30196 9512 30248 9518
rect 30196 9454 30248 9460
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 30012 3460 30064 3466
rect 30012 3402 30064 3408
rect 29460 2848 29512 2854
rect 29460 2790 29512 2796
rect 29920 2644 29972 2650
rect 29920 2586 29972 2592
rect 29932 2446 29960 2586
rect 29920 2440 29972 2446
rect 29920 2382 29972 2388
rect 29184 2304 29236 2310
rect 29184 2246 29236 2252
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 29092 1352 29144 1358
rect 29092 1294 29144 1300
rect 29656 800 29684 2246
rect 30208 1562 30236 9454
rect 30668 5302 30696 13126
rect 30932 12844 30984 12850
rect 30932 12786 30984 12792
rect 30944 12442 30972 12786
rect 30932 12436 30984 12442
rect 30932 12378 30984 12384
rect 30840 11756 30892 11762
rect 30840 11698 30892 11704
rect 30748 11144 30800 11150
rect 30746 11112 30748 11121
rect 30800 11112 30802 11121
rect 30746 11047 30802 11056
rect 30748 10804 30800 10810
rect 30748 10746 30800 10752
rect 30656 5296 30708 5302
rect 30656 5238 30708 5244
rect 30668 4214 30696 5238
rect 30656 4208 30708 4214
rect 30656 4150 30708 4156
rect 30760 3534 30788 10746
rect 30852 3738 30880 11698
rect 31036 11286 31064 26318
rect 31128 22681 31156 27406
rect 31206 27367 31262 27376
rect 31114 22672 31170 22681
rect 31114 22607 31170 22616
rect 31220 17746 31248 27367
rect 31312 26382 31340 27610
rect 31680 27554 31708 29294
rect 32862 29294 32996 29322
rect 32862 29200 32918 29294
rect 31576 27532 31628 27538
rect 31680 27526 31892 27554
rect 31576 27474 31628 27480
rect 31300 26376 31352 26382
rect 31300 26318 31352 26324
rect 31392 19372 31444 19378
rect 31392 19314 31444 19320
rect 31116 17740 31168 17746
rect 31116 17682 31168 17688
rect 31208 17740 31260 17746
rect 31208 17682 31260 17688
rect 31128 17513 31156 17682
rect 31114 17504 31170 17513
rect 31114 17439 31170 17448
rect 31116 16584 31168 16590
rect 31116 16526 31168 16532
rect 31128 15502 31156 16526
rect 31116 15496 31168 15502
rect 31116 15438 31168 15444
rect 31404 15144 31432 19314
rect 31484 16992 31536 16998
rect 31484 16934 31536 16940
rect 31496 16522 31524 16934
rect 31484 16516 31536 16522
rect 31484 16458 31536 16464
rect 31588 16182 31616 27474
rect 31864 27470 31892 27526
rect 32680 27532 32732 27538
rect 32680 27474 32732 27480
rect 31852 27464 31904 27470
rect 31852 27406 31904 27412
rect 31944 27396 31996 27402
rect 31944 27338 31996 27344
rect 31956 26602 31984 27338
rect 32692 27062 32720 27474
rect 32968 27130 32996 29294
rect 33506 29200 33562 30000
rect 34150 29322 34206 30000
rect 34794 29322 34850 30000
rect 35438 29322 35494 30000
rect 34150 29294 34284 29322
rect 34150 29200 34206 29294
rect 33520 27606 33548 29200
rect 33872 27772 34180 27781
rect 33872 27770 33878 27772
rect 33934 27770 33958 27772
rect 34014 27770 34038 27772
rect 34094 27770 34118 27772
rect 34174 27770 34180 27772
rect 33934 27718 33936 27770
rect 34116 27718 34118 27770
rect 33872 27716 33878 27718
rect 33934 27716 33958 27718
rect 34014 27716 34038 27718
rect 34094 27716 34118 27718
rect 34174 27716 34180 27718
rect 33872 27707 34180 27716
rect 34256 27606 34284 29294
rect 34794 29294 34928 29322
rect 34794 29200 34850 29294
rect 34900 27606 34928 29294
rect 35438 29294 35572 29322
rect 35438 29200 35494 29294
rect 35544 27606 35572 29294
rect 36082 29200 36138 30000
rect 36726 29322 36782 30000
rect 37370 29322 37426 30000
rect 38014 29322 38070 30000
rect 38658 29322 38714 30000
rect 36726 29294 36860 29322
rect 36726 29200 36782 29294
rect 36096 27606 36124 29200
rect 36544 27668 36596 27674
rect 36544 27610 36596 27616
rect 33508 27600 33560 27606
rect 33508 27542 33560 27548
rect 34244 27600 34296 27606
rect 34244 27542 34296 27548
rect 34888 27600 34940 27606
rect 34888 27542 34940 27548
rect 35532 27600 35584 27606
rect 35532 27542 35584 27548
rect 36084 27600 36136 27606
rect 36084 27542 36136 27548
rect 36176 27600 36228 27606
rect 36176 27542 36228 27548
rect 33692 27464 33744 27470
rect 33692 27406 33744 27412
rect 34244 27464 34296 27470
rect 34244 27406 34296 27412
rect 35072 27464 35124 27470
rect 35072 27406 35124 27412
rect 35716 27464 35768 27470
rect 35716 27406 35768 27412
rect 32956 27124 33008 27130
rect 32956 27066 33008 27072
rect 33048 27124 33100 27130
rect 33048 27066 33100 27072
rect 32680 27056 32732 27062
rect 32680 26998 32732 27004
rect 32864 26988 32916 26994
rect 32864 26930 32916 26936
rect 32876 26790 32904 26930
rect 32864 26784 32916 26790
rect 32864 26726 32916 26732
rect 31772 26574 31984 26602
rect 31772 26518 31800 26574
rect 31760 26512 31812 26518
rect 33060 26489 33088 27066
rect 33232 26988 33284 26994
rect 33232 26930 33284 26936
rect 31760 26454 31812 26460
rect 33046 26480 33102 26489
rect 33046 26415 33102 26424
rect 32220 26036 32272 26042
rect 32220 25978 32272 25984
rect 31944 17876 31996 17882
rect 31944 17818 31996 17824
rect 31760 17808 31812 17814
rect 31760 17750 31812 17756
rect 31772 17490 31800 17750
rect 31956 17610 31984 17818
rect 31944 17604 31996 17610
rect 31944 17546 31996 17552
rect 32128 17604 32180 17610
rect 32128 17546 32180 17552
rect 31772 17462 32076 17490
rect 31758 17368 31814 17377
rect 31758 17303 31814 17312
rect 31772 17134 31800 17303
rect 32048 17134 32076 17462
rect 32140 17270 32168 17546
rect 32232 17270 32260 25978
rect 32864 25764 32916 25770
rect 32864 25706 32916 25712
rect 32312 22976 32364 22982
rect 32312 22918 32364 22924
rect 32128 17264 32180 17270
rect 32128 17206 32180 17212
rect 32220 17264 32272 17270
rect 32220 17206 32272 17212
rect 31760 17128 31812 17134
rect 31760 17070 31812 17076
rect 32036 17128 32088 17134
rect 32036 17070 32088 17076
rect 31576 16176 31628 16182
rect 31576 16118 31628 16124
rect 31220 15116 31432 15144
rect 31482 15192 31538 15201
rect 31482 15127 31538 15136
rect 31116 14408 31168 14414
rect 31116 14350 31168 14356
rect 31128 13938 31156 14350
rect 31220 14278 31248 15116
rect 31300 15020 31352 15026
rect 31300 14962 31352 14968
rect 31312 14618 31340 14962
rect 31300 14612 31352 14618
rect 31300 14554 31352 14560
rect 31496 14550 31524 15127
rect 31772 14940 31800 17070
rect 32128 16040 32180 16046
rect 32128 15982 32180 15988
rect 32220 16040 32272 16046
rect 32220 15982 32272 15988
rect 31944 15972 31996 15978
rect 31944 15914 31996 15920
rect 31956 15609 31984 15914
rect 31942 15600 31998 15609
rect 31942 15535 31998 15544
rect 32036 15496 32088 15502
rect 32036 15438 32088 15444
rect 31944 15156 31996 15162
rect 31944 15098 31996 15104
rect 31772 14912 31892 14940
rect 31864 14822 31892 14912
rect 31760 14816 31812 14822
rect 31760 14758 31812 14764
rect 31852 14816 31904 14822
rect 31852 14758 31904 14764
rect 31484 14544 31536 14550
rect 31484 14486 31536 14492
rect 31208 14272 31260 14278
rect 31260 14232 31340 14260
rect 31208 14214 31260 14220
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 31114 13832 31170 13841
rect 31114 13767 31116 13776
rect 31168 13767 31170 13776
rect 31116 13738 31168 13744
rect 31312 13546 31340 14232
rect 31496 14006 31524 14486
rect 31668 14476 31720 14482
rect 31668 14418 31720 14424
rect 31576 14340 31628 14346
rect 31576 14282 31628 14288
rect 31484 14000 31536 14006
rect 31484 13942 31536 13948
rect 31312 13518 31432 13546
rect 31300 13388 31352 13394
rect 31300 13330 31352 13336
rect 31116 11824 31168 11830
rect 31116 11766 31168 11772
rect 31128 11626 31156 11766
rect 31116 11620 31168 11626
rect 31116 11562 31168 11568
rect 31024 11280 31076 11286
rect 31024 11222 31076 11228
rect 31116 10464 31168 10470
rect 31116 10406 31168 10412
rect 31128 9586 31156 10406
rect 31116 9580 31168 9586
rect 31116 9522 31168 9528
rect 31128 8906 31156 9522
rect 31116 8900 31168 8906
rect 31116 8842 31168 8848
rect 31208 4208 31260 4214
rect 31208 4150 31260 4156
rect 30840 3732 30892 3738
rect 30840 3674 30892 3680
rect 31220 3534 31248 4150
rect 30748 3528 30800 3534
rect 30748 3470 30800 3476
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31312 3466 31340 13330
rect 31404 6730 31432 13518
rect 31588 12442 31616 14282
rect 31680 14006 31708 14418
rect 31668 14000 31720 14006
rect 31668 13942 31720 13948
rect 31668 13320 31720 13326
rect 31668 13262 31720 13268
rect 31576 12436 31628 12442
rect 31576 12378 31628 12384
rect 31484 11756 31536 11762
rect 31484 11698 31536 11704
rect 31496 10849 31524 11698
rect 31680 11626 31708 13262
rect 31772 12238 31800 14758
rect 31956 14618 31984 15098
rect 31852 14612 31904 14618
rect 31852 14554 31904 14560
rect 31944 14612 31996 14618
rect 31944 14554 31996 14560
rect 31864 14521 31892 14554
rect 31850 14512 31906 14521
rect 32048 14482 32076 15438
rect 32140 15162 32168 15982
rect 32232 15706 32260 15982
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32324 15162 32352 22918
rect 32404 17740 32456 17746
rect 32404 17682 32456 17688
rect 32416 17134 32444 17682
rect 32496 17536 32548 17542
rect 32496 17478 32548 17484
rect 32770 17504 32826 17513
rect 32404 17128 32456 17134
rect 32404 17070 32456 17076
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32128 15156 32180 15162
rect 32128 15098 32180 15104
rect 32312 15156 32364 15162
rect 32312 15098 32364 15104
rect 32416 15042 32444 16050
rect 32508 15706 32536 17478
rect 32770 17439 32826 17448
rect 32784 17270 32812 17439
rect 32772 17264 32824 17270
rect 32772 17206 32824 17212
rect 32680 17196 32732 17202
rect 32680 17138 32732 17144
rect 32692 16454 32720 17138
rect 32772 17128 32824 17134
rect 32772 17070 32824 17076
rect 32784 16726 32812 17070
rect 32772 16720 32824 16726
rect 32772 16662 32824 16668
rect 32876 16658 32904 25706
rect 33048 17060 33100 17066
rect 33048 17002 33100 17008
rect 32864 16652 32916 16658
rect 32864 16594 32916 16600
rect 32864 16516 32916 16522
rect 32864 16458 32916 16464
rect 32680 16448 32732 16454
rect 32680 16390 32732 16396
rect 32496 15700 32548 15706
rect 32548 15660 32628 15688
rect 32496 15642 32548 15648
rect 32494 15600 32550 15609
rect 32494 15535 32550 15544
rect 32508 15502 32536 15535
rect 32496 15496 32548 15502
rect 32496 15438 32548 15444
rect 32496 15360 32548 15366
rect 32496 15302 32548 15308
rect 32508 15094 32536 15302
rect 32324 15014 32444 15042
rect 32496 15088 32548 15094
rect 32496 15030 32548 15036
rect 32600 15026 32628 15660
rect 32692 15094 32720 16390
rect 32876 16114 32904 16458
rect 33060 16114 33088 17002
rect 33140 16448 33192 16454
rect 33140 16390 33192 16396
rect 33152 16182 33180 16390
rect 33140 16176 33192 16182
rect 33140 16118 33192 16124
rect 32864 16108 32916 16114
rect 33048 16108 33100 16114
rect 32916 16068 32996 16096
rect 32864 16050 32916 16056
rect 32864 15972 32916 15978
rect 32864 15914 32916 15920
rect 32680 15088 32732 15094
rect 32680 15030 32732 15036
rect 32588 15020 32640 15026
rect 32128 14816 32180 14822
rect 32128 14758 32180 14764
rect 31850 14447 31906 14456
rect 32036 14476 32088 14482
rect 32036 14418 32088 14424
rect 31852 14408 31904 14414
rect 31852 14350 31904 14356
rect 31864 13394 31892 14350
rect 31944 13524 31996 13530
rect 31944 13466 31996 13472
rect 31852 13388 31904 13394
rect 31852 13330 31904 13336
rect 31956 12850 31984 13466
rect 31944 12844 31996 12850
rect 31944 12786 31996 12792
rect 32036 12844 32088 12850
rect 32036 12786 32088 12792
rect 32048 12646 32076 12786
rect 32036 12640 32088 12646
rect 32036 12582 32088 12588
rect 32140 12374 32168 14758
rect 32324 14006 32352 15014
rect 32588 14962 32640 14968
rect 32402 14784 32458 14793
rect 32402 14719 32458 14728
rect 32312 14000 32364 14006
rect 32312 13942 32364 13948
rect 32324 13326 32352 13942
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 32416 12850 32444 14719
rect 32772 14408 32824 14414
rect 32772 14350 32824 14356
rect 32496 13932 32548 13938
rect 32496 13874 32548 13880
rect 32508 12918 32536 13874
rect 32588 13456 32640 13462
rect 32588 13398 32640 13404
rect 32496 12912 32548 12918
rect 32496 12854 32548 12860
rect 32600 12850 32628 13398
rect 32784 13394 32812 14350
rect 32876 13705 32904 15914
rect 32862 13696 32918 13705
rect 32862 13631 32918 13640
rect 32772 13388 32824 13394
rect 32772 13330 32824 13336
rect 32680 13252 32732 13258
rect 32680 13194 32732 13200
rect 32404 12844 32456 12850
rect 32404 12786 32456 12792
rect 32588 12844 32640 12850
rect 32588 12786 32640 12792
rect 32220 12640 32272 12646
rect 32220 12582 32272 12588
rect 32232 12434 32260 12582
rect 32232 12406 32352 12434
rect 32128 12368 32180 12374
rect 32128 12310 32180 12316
rect 32220 12300 32272 12306
rect 32220 12242 32272 12248
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 32232 12102 32260 12242
rect 32220 12096 32272 12102
rect 32220 12038 32272 12044
rect 31758 11792 31814 11801
rect 31758 11727 31814 11736
rect 31668 11620 31720 11626
rect 31668 11562 31720 11568
rect 31772 11150 31800 11727
rect 31760 11144 31812 11150
rect 31760 11086 31812 11092
rect 31482 10840 31538 10849
rect 31482 10775 31484 10784
rect 31536 10775 31538 10784
rect 31484 10746 31536 10752
rect 31496 10715 31524 10746
rect 32324 10470 32352 12406
rect 32588 11552 32640 11558
rect 32588 11494 32640 11500
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32508 10742 32536 11086
rect 32496 10736 32548 10742
rect 32496 10678 32548 10684
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 32600 10282 32628 11494
rect 32508 10266 32628 10282
rect 32496 10260 32628 10266
rect 32548 10254 32628 10260
rect 32496 10202 32548 10208
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31392 6724 31444 6730
rect 31392 6666 31444 6672
rect 31576 6180 31628 6186
rect 31576 6122 31628 6128
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 31484 3732 31536 3738
rect 31484 3674 31536 3680
rect 31404 3534 31432 3674
rect 31392 3528 31444 3534
rect 31392 3470 31444 3476
rect 30288 3460 30340 3466
rect 30288 3402 30340 3408
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 30300 2009 30328 3402
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30392 2650 30420 2790
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 31116 2644 31168 2650
rect 31116 2586 31168 2592
rect 31128 2378 31156 2586
rect 31116 2372 31168 2378
rect 31116 2314 31168 2320
rect 31300 2372 31352 2378
rect 31300 2314 31352 2320
rect 30286 2000 30342 2009
rect 30286 1935 30342 1944
rect 30196 1556 30248 1562
rect 30196 1498 30248 1504
rect 30288 1556 30340 1562
rect 30288 1498 30340 1504
rect 30300 1426 30328 1498
rect 30288 1420 30340 1426
rect 30288 1362 30340 1368
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 31312 762 31340 2314
rect 31404 1834 31432 3470
rect 31496 3398 31524 3674
rect 31484 3392 31536 3398
rect 31484 3334 31536 3340
rect 31484 2848 31536 2854
rect 31484 2790 31536 2796
rect 31496 2446 31524 2790
rect 31588 2514 31616 6122
rect 31668 3392 31720 3398
rect 31668 3334 31720 3340
rect 31680 3058 31708 3334
rect 31772 3126 31800 9998
rect 32600 9722 32628 10254
rect 32588 9716 32640 9722
rect 32588 9658 32640 9664
rect 31852 4820 31904 4826
rect 31852 4762 31904 4768
rect 31760 3120 31812 3126
rect 31760 3062 31812 3068
rect 31668 3052 31720 3058
rect 31668 2994 31720 3000
rect 31864 2774 31892 4762
rect 32588 3392 32640 3398
rect 32588 3334 32640 3340
rect 32600 3058 32628 3334
rect 32588 3052 32640 3058
rect 32588 2994 32640 3000
rect 31772 2746 31892 2774
rect 31668 2576 31720 2582
rect 31772 2530 31800 2746
rect 31720 2524 31800 2530
rect 31668 2518 31800 2524
rect 31852 2576 31904 2582
rect 31852 2518 31904 2524
rect 31576 2508 31628 2514
rect 31680 2502 31800 2518
rect 31576 2450 31628 2456
rect 31484 2440 31536 2446
rect 31484 2382 31536 2388
rect 31864 2009 31892 2518
rect 32692 2378 32720 13194
rect 32784 12850 32812 13330
rect 32772 12844 32824 12850
rect 32772 12786 32824 12792
rect 32876 12782 32904 13631
rect 32968 13462 32996 16068
rect 33048 16050 33100 16056
rect 33060 15706 33088 16050
rect 33140 16040 33192 16046
rect 33140 15982 33192 15988
rect 33152 15881 33180 15982
rect 33138 15872 33194 15881
rect 33138 15807 33194 15816
rect 33048 15700 33100 15706
rect 33048 15642 33100 15648
rect 33060 13462 33088 15642
rect 33152 13938 33180 15807
rect 33244 15162 33272 26930
rect 33416 26920 33468 26926
rect 33416 26862 33468 26868
rect 33324 16584 33376 16590
rect 33324 16526 33376 16532
rect 33336 15978 33364 16526
rect 33324 15972 33376 15978
rect 33324 15914 33376 15920
rect 33232 15156 33284 15162
rect 33232 15098 33284 15104
rect 33324 15156 33376 15162
rect 33324 15098 33376 15104
rect 33336 14929 33364 15098
rect 33322 14920 33378 14929
rect 33322 14855 33378 14864
rect 33232 14816 33284 14822
rect 33232 14758 33284 14764
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 32956 13456 33008 13462
rect 32956 13398 33008 13404
rect 33048 13456 33100 13462
rect 33048 13398 33100 13404
rect 32968 13190 32996 13398
rect 32956 13184 33008 13190
rect 32956 13126 33008 13132
rect 33140 12844 33192 12850
rect 33060 12804 33140 12832
rect 32864 12776 32916 12782
rect 32864 12718 32916 12724
rect 32956 12640 33008 12646
rect 32956 12582 33008 12588
rect 32864 12368 32916 12374
rect 32864 12310 32916 12316
rect 32876 12170 32904 12310
rect 32864 12164 32916 12170
rect 32864 12106 32916 12112
rect 32968 12102 32996 12582
rect 33060 12442 33088 12804
rect 33140 12786 33192 12792
rect 33048 12436 33100 12442
rect 33048 12378 33100 12384
rect 33060 12238 33088 12378
rect 33244 12345 33272 14758
rect 33322 14240 33378 14249
rect 33322 14175 33378 14184
rect 33336 13802 33364 14175
rect 33428 14006 33456 26862
rect 33704 25770 33732 27406
rect 33872 26684 34180 26693
rect 33872 26682 33878 26684
rect 33934 26682 33958 26684
rect 34014 26682 34038 26684
rect 34094 26682 34118 26684
rect 34174 26682 34180 26684
rect 33934 26630 33936 26682
rect 34116 26630 34118 26682
rect 33872 26628 33878 26630
rect 33934 26628 33958 26630
rect 34014 26628 34038 26630
rect 34094 26628 34118 26630
rect 34174 26628 34180 26630
rect 33872 26619 34180 26628
rect 33692 25764 33744 25770
rect 33692 25706 33744 25712
rect 33872 25596 34180 25605
rect 33872 25594 33878 25596
rect 33934 25594 33958 25596
rect 34014 25594 34038 25596
rect 34094 25594 34118 25596
rect 34174 25594 34180 25596
rect 33934 25542 33936 25594
rect 34116 25542 34118 25594
rect 33872 25540 33878 25542
rect 33934 25540 33958 25542
rect 34014 25540 34038 25542
rect 34094 25540 34118 25542
rect 34174 25540 34180 25542
rect 33872 25531 34180 25540
rect 33872 24508 34180 24517
rect 33872 24506 33878 24508
rect 33934 24506 33958 24508
rect 34014 24506 34038 24508
rect 34094 24506 34118 24508
rect 34174 24506 34180 24508
rect 33934 24454 33936 24506
rect 34116 24454 34118 24506
rect 33872 24452 33878 24454
rect 33934 24452 33958 24454
rect 34014 24452 34038 24454
rect 34094 24452 34118 24454
rect 34174 24452 34180 24454
rect 33872 24443 34180 24452
rect 33872 23420 34180 23429
rect 33872 23418 33878 23420
rect 33934 23418 33958 23420
rect 34014 23418 34038 23420
rect 34094 23418 34118 23420
rect 34174 23418 34180 23420
rect 33934 23366 33936 23418
rect 34116 23366 34118 23418
rect 33872 23364 33878 23366
rect 33934 23364 33958 23366
rect 34014 23364 34038 23366
rect 34094 23364 34118 23366
rect 34174 23364 34180 23366
rect 33872 23355 34180 23364
rect 33872 22332 34180 22341
rect 33872 22330 33878 22332
rect 33934 22330 33958 22332
rect 34014 22330 34038 22332
rect 34094 22330 34118 22332
rect 34174 22330 34180 22332
rect 33934 22278 33936 22330
rect 34116 22278 34118 22330
rect 33872 22276 33878 22278
rect 33934 22276 33958 22278
rect 34014 22276 34038 22278
rect 34094 22276 34118 22278
rect 34174 22276 34180 22278
rect 33872 22267 34180 22276
rect 33872 21244 34180 21253
rect 33872 21242 33878 21244
rect 33934 21242 33958 21244
rect 34014 21242 34038 21244
rect 34094 21242 34118 21244
rect 34174 21242 34180 21244
rect 33934 21190 33936 21242
rect 34116 21190 34118 21242
rect 33872 21188 33878 21190
rect 33934 21188 33958 21190
rect 34014 21188 34038 21190
rect 34094 21188 34118 21190
rect 34174 21188 34180 21190
rect 33872 21179 34180 21188
rect 33872 20156 34180 20165
rect 33872 20154 33878 20156
rect 33934 20154 33958 20156
rect 34014 20154 34038 20156
rect 34094 20154 34118 20156
rect 34174 20154 34180 20156
rect 33934 20102 33936 20154
rect 34116 20102 34118 20154
rect 33872 20100 33878 20102
rect 33934 20100 33958 20102
rect 34014 20100 34038 20102
rect 34094 20100 34118 20102
rect 34174 20100 34180 20102
rect 33872 20091 34180 20100
rect 33872 19068 34180 19077
rect 33872 19066 33878 19068
rect 33934 19066 33958 19068
rect 34014 19066 34038 19068
rect 34094 19066 34118 19068
rect 34174 19066 34180 19068
rect 33934 19014 33936 19066
rect 34116 19014 34118 19066
rect 33872 19012 33878 19014
rect 33934 19012 33958 19014
rect 34014 19012 34038 19014
rect 34094 19012 34118 19014
rect 34174 19012 34180 19014
rect 33872 19003 34180 19012
rect 33692 18964 33744 18970
rect 33692 18906 33744 18912
rect 33600 17672 33652 17678
rect 33600 17614 33652 17620
rect 33612 17241 33640 17614
rect 33598 17232 33654 17241
rect 33598 17167 33600 17176
rect 33652 17167 33654 17176
rect 33600 17138 33652 17144
rect 33598 15736 33654 15745
rect 33598 15671 33654 15680
rect 33612 15026 33640 15671
rect 33508 15020 33560 15026
rect 33508 14962 33560 14968
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 33520 14793 33548 14962
rect 33506 14784 33562 14793
rect 33506 14719 33562 14728
rect 33704 14090 33732 18906
rect 33872 17980 34180 17989
rect 33872 17978 33878 17980
rect 33934 17978 33958 17980
rect 34014 17978 34038 17980
rect 34094 17978 34118 17980
rect 34174 17978 34180 17980
rect 33934 17926 33936 17978
rect 34116 17926 34118 17978
rect 33872 17924 33878 17926
rect 33934 17924 33958 17926
rect 34014 17924 34038 17926
rect 34094 17924 34118 17926
rect 34174 17924 34180 17926
rect 33872 17915 34180 17924
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 33796 17202 33824 17478
rect 33784 17196 33836 17202
rect 33784 17138 33836 17144
rect 33796 16658 33824 17138
rect 33872 16892 34180 16901
rect 33872 16890 33878 16892
rect 33934 16890 33958 16892
rect 34014 16890 34038 16892
rect 34094 16890 34118 16892
rect 34174 16890 34180 16892
rect 33934 16838 33936 16890
rect 34116 16838 34118 16890
rect 33872 16836 33878 16838
rect 33934 16836 33958 16838
rect 34014 16836 34038 16838
rect 34094 16836 34118 16838
rect 34174 16836 34180 16838
rect 33872 16827 34180 16836
rect 33784 16652 33836 16658
rect 33784 16594 33836 16600
rect 34256 15910 34284 27406
rect 35084 22982 35112 27406
rect 35532 27056 35584 27062
rect 35532 26998 35584 27004
rect 35256 26988 35308 26994
rect 35256 26930 35308 26936
rect 35072 22976 35124 22982
rect 35072 22918 35124 22924
rect 34520 18964 34572 18970
rect 34520 18906 34572 18912
rect 34336 18896 34388 18902
rect 34336 18838 34388 18844
rect 34348 18290 34376 18838
rect 34336 18284 34388 18290
rect 34336 18226 34388 18232
rect 34532 18222 34560 18906
rect 34520 18216 34572 18222
rect 34520 18158 34572 18164
rect 34980 18080 35032 18086
rect 34980 18022 35032 18028
rect 34428 17672 34480 17678
rect 34428 17614 34480 17620
rect 34704 17672 34756 17678
rect 34704 17614 34756 17620
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34348 16561 34376 17070
rect 34334 16552 34390 16561
rect 34334 16487 34390 16496
rect 34244 15904 34296 15910
rect 34244 15846 34296 15852
rect 33872 15804 34180 15813
rect 33872 15802 33878 15804
rect 33934 15802 33958 15804
rect 34014 15802 34038 15804
rect 34094 15802 34118 15804
rect 34174 15802 34180 15804
rect 33934 15750 33936 15802
rect 34116 15750 34118 15802
rect 33872 15748 33878 15750
rect 33934 15748 33958 15750
rect 34014 15748 34038 15750
rect 34094 15748 34118 15750
rect 34174 15748 34180 15750
rect 33872 15739 34180 15748
rect 34440 15706 34468 17614
rect 34716 17066 34744 17614
rect 34992 17610 35020 18022
rect 34796 17604 34848 17610
rect 34796 17546 34848 17552
rect 34980 17604 35032 17610
rect 34980 17546 35032 17552
rect 34808 17490 34836 17546
rect 35164 17536 35216 17542
rect 34808 17484 35164 17490
rect 34808 17478 35216 17484
rect 34808 17462 35204 17478
rect 35070 17232 35126 17241
rect 35070 17167 35126 17176
rect 34704 17060 34756 17066
rect 34704 17002 34756 17008
rect 34704 16516 34756 16522
rect 34704 16458 34756 16464
rect 34716 16250 34744 16458
rect 34704 16244 34756 16250
rect 34704 16186 34756 16192
rect 34428 15700 34480 15706
rect 34428 15642 34480 15648
rect 34244 15088 34296 15094
rect 34244 15030 34296 15036
rect 33968 15020 34020 15026
rect 33968 14962 34020 14968
rect 33980 14929 34008 14962
rect 33966 14920 34022 14929
rect 33966 14855 34022 14864
rect 33872 14716 34180 14725
rect 33872 14714 33878 14716
rect 33934 14714 33958 14716
rect 34014 14714 34038 14716
rect 34094 14714 34118 14716
rect 34174 14714 34180 14716
rect 33934 14662 33936 14714
rect 34116 14662 34118 14714
rect 33872 14660 33878 14662
rect 33934 14660 33958 14662
rect 34014 14660 34038 14662
rect 34094 14660 34118 14662
rect 34174 14660 34180 14662
rect 33872 14651 34180 14660
rect 34256 14600 34284 15030
rect 34164 14572 34284 14600
rect 33876 14408 33928 14414
rect 33876 14350 33928 14356
rect 33888 14113 33916 14350
rect 34164 14278 34192 14572
rect 34242 14512 34298 14521
rect 34242 14447 34298 14456
rect 34256 14346 34284 14447
rect 34440 14362 34468 15642
rect 35084 15502 35112 17167
rect 35072 15496 35124 15502
rect 35072 15438 35124 15444
rect 35268 15144 35296 26930
rect 35348 26512 35400 26518
rect 35348 26454 35400 26460
rect 35360 25838 35388 26454
rect 35544 26450 35572 26998
rect 35532 26444 35584 26450
rect 35532 26386 35584 26392
rect 35348 25832 35400 25838
rect 35348 25774 35400 25780
rect 35728 24206 35756 27406
rect 36188 27402 36216 27542
rect 36176 27396 36228 27402
rect 36176 27338 36228 27344
rect 35716 24200 35768 24206
rect 35716 24142 35768 24148
rect 36360 22772 36412 22778
rect 36360 22714 36412 22720
rect 36176 22636 36228 22642
rect 36176 22578 36228 22584
rect 35992 18760 36044 18766
rect 35992 18702 36044 18708
rect 35716 18624 35768 18630
rect 35716 18566 35768 18572
rect 35728 17270 35756 18566
rect 36004 18426 36032 18702
rect 35992 18420 36044 18426
rect 35992 18362 36044 18368
rect 35992 18284 36044 18290
rect 35992 18226 36044 18232
rect 35716 17264 35768 17270
rect 35716 17206 35768 17212
rect 35440 17128 35492 17134
rect 35440 17070 35492 17076
rect 35348 15972 35400 15978
rect 35348 15914 35400 15920
rect 35360 15502 35388 15914
rect 35452 15638 35480 17070
rect 35900 16584 35952 16590
rect 35900 16526 35952 16532
rect 35532 16448 35584 16454
rect 35532 16390 35584 16396
rect 35440 15632 35492 15638
rect 35440 15574 35492 15580
rect 35348 15496 35400 15502
rect 35348 15438 35400 15444
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 35176 15116 35296 15144
rect 34520 14952 34572 14958
rect 34520 14894 34572 14900
rect 34532 14822 34560 14894
rect 34520 14816 34572 14822
rect 34520 14758 34572 14764
rect 34704 14816 34756 14822
rect 34704 14758 34756 14764
rect 34520 14544 34572 14550
rect 34520 14486 34572 14492
rect 34244 14340 34296 14346
rect 34244 14282 34296 14288
rect 34348 14334 34468 14362
rect 34152 14272 34204 14278
rect 34152 14214 34204 14220
rect 33520 14062 33732 14090
rect 33874 14104 33930 14113
rect 33416 14000 33468 14006
rect 33416 13942 33468 13948
rect 33414 13832 33470 13841
rect 33324 13796 33376 13802
rect 33414 13767 33416 13776
rect 33324 13738 33376 13744
rect 33468 13767 33470 13776
rect 33416 13738 33468 13744
rect 33520 12646 33548 14062
rect 33874 14039 33930 14048
rect 33692 14000 33744 14006
rect 33692 13942 33744 13948
rect 33600 13252 33652 13258
rect 33600 13194 33652 13200
rect 33612 12782 33640 13194
rect 33600 12776 33652 12782
rect 33600 12718 33652 12724
rect 33508 12640 33560 12646
rect 33428 12600 33508 12628
rect 33230 12336 33286 12345
rect 33230 12271 33286 12280
rect 33048 12232 33100 12238
rect 33048 12174 33100 12180
rect 33324 12232 33376 12238
rect 33324 12174 33376 12180
rect 32956 12096 33008 12102
rect 32956 12038 33008 12044
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 32876 11665 32904 11698
rect 32862 11656 32918 11665
rect 32862 11591 32918 11600
rect 32772 11552 32824 11558
rect 32772 11494 32824 11500
rect 32784 11014 32812 11494
rect 32772 11008 32824 11014
rect 32772 10950 32824 10956
rect 32968 4554 32996 12038
rect 33060 11830 33088 12174
rect 33336 12073 33364 12174
rect 33322 12064 33378 12073
rect 33322 11999 33378 12008
rect 33048 11824 33100 11830
rect 33048 11766 33100 11772
rect 33324 11688 33376 11694
rect 33244 11648 33324 11676
rect 33244 11082 33272 11648
rect 33324 11630 33376 11636
rect 33140 11076 33192 11082
rect 33140 11018 33192 11024
rect 33232 11076 33284 11082
rect 33232 11018 33284 11024
rect 33152 10810 33180 11018
rect 33140 10804 33192 10810
rect 33140 10746 33192 10752
rect 33244 10062 33272 11018
rect 33232 10056 33284 10062
rect 33232 9998 33284 10004
rect 32956 4548 33008 4554
rect 32956 4490 33008 4496
rect 33428 3584 33456 12600
rect 33508 12582 33560 12588
rect 33508 12300 33560 12306
rect 33508 12242 33560 12248
rect 33520 10674 33548 12242
rect 33600 11756 33652 11762
rect 33600 11698 33652 11704
rect 33612 10810 33640 11698
rect 33600 10804 33652 10810
rect 33600 10746 33652 10752
rect 33508 10668 33560 10674
rect 33508 10610 33560 10616
rect 33508 10260 33560 10266
rect 33508 10202 33560 10208
rect 33520 9654 33548 10202
rect 33508 9648 33560 9654
rect 33508 9590 33560 9596
rect 33704 8430 33732 13942
rect 33872 13628 34180 13637
rect 33872 13626 33878 13628
rect 33934 13626 33958 13628
rect 34014 13626 34038 13628
rect 34094 13626 34118 13628
rect 34174 13626 34180 13628
rect 33934 13574 33936 13626
rect 34116 13574 34118 13626
rect 33872 13572 33878 13574
rect 33934 13572 33958 13574
rect 34014 13572 34038 13574
rect 34094 13572 34118 13574
rect 34174 13572 34180 13574
rect 33872 13563 34180 13572
rect 33784 13320 33836 13326
rect 33784 13262 33836 13268
rect 34152 13320 34204 13326
rect 34152 13262 34204 13268
rect 33796 12238 33824 13262
rect 34164 13161 34192 13262
rect 34150 13152 34206 13161
rect 34150 13087 34206 13096
rect 33876 12980 33928 12986
rect 33876 12922 33928 12928
rect 33888 12646 33916 12922
rect 34244 12912 34296 12918
rect 34244 12854 34296 12860
rect 33876 12640 33928 12646
rect 33876 12582 33928 12588
rect 33872 12540 34180 12549
rect 33872 12538 33878 12540
rect 33934 12538 33958 12540
rect 34014 12538 34038 12540
rect 34094 12538 34118 12540
rect 34174 12538 34180 12540
rect 33934 12486 33936 12538
rect 34116 12486 34118 12538
rect 33872 12484 33878 12486
rect 33934 12484 33958 12486
rect 34014 12484 34038 12486
rect 34094 12484 34118 12486
rect 34174 12484 34180 12486
rect 33872 12475 34180 12484
rect 33784 12232 33836 12238
rect 33784 12174 33836 12180
rect 33874 11928 33930 11937
rect 33874 11863 33930 11872
rect 33888 11830 33916 11863
rect 33876 11824 33928 11830
rect 33876 11766 33928 11772
rect 33872 11452 34180 11461
rect 33872 11450 33878 11452
rect 33934 11450 33958 11452
rect 34014 11450 34038 11452
rect 34094 11450 34118 11452
rect 34174 11450 34180 11452
rect 33934 11398 33936 11450
rect 34116 11398 34118 11450
rect 33872 11396 33878 11398
rect 33934 11396 33958 11398
rect 34014 11396 34038 11398
rect 34094 11396 34118 11398
rect 34174 11396 34180 11398
rect 33872 11387 34180 11396
rect 34256 11354 34284 12854
rect 34348 12434 34376 14334
rect 34428 14272 34480 14278
rect 34428 14214 34480 14220
rect 34440 13938 34468 14214
rect 34428 13932 34480 13938
rect 34428 13874 34480 13880
rect 34428 13184 34480 13190
rect 34428 13126 34480 13132
rect 34440 12714 34468 13126
rect 34532 12850 34560 14486
rect 34716 14414 34744 14758
rect 35072 14544 35124 14550
rect 35072 14486 35124 14492
rect 34704 14408 34756 14414
rect 34980 14408 35032 14414
rect 34704 14350 34756 14356
rect 34978 14376 34980 14385
rect 35032 14376 35034 14385
rect 34888 14340 34940 14346
rect 34978 14311 35034 14320
rect 34888 14282 34940 14288
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34610 13560 34666 13569
rect 34610 13495 34612 13504
rect 34664 13495 34666 13504
rect 34612 13466 34664 13472
rect 34612 13388 34664 13394
rect 34664 13348 34744 13376
rect 34612 13330 34664 13336
rect 34612 13184 34664 13190
rect 34612 13126 34664 13132
rect 34624 12918 34652 13126
rect 34612 12912 34664 12918
rect 34612 12854 34664 12860
rect 34520 12844 34572 12850
rect 34716 12798 34744 13348
rect 34808 13326 34836 14010
rect 34900 13938 34928 14282
rect 34888 13932 34940 13938
rect 34888 13874 34940 13880
rect 34886 13696 34942 13705
rect 34886 13631 34942 13640
rect 34796 13320 34848 13326
rect 34796 13262 34848 13268
rect 34900 12850 34928 13631
rect 34888 12844 34940 12850
rect 34520 12786 34572 12792
rect 34624 12770 34744 12798
rect 34808 12804 34888 12832
rect 34428 12708 34480 12714
rect 34428 12650 34480 12656
rect 34440 12594 34468 12650
rect 34440 12566 34560 12594
rect 34532 12442 34560 12566
rect 34520 12436 34572 12442
rect 34348 12406 34468 12434
rect 34336 12300 34388 12306
rect 34336 12242 34388 12248
rect 34348 11801 34376 12242
rect 34334 11792 34390 11801
rect 34334 11727 34390 11736
rect 34244 11348 34296 11354
rect 34244 11290 34296 11296
rect 33876 10804 33928 10810
rect 33876 10746 33928 10752
rect 33784 10736 33836 10742
rect 33784 10678 33836 10684
rect 33796 10130 33824 10678
rect 33888 10470 33916 10746
rect 34244 10668 34296 10674
rect 34244 10610 34296 10616
rect 33876 10464 33928 10470
rect 33876 10406 33928 10412
rect 33872 10364 34180 10373
rect 33872 10362 33878 10364
rect 33934 10362 33958 10364
rect 34014 10362 34038 10364
rect 34094 10362 34118 10364
rect 34174 10362 34180 10364
rect 33934 10310 33936 10362
rect 34116 10310 34118 10362
rect 33872 10308 33878 10310
rect 33934 10308 33958 10310
rect 34014 10308 34038 10310
rect 34094 10308 34118 10310
rect 34174 10308 34180 10310
rect 33872 10299 34180 10308
rect 34256 10266 34284 10610
rect 34336 10464 34388 10470
rect 34336 10406 34388 10412
rect 34348 10266 34376 10406
rect 34244 10260 34296 10266
rect 34244 10202 34296 10208
rect 34336 10260 34388 10266
rect 34336 10202 34388 10208
rect 33784 10124 33836 10130
rect 33784 10066 33836 10072
rect 33784 9512 33836 9518
rect 33784 9454 33836 9460
rect 33796 9042 33824 9454
rect 33872 9276 34180 9285
rect 33872 9274 33878 9276
rect 33934 9274 33958 9276
rect 34014 9274 34038 9276
rect 34094 9274 34118 9276
rect 34174 9274 34180 9276
rect 33934 9222 33936 9274
rect 34116 9222 34118 9274
rect 33872 9220 33878 9222
rect 33934 9220 33958 9222
rect 34014 9220 34038 9222
rect 34094 9220 34118 9222
rect 34174 9220 34180 9222
rect 33872 9211 34180 9220
rect 33784 9036 33836 9042
rect 33784 8978 33836 8984
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 33872 8188 34180 8197
rect 33872 8186 33878 8188
rect 33934 8186 33958 8188
rect 34014 8186 34038 8188
rect 34094 8186 34118 8188
rect 34174 8186 34180 8188
rect 33934 8134 33936 8186
rect 34116 8134 34118 8186
rect 33872 8132 33878 8134
rect 33934 8132 33958 8134
rect 34014 8132 34038 8134
rect 34094 8132 34118 8134
rect 34174 8132 34180 8134
rect 33872 8123 34180 8132
rect 34440 7750 34468 12406
rect 34520 12378 34572 12384
rect 34624 12238 34652 12770
rect 34612 12232 34664 12238
rect 34612 12174 34664 12180
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34532 9722 34560 9998
rect 34612 9920 34664 9926
rect 34612 9862 34664 9868
rect 34520 9716 34572 9722
rect 34520 9658 34572 9664
rect 34624 9654 34652 9862
rect 34612 9648 34664 9654
rect 34612 9590 34664 9596
rect 34428 7744 34480 7750
rect 34428 7686 34480 7692
rect 33872 7100 34180 7109
rect 33872 7098 33878 7100
rect 33934 7098 33958 7100
rect 34014 7098 34038 7100
rect 34094 7098 34118 7100
rect 34174 7098 34180 7100
rect 33934 7046 33936 7098
rect 34116 7046 34118 7098
rect 33872 7044 33878 7046
rect 33934 7044 33958 7046
rect 34014 7044 34038 7046
rect 34094 7044 34118 7046
rect 34174 7044 34180 7046
rect 33872 7035 34180 7044
rect 34808 6186 34836 12804
rect 34888 12786 34940 12792
rect 34992 12102 35020 14311
rect 35084 13938 35112 14486
rect 35072 13932 35124 13938
rect 35072 13874 35124 13880
rect 35176 13802 35204 15116
rect 35256 15020 35308 15026
rect 35256 14962 35308 14968
rect 35268 14113 35296 14962
rect 35254 14104 35310 14113
rect 35254 14039 35310 14048
rect 35256 13932 35308 13938
rect 35256 13874 35308 13880
rect 35164 13796 35216 13802
rect 35164 13738 35216 13744
rect 35072 12640 35124 12646
rect 35072 12582 35124 12588
rect 34980 12096 35032 12102
rect 35084 12073 35112 12582
rect 35176 12102 35204 13738
rect 35268 12374 35296 13874
rect 35256 12368 35308 12374
rect 35256 12310 35308 12316
rect 35256 12164 35308 12170
rect 35256 12106 35308 12112
rect 35164 12096 35216 12102
rect 34980 12038 35032 12044
rect 35070 12064 35126 12073
rect 34992 11218 35020 12038
rect 35268 12073 35296 12106
rect 35164 12038 35216 12044
rect 35254 12064 35310 12073
rect 35070 11999 35126 12008
rect 35176 11914 35204 12038
rect 35254 11999 35310 12008
rect 35176 11886 35296 11914
rect 34980 11212 35032 11218
rect 34980 11154 35032 11160
rect 35072 11008 35124 11014
rect 35072 10950 35124 10956
rect 35164 11008 35216 11014
rect 35164 10950 35216 10956
rect 35084 10742 35112 10950
rect 35176 10810 35204 10950
rect 35164 10804 35216 10810
rect 35164 10746 35216 10752
rect 35072 10736 35124 10742
rect 35072 10678 35124 10684
rect 35164 10192 35216 10198
rect 35164 10134 35216 10140
rect 34888 10056 34940 10062
rect 34888 9998 34940 10004
rect 34900 9450 34928 9998
rect 35176 9586 35204 10134
rect 35164 9580 35216 9586
rect 35164 9522 35216 9528
rect 34888 9444 34940 9450
rect 34888 9386 34940 9392
rect 35268 6662 35296 11886
rect 35256 6656 35308 6662
rect 35256 6598 35308 6604
rect 34796 6180 34848 6186
rect 34796 6122 34848 6128
rect 33872 6012 34180 6021
rect 33872 6010 33878 6012
rect 33934 6010 33958 6012
rect 34014 6010 34038 6012
rect 34094 6010 34118 6012
rect 34174 6010 34180 6012
rect 33934 5958 33936 6010
rect 34116 5958 34118 6010
rect 33872 5956 33878 5958
rect 33934 5956 33958 5958
rect 34014 5956 34038 5958
rect 34094 5956 34118 5958
rect 34174 5956 34180 5958
rect 33872 5947 34180 5956
rect 33872 4924 34180 4933
rect 33872 4922 33878 4924
rect 33934 4922 33958 4924
rect 34014 4922 34038 4924
rect 34094 4922 34118 4924
rect 34174 4922 34180 4924
rect 33934 4870 33936 4922
rect 34116 4870 34118 4922
rect 33872 4868 33878 4870
rect 33934 4868 33958 4870
rect 34014 4868 34038 4870
rect 34094 4868 34118 4870
rect 34174 4868 34180 4870
rect 33872 4859 34180 4868
rect 33600 4548 33652 4554
rect 33600 4490 33652 4496
rect 33612 4214 33640 4490
rect 33600 4208 33652 4214
rect 33600 4150 33652 4156
rect 33872 3836 34180 3845
rect 33872 3834 33878 3836
rect 33934 3834 33958 3836
rect 34014 3834 34038 3836
rect 34094 3834 34118 3836
rect 34174 3834 34180 3836
rect 33934 3782 33936 3834
rect 34116 3782 34118 3834
rect 33872 3780 33878 3782
rect 33934 3780 33958 3782
rect 34014 3780 34038 3782
rect 34094 3780 34118 3782
rect 34174 3780 34180 3782
rect 33872 3771 34180 3780
rect 34704 3732 34756 3738
rect 34704 3674 34756 3680
rect 34888 3732 34940 3738
rect 34888 3674 34940 3680
rect 33508 3596 33560 3602
rect 33428 3556 33508 3584
rect 33508 3538 33560 3544
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33060 3398 33088 3470
rect 33968 3460 34020 3466
rect 33968 3402 34020 3408
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 33980 3126 34008 3402
rect 34716 3126 34744 3674
rect 33968 3120 34020 3126
rect 33968 3062 34020 3068
rect 34704 3120 34756 3126
rect 34704 3062 34756 3068
rect 34900 3058 34928 3674
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 33508 2916 33560 2922
rect 33508 2858 33560 2864
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32680 2372 32732 2378
rect 32680 2314 32732 2320
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 31850 2000 31906 2009
rect 31850 1935 31906 1944
rect 31668 1896 31720 1902
rect 31666 1864 31668 1873
rect 31720 1864 31722 1873
rect 31392 1828 31444 1834
rect 31666 1799 31722 1808
rect 31392 1770 31444 1776
rect 31758 1728 31814 1737
rect 31758 1663 31814 1672
rect 31772 1562 31800 1663
rect 31850 1592 31906 1601
rect 31760 1556 31812 1562
rect 31850 1527 31852 1536
rect 31760 1498 31812 1504
rect 31904 1527 31906 1536
rect 31852 1498 31904 1504
rect 31496 870 31616 898
rect 31496 762 31524 870
rect 31588 800 31616 870
rect 32232 800 32260 2246
rect 32876 800 32904 2382
rect 33520 800 33548 2858
rect 33872 2748 34180 2757
rect 33872 2746 33878 2748
rect 33934 2746 33958 2748
rect 34014 2746 34038 2748
rect 34094 2746 34118 2748
rect 34174 2746 34180 2748
rect 33934 2694 33936 2746
rect 34116 2694 34118 2746
rect 33872 2692 33878 2694
rect 33934 2692 33958 2694
rect 34014 2692 34038 2694
rect 34094 2692 34118 2694
rect 34174 2692 34180 2694
rect 33872 2683 34180 2692
rect 34888 2576 34940 2582
rect 34808 2536 34888 2564
rect 34808 2446 34836 2536
rect 34888 2518 34940 2524
rect 35360 2446 35388 15302
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 35452 14346 35480 14962
rect 35440 14340 35492 14346
rect 35440 14282 35492 14288
rect 35440 14068 35492 14074
rect 35440 14010 35492 14016
rect 35452 13938 35480 14010
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 35544 12889 35572 16390
rect 35716 16108 35768 16114
rect 35636 16068 35716 16096
rect 35636 15366 35664 16068
rect 35716 16050 35768 16056
rect 35912 15570 35940 16526
rect 36004 16454 36032 18226
rect 35992 16448 36044 16454
rect 35992 16390 36044 16396
rect 35900 15564 35952 15570
rect 35900 15506 35952 15512
rect 35624 15360 35676 15366
rect 36188 15314 36216 22578
rect 36268 18216 36320 18222
rect 36268 18158 36320 18164
rect 36280 17814 36308 18158
rect 36268 17808 36320 17814
rect 36268 17750 36320 17756
rect 35624 15302 35676 15308
rect 35636 14482 35664 15302
rect 36004 15286 36216 15314
rect 36280 15314 36308 17750
rect 36372 16658 36400 22714
rect 36452 18352 36504 18358
rect 36450 18320 36452 18329
rect 36504 18320 36506 18329
rect 36450 18255 36506 18264
rect 36452 17060 36504 17066
rect 36452 17002 36504 17008
rect 36464 16726 36492 17002
rect 36452 16720 36504 16726
rect 36452 16662 36504 16668
rect 36360 16652 36412 16658
rect 36360 16594 36412 16600
rect 36556 16250 36584 27610
rect 36832 27470 36860 29294
rect 37370 29294 37504 29322
rect 37370 29200 37426 29294
rect 37476 27606 37504 29294
rect 38014 29294 38148 29322
rect 38014 29200 38070 29294
rect 38120 27606 38148 29294
rect 38658 29294 38792 29322
rect 38658 29200 38714 29294
rect 38764 27606 38792 29294
rect 39302 29200 39358 30000
rect 40590 29322 40646 30000
rect 40590 29294 40724 29322
rect 40590 29200 40646 29294
rect 39316 27606 39344 29200
rect 40696 27606 40724 29294
rect 41234 29200 41290 30000
rect 41878 29322 41934 30000
rect 42522 29322 42578 30000
rect 43166 29322 43222 30000
rect 41878 29294 42012 29322
rect 41878 29200 41934 29294
rect 37280 27600 37332 27606
rect 37280 27542 37332 27548
rect 37464 27600 37516 27606
rect 37464 27542 37516 27548
rect 37556 27600 37608 27606
rect 37556 27542 37608 27548
rect 38108 27600 38160 27606
rect 38108 27542 38160 27548
rect 38752 27600 38804 27606
rect 38752 27542 38804 27548
rect 39304 27600 39356 27606
rect 39304 27542 39356 27548
rect 40684 27600 40736 27606
rect 40684 27542 40736 27548
rect 37292 27470 37320 27542
rect 36820 27464 36872 27470
rect 36820 27406 36872 27412
rect 37280 27464 37332 27470
rect 37280 27406 37332 27412
rect 37568 27130 37596 27542
rect 37832 27464 37884 27470
rect 37832 27406 37884 27412
rect 37924 27464 37976 27470
rect 37924 27406 37976 27412
rect 39120 27464 39172 27470
rect 39120 27406 39172 27412
rect 39856 27464 39908 27470
rect 39856 27406 39908 27412
rect 40684 27464 40736 27470
rect 40684 27406 40736 27412
rect 37556 27124 37608 27130
rect 37556 27066 37608 27072
rect 36820 23588 36872 23594
rect 36820 23530 36872 23536
rect 36832 20806 36860 23530
rect 37844 22094 37872 27406
rect 37936 27130 37964 27406
rect 37924 27124 37976 27130
rect 37924 27066 37976 27072
rect 38016 27124 38068 27130
rect 38016 27066 38068 27072
rect 38028 26994 38056 27066
rect 38568 27056 38620 27062
rect 38568 26998 38620 27004
rect 38016 26988 38068 26994
rect 38016 26930 38068 26936
rect 38108 26988 38160 26994
rect 38108 26930 38160 26936
rect 37844 22066 37964 22094
rect 36820 20800 36872 20806
rect 36820 20742 36872 20748
rect 37740 20800 37792 20806
rect 37740 20742 37792 20748
rect 36820 18284 36872 18290
rect 36820 18226 36872 18232
rect 36728 18216 36780 18222
rect 36728 18158 36780 18164
rect 36636 18080 36688 18086
rect 36636 18022 36688 18028
rect 36648 17678 36676 18022
rect 36636 17672 36688 17678
rect 36636 17614 36688 17620
rect 36740 16726 36768 18158
rect 36832 16998 36860 18226
rect 37556 17808 37608 17814
rect 37556 17750 37608 17756
rect 37568 17202 37596 17750
rect 37646 17232 37702 17241
rect 37556 17196 37608 17202
rect 37646 17167 37648 17176
rect 37556 17138 37608 17144
rect 37700 17167 37702 17176
rect 37648 17138 37700 17144
rect 36820 16992 36872 16998
rect 36820 16934 36872 16940
rect 36728 16720 36780 16726
rect 36728 16662 36780 16668
rect 36832 16658 36860 16934
rect 36820 16652 36872 16658
rect 36820 16594 36872 16600
rect 37556 16448 37608 16454
rect 37556 16390 37608 16396
rect 36544 16244 36596 16250
rect 36544 16186 36596 16192
rect 37568 16114 37596 16390
rect 37752 16114 37780 20742
rect 37832 17740 37884 17746
rect 37832 17682 37884 17688
rect 37844 17270 37872 17682
rect 37832 17264 37884 17270
rect 37832 17206 37884 17212
rect 37844 16250 37872 17206
rect 37832 16244 37884 16250
rect 37832 16186 37884 16192
rect 37556 16108 37608 16114
rect 37384 16068 37556 16096
rect 36360 15904 36412 15910
rect 36360 15846 36412 15852
rect 36372 15434 36400 15846
rect 37384 15570 37412 16068
rect 37556 16050 37608 16056
rect 37740 16108 37792 16114
rect 37740 16050 37792 16056
rect 37464 15904 37516 15910
rect 37464 15846 37516 15852
rect 37372 15564 37424 15570
rect 37372 15506 37424 15512
rect 37280 15496 37332 15502
rect 37280 15438 37332 15444
rect 36360 15428 36412 15434
rect 36360 15370 36412 15376
rect 36280 15286 36400 15314
rect 35900 14816 35952 14822
rect 35900 14758 35952 14764
rect 35624 14476 35676 14482
rect 35624 14418 35676 14424
rect 35808 14340 35860 14346
rect 35808 14282 35860 14288
rect 35820 14113 35848 14282
rect 35806 14104 35862 14113
rect 35806 14039 35862 14048
rect 35912 13938 35940 14758
rect 35900 13932 35952 13938
rect 35900 13874 35952 13880
rect 35808 13796 35860 13802
rect 35808 13738 35860 13744
rect 35714 13560 35770 13569
rect 35714 13495 35770 13504
rect 35728 13462 35756 13495
rect 35716 13456 35768 13462
rect 35716 13398 35768 13404
rect 35820 12918 35848 13738
rect 35900 13184 35952 13190
rect 35900 13126 35952 13132
rect 35808 12912 35860 12918
rect 35530 12880 35586 12889
rect 35440 12844 35492 12850
rect 35808 12854 35860 12860
rect 35530 12815 35586 12824
rect 35716 12844 35768 12850
rect 35440 12786 35492 12792
rect 35716 12786 35768 12792
rect 35452 12209 35480 12786
rect 35532 12300 35584 12306
rect 35532 12242 35584 12248
rect 35624 12300 35676 12306
rect 35624 12242 35676 12248
rect 35438 12200 35494 12209
rect 35438 12135 35494 12144
rect 35438 11792 35494 11801
rect 35438 11727 35494 11736
rect 35452 11626 35480 11727
rect 35440 11620 35492 11626
rect 35440 11562 35492 11568
rect 35544 3602 35572 12242
rect 35636 10962 35664 12242
rect 35728 11354 35756 12786
rect 35808 12436 35860 12442
rect 35808 12378 35860 12384
rect 35820 11937 35848 12378
rect 35912 12288 35940 13126
rect 36004 12442 36032 15286
rect 36174 15192 36230 15201
rect 36174 15127 36230 15136
rect 36188 15026 36216 15127
rect 36176 15020 36228 15026
rect 36176 14962 36228 14968
rect 36268 14952 36320 14958
rect 36266 14920 36268 14929
rect 36320 14920 36322 14929
rect 36266 14855 36322 14864
rect 36176 14340 36228 14346
rect 36176 14282 36228 14288
rect 36188 14074 36216 14282
rect 36176 14068 36228 14074
rect 36176 14010 36228 14016
rect 35992 12436 36044 12442
rect 35992 12378 36044 12384
rect 36176 12436 36228 12442
rect 36176 12378 36228 12384
rect 36084 12300 36136 12306
rect 35912 12260 36084 12288
rect 36084 12242 36136 12248
rect 35900 12096 35952 12102
rect 35900 12038 35952 12044
rect 35806 11928 35862 11937
rect 35806 11863 35862 11872
rect 35808 11756 35860 11762
rect 35912 11744 35940 12038
rect 35860 11716 35940 11744
rect 35808 11698 35860 11704
rect 35806 11656 35862 11665
rect 35806 11591 35862 11600
rect 35820 11354 35848 11591
rect 35992 11552 36044 11558
rect 35992 11494 36044 11500
rect 35716 11348 35768 11354
rect 35716 11290 35768 11296
rect 35808 11348 35860 11354
rect 35808 11290 35860 11296
rect 36004 11150 36032 11494
rect 36096 11150 36124 12242
rect 36188 12102 36216 12378
rect 36176 12096 36228 12102
rect 36268 12096 36320 12102
rect 36176 12038 36228 12044
rect 36266 12064 36268 12073
rect 36320 12064 36322 12073
rect 36266 11999 36322 12008
rect 36268 11688 36320 11694
rect 36266 11656 36268 11665
rect 36320 11656 36322 11665
rect 36266 11591 36322 11600
rect 36176 11552 36228 11558
rect 36176 11494 36228 11500
rect 35716 11144 35768 11150
rect 35992 11144 36044 11150
rect 35768 11092 35940 11098
rect 35716 11086 35940 11092
rect 35992 11086 36044 11092
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 35728 11070 35940 11086
rect 35912 10962 35940 11070
rect 36188 10962 36216 11494
rect 35636 10934 35756 10962
rect 35912 10934 36216 10962
rect 35728 9586 35756 10934
rect 36268 10668 36320 10674
rect 36268 10610 36320 10616
rect 35992 10056 36044 10062
rect 35992 9998 36044 10004
rect 35808 9920 35860 9926
rect 35808 9862 35860 9868
rect 35820 9654 35848 9862
rect 35808 9648 35860 9654
rect 35808 9590 35860 9596
rect 35716 9580 35768 9586
rect 35716 9522 35768 9528
rect 36004 9178 36032 9998
rect 36280 9722 36308 10610
rect 36268 9716 36320 9722
rect 36268 9658 36320 9664
rect 35992 9172 36044 9178
rect 35992 9114 36044 9120
rect 36280 8974 36308 9658
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 35532 3596 35584 3602
rect 35532 3538 35584 3544
rect 35716 2848 35768 2854
rect 35716 2790 35768 2796
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 34060 2304 34112 2310
rect 34060 2246 34112 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 34072 2145 34100 2246
rect 34058 2136 34114 2145
rect 34058 2071 34114 2080
rect 34164 800 34192 2246
rect 35452 800 35480 2382
rect 35728 1737 35756 2790
rect 36372 2514 36400 15286
rect 36452 15020 36504 15026
rect 36452 14962 36504 14968
rect 37096 15020 37148 15026
rect 37096 14962 37148 14968
rect 36464 13705 36492 14962
rect 37108 14618 37136 14962
rect 37292 14958 37320 15438
rect 37280 14952 37332 14958
rect 37200 14912 37280 14940
rect 37096 14612 37148 14618
rect 37096 14554 37148 14560
rect 36634 14376 36690 14385
rect 36634 14311 36690 14320
rect 36450 13696 36506 13705
rect 36450 13631 36506 13640
rect 36452 12980 36504 12986
rect 36452 12922 36504 12928
rect 36464 12356 36492 12922
rect 36544 12844 36596 12850
rect 36648 12832 36676 14311
rect 37004 14272 37056 14278
rect 37002 14240 37004 14249
rect 37096 14272 37148 14278
rect 37056 14240 37058 14249
rect 37096 14214 37148 14220
rect 37002 14175 37058 14184
rect 37002 13832 37058 13841
rect 37002 13767 37058 13776
rect 36820 13388 36872 13394
rect 36820 13330 36872 13336
rect 36728 13184 36780 13190
rect 36728 13126 36780 13132
rect 36596 12804 36676 12832
rect 36544 12786 36596 12792
rect 36648 12646 36676 12804
rect 36544 12640 36596 12646
rect 36544 12582 36596 12588
rect 36636 12640 36688 12646
rect 36636 12582 36688 12588
rect 36556 12434 36584 12582
rect 36556 12406 36676 12434
rect 36544 12368 36596 12374
rect 36464 12328 36544 12356
rect 36544 12310 36596 12316
rect 36556 12238 36584 12310
rect 36544 12232 36596 12238
rect 36544 12174 36596 12180
rect 36452 11756 36504 11762
rect 36452 11698 36504 11704
rect 36464 11150 36492 11698
rect 36556 11218 36584 12174
rect 36648 12050 36676 12406
rect 36740 12238 36768 13126
rect 36832 12238 36860 13330
rect 36912 13184 36964 13190
rect 36910 13152 36912 13161
rect 36964 13152 36966 13161
rect 36910 13087 36966 13096
rect 37016 12918 37044 13767
rect 37004 12912 37056 12918
rect 37004 12854 37056 12860
rect 37108 12238 37136 14214
rect 37200 13530 37228 14912
rect 37384 14929 37412 15506
rect 37280 14894 37332 14900
rect 37370 14920 37426 14929
rect 37370 14855 37426 14864
rect 37370 14240 37426 14249
rect 37370 14175 37426 14184
rect 37278 14104 37334 14113
rect 37278 14039 37334 14048
rect 37188 13524 37240 13530
rect 37188 13466 37240 13472
rect 37292 13161 37320 14039
rect 37278 13152 37334 13161
rect 37278 13087 37334 13096
rect 36728 12232 36780 12238
rect 36728 12174 36780 12180
rect 36820 12232 36872 12238
rect 36820 12174 36872 12180
rect 37096 12232 37148 12238
rect 37096 12174 37148 12180
rect 37186 12200 37242 12209
rect 37186 12135 37242 12144
rect 36648 12022 36952 12050
rect 36726 11792 36782 11801
rect 36726 11727 36728 11736
rect 36780 11727 36782 11736
rect 36728 11698 36780 11704
rect 36636 11688 36688 11694
rect 36688 11636 36768 11642
rect 36636 11630 36768 11636
rect 36648 11626 36768 11630
rect 36648 11620 36780 11626
rect 36648 11614 36728 11620
rect 36728 11562 36780 11568
rect 36924 11558 36952 12022
rect 37004 11688 37056 11694
rect 37004 11630 37056 11636
rect 36912 11552 36964 11558
rect 36912 11494 36964 11500
rect 36544 11212 36596 11218
rect 36544 11154 36596 11160
rect 36452 11144 36504 11150
rect 36452 11086 36504 11092
rect 36464 10674 36492 11086
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36728 8832 36780 8838
rect 36728 8774 36780 8780
rect 36740 7274 36768 8774
rect 36728 7268 36780 7274
rect 36728 7210 36780 7216
rect 36544 4004 36596 4010
rect 36544 3946 36596 3952
rect 36556 3534 36584 3946
rect 36544 3528 36596 3534
rect 36544 3470 36596 3476
rect 36924 2774 36952 11494
rect 37016 10810 37044 11630
rect 37200 11626 37228 12135
rect 37292 11830 37320 13087
rect 37384 11898 37412 14175
rect 37372 11892 37424 11898
rect 37372 11834 37424 11840
rect 37280 11824 37332 11830
rect 37280 11766 37332 11772
rect 37188 11620 37240 11626
rect 37372 11620 37424 11626
rect 37188 11562 37240 11568
rect 37292 11580 37372 11608
rect 37094 11248 37150 11257
rect 37094 11183 37150 11192
rect 37108 11150 37136 11183
rect 37096 11144 37148 11150
rect 37096 11086 37148 11092
rect 37094 10840 37150 10849
rect 37004 10804 37056 10810
rect 37094 10775 37150 10784
rect 37004 10746 37056 10752
rect 37108 10606 37136 10775
rect 37096 10600 37148 10606
rect 37096 10542 37148 10548
rect 37292 3466 37320 11580
rect 37372 11562 37424 11568
rect 37372 10668 37424 10674
rect 37372 10610 37424 10616
rect 37384 9178 37412 10610
rect 37372 9172 37424 9178
rect 37372 9114 37424 9120
rect 37280 3460 37332 3466
rect 37280 3402 37332 3408
rect 37476 2854 37504 15846
rect 37648 15496 37700 15502
rect 37648 15438 37700 15444
rect 37556 15360 37608 15366
rect 37556 15302 37608 15308
rect 37568 14414 37596 15302
rect 37556 14408 37608 14414
rect 37556 14350 37608 14356
rect 37556 13932 37608 13938
rect 37556 13874 37608 13880
rect 37568 13841 37596 13874
rect 37554 13832 37610 13841
rect 37554 13767 37556 13776
rect 37608 13767 37610 13776
rect 37556 13738 37608 13744
rect 37568 13707 37596 13738
rect 37660 12850 37688 15438
rect 37752 13938 37780 16050
rect 37832 16040 37884 16046
rect 37832 15982 37884 15988
rect 37844 15434 37872 15982
rect 37832 15428 37884 15434
rect 37832 15370 37884 15376
rect 37832 15020 37884 15026
rect 37832 14962 37884 14968
rect 37844 14618 37872 14962
rect 37936 14929 37964 22066
rect 38120 19378 38148 26930
rect 38292 26920 38344 26926
rect 38198 26888 38254 26897
rect 38292 26862 38344 26868
rect 38198 26823 38254 26832
rect 38212 26382 38240 26823
rect 38304 26518 38332 26862
rect 38292 26512 38344 26518
rect 38292 26454 38344 26460
rect 38200 26376 38252 26382
rect 38200 26318 38252 26324
rect 38580 22642 38608 26998
rect 38568 22636 38620 22642
rect 38568 22578 38620 22584
rect 38384 19984 38436 19990
rect 38384 19926 38436 19932
rect 38108 19372 38160 19378
rect 38108 19314 38160 19320
rect 38200 17536 38252 17542
rect 38200 17478 38252 17484
rect 38212 17202 38240 17478
rect 38200 17196 38252 17202
rect 38200 17138 38252 17144
rect 38212 16590 38240 17138
rect 38200 16584 38252 16590
rect 38200 16526 38252 16532
rect 38396 15570 38424 19926
rect 39132 18698 39160 27406
rect 39396 26444 39448 26450
rect 39396 26386 39448 26392
rect 39120 18692 39172 18698
rect 39120 18634 39172 18640
rect 38750 16688 38806 16697
rect 38750 16623 38752 16632
rect 38804 16623 38806 16632
rect 38752 16594 38804 16600
rect 38660 16448 38712 16454
rect 38660 16390 38712 16396
rect 38672 16250 38700 16390
rect 38660 16244 38712 16250
rect 38660 16186 38712 16192
rect 38384 15564 38436 15570
rect 38384 15506 38436 15512
rect 38568 15428 38620 15434
rect 38568 15370 38620 15376
rect 37922 14920 37978 14929
rect 37922 14855 37978 14864
rect 38580 14822 38608 15370
rect 39302 15192 39358 15201
rect 39302 15127 39358 15136
rect 38568 14816 38620 14822
rect 38568 14758 38620 14764
rect 37832 14612 37884 14618
rect 37832 14554 37884 14560
rect 38580 14482 38608 14758
rect 38568 14476 38620 14482
rect 38568 14418 38620 14424
rect 37924 14408 37976 14414
rect 38292 14408 38344 14414
rect 37924 14350 37976 14356
rect 38290 14376 38292 14385
rect 38476 14408 38528 14414
rect 38344 14376 38346 14385
rect 37936 14074 37964 14350
rect 38476 14350 38528 14356
rect 38290 14311 38346 14320
rect 37924 14068 37976 14074
rect 37924 14010 37976 14016
rect 38212 14062 38424 14090
rect 38212 13954 38240 14062
rect 37740 13932 37792 13938
rect 37740 13874 37792 13880
rect 37844 13926 38240 13954
rect 38396 13938 38424 14062
rect 38292 13932 38344 13938
rect 37648 12844 37700 12850
rect 37648 12786 37700 12792
rect 37556 12300 37608 12306
rect 37556 12242 37608 12248
rect 37568 11626 37596 12242
rect 37556 11620 37608 11626
rect 37556 11562 37608 11568
rect 37556 11076 37608 11082
rect 37556 11018 37608 11024
rect 37568 10810 37596 11018
rect 37556 10804 37608 10810
rect 37556 10746 37608 10752
rect 37660 10674 37688 12786
rect 37738 11928 37794 11937
rect 37738 11863 37794 11872
rect 37752 11218 37780 11863
rect 37740 11212 37792 11218
rect 37740 11154 37792 11160
rect 37740 11008 37792 11014
rect 37738 10976 37740 10985
rect 37792 10976 37794 10985
rect 37738 10911 37794 10920
rect 37648 10668 37700 10674
rect 37648 10610 37700 10616
rect 37556 10600 37608 10606
rect 37556 10542 37608 10548
rect 37568 10062 37596 10542
rect 37660 10418 37688 10610
rect 37660 10390 37780 10418
rect 37556 10056 37608 10062
rect 37556 9998 37608 10004
rect 37568 9586 37596 9998
rect 37648 9716 37700 9722
rect 37648 9658 37700 9664
rect 37556 9580 37608 9586
rect 37556 9522 37608 9528
rect 37568 8974 37596 9522
rect 37660 8974 37688 9658
rect 37752 9110 37780 10390
rect 37740 9104 37792 9110
rect 37740 9046 37792 9052
rect 37556 8968 37608 8974
rect 37556 8910 37608 8916
rect 37648 8968 37700 8974
rect 37648 8910 37700 8916
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 37844 2774 37872 13926
rect 38292 13874 38344 13880
rect 38384 13932 38436 13938
rect 38384 13874 38436 13880
rect 37924 13728 37976 13734
rect 37924 13670 37976 13676
rect 38108 13728 38160 13734
rect 38108 13670 38160 13676
rect 37936 12782 37964 13670
rect 37924 12776 37976 12782
rect 37924 12718 37976 12724
rect 38016 12776 38068 12782
rect 38016 12718 38068 12724
rect 37936 4758 37964 12718
rect 38028 12374 38056 12718
rect 38016 12368 38068 12374
rect 38016 12310 38068 12316
rect 38120 12238 38148 13670
rect 38304 12986 38332 13874
rect 38488 12986 38516 14350
rect 39316 14074 39344 15127
rect 39408 15042 39436 26386
rect 39488 18352 39540 18358
rect 39488 18294 39540 18300
rect 39500 17270 39528 18294
rect 39488 17264 39540 17270
rect 39488 17206 39540 17212
rect 39580 17060 39632 17066
rect 39580 17002 39632 17008
rect 39592 16833 39620 17002
rect 39578 16824 39634 16833
rect 39578 16759 39634 16768
rect 39408 15014 39528 15042
rect 39396 14952 39448 14958
rect 39396 14894 39448 14900
rect 39408 14550 39436 14894
rect 39396 14544 39448 14550
rect 39396 14486 39448 14492
rect 39396 14408 39448 14414
rect 39396 14350 39448 14356
rect 39408 14074 39436 14350
rect 38752 14068 38804 14074
rect 38752 14010 38804 14016
rect 39304 14068 39356 14074
rect 39304 14010 39356 14016
rect 39396 14068 39448 14074
rect 39396 14010 39448 14016
rect 38764 13734 38792 14010
rect 38844 14000 38896 14006
rect 38844 13942 38896 13948
rect 38752 13728 38804 13734
rect 38752 13670 38804 13676
rect 38750 13560 38806 13569
rect 38856 13530 38884 13942
rect 39396 13864 39448 13870
rect 39500 13852 39528 15014
rect 39764 14476 39816 14482
rect 39764 14418 39816 14424
rect 39776 13870 39804 14418
rect 39448 13824 39528 13852
rect 39764 13864 39816 13870
rect 39396 13806 39448 13812
rect 39764 13806 39816 13812
rect 39408 13705 39436 13806
rect 39394 13696 39450 13705
rect 39394 13631 39450 13640
rect 39394 13560 39450 13569
rect 38750 13495 38806 13504
rect 38844 13524 38896 13530
rect 38660 13456 38712 13462
rect 38660 13398 38712 13404
rect 38292 12980 38344 12986
rect 38292 12922 38344 12928
rect 38476 12980 38528 12986
rect 38476 12922 38528 12928
rect 38384 12912 38436 12918
rect 38384 12854 38436 12860
rect 38016 12232 38068 12238
rect 38016 12174 38068 12180
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 38028 9586 38056 12174
rect 38396 11830 38424 12854
rect 38384 11824 38436 11830
rect 38384 11766 38436 11772
rect 38488 11694 38516 12922
rect 38566 12336 38622 12345
rect 38566 12271 38622 12280
rect 38580 12238 38608 12271
rect 38568 12232 38620 12238
rect 38568 12174 38620 12180
rect 38200 11688 38252 11694
rect 38200 11630 38252 11636
rect 38476 11688 38528 11694
rect 38476 11630 38528 11636
rect 38212 11218 38240 11630
rect 38292 11620 38344 11626
rect 38292 11562 38344 11568
rect 38304 11393 38332 11562
rect 38290 11384 38346 11393
rect 38290 11319 38346 11328
rect 38568 11348 38620 11354
rect 38568 11290 38620 11296
rect 38200 11212 38252 11218
rect 38200 11154 38252 11160
rect 38476 11212 38528 11218
rect 38476 11154 38528 11160
rect 38108 11144 38160 11150
rect 38106 11112 38108 11121
rect 38160 11112 38162 11121
rect 38106 11047 38162 11056
rect 38212 10742 38240 11154
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38200 10736 38252 10742
rect 38200 10678 38252 10684
rect 38108 10260 38160 10266
rect 38108 10202 38160 10208
rect 38120 9926 38148 10202
rect 38108 9920 38160 9926
rect 38108 9862 38160 9868
rect 38200 9920 38252 9926
rect 38200 9862 38252 9868
rect 38016 9580 38068 9586
rect 38016 9522 38068 9528
rect 38212 8498 38240 9862
rect 38304 9654 38332 11086
rect 38488 10810 38516 11154
rect 38580 11082 38608 11290
rect 38568 11076 38620 11082
rect 38568 11018 38620 11024
rect 38476 10804 38528 10810
rect 38476 10746 38528 10752
rect 38568 10668 38620 10674
rect 38568 10610 38620 10616
rect 38384 10600 38436 10606
rect 38580 10577 38608 10610
rect 38384 10542 38436 10548
rect 38566 10568 38622 10577
rect 38396 9722 38424 10542
rect 38566 10503 38622 10512
rect 38672 10112 38700 13398
rect 38764 13394 38792 13495
rect 39394 13495 39450 13504
rect 38844 13466 38896 13472
rect 38752 13388 38804 13394
rect 38752 13330 38804 13336
rect 39408 13326 39436 13495
rect 39304 13320 39356 13326
rect 39304 13262 39356 13268
rect 39396 13320 39448 13326
rect 39396 13262 39448 13268
rect 38936 13252 38988 13258
rect 38936 13194 38988 13200
rect 38948 12918 38976 13194
rect 38936 12912 38988 12918
rect 38936 12854 38988 12860
rect 39120 12912 39172 12918
rect 39120 12854 39172 12860
rect 38842 12336 38898 12345
rect 38842 12271 38898 12280
rect 38752 11620 38804 11626
rect 38752 11562 38804 11568
rect 38764 11354 38792 11562
rect 38856 11354 38884 12271
rect 39026 12064 39082 12073
rect 39026 11999 39082 12008
rect 38936 11688 38988 11694
rect 38936 11630 38988 11636
rect 38752 11348 38804 11354
rect 38752 11290 38804 11296
rect 38844 11348 38896 11354
rect 38844 11290 38896 11296
rect 38948 11257 38976 11630
rect 39040 11558 39068 11999
rect 39028 11552 39080 11558
rect 39028 11494 39080 11500
rect 39040 11286 39068 11494
rect 39028 11280 39080 11286
rect 38934 11248 38990 11257
rect 38844 11212 38896 11218
rect 39028 11222 39080 11228
rect 38934 11183 38990 11192
rect 38844 11154 38896 11160
rect 38856 10849 38884 11154
rect 38948 11150 38976 11183
rect 38936 11144 38988 11150
rect 38936 11086 38988 11092
rect 39028 11144 39080 11150
rect 39028 11086 39080 11092
rect 38842 10840 38898 10849
rect 38842 10775 38898 10784
rect 38752 10464 38804 10470
rect 38752 10406 38804 10412
rect 38936 10464 38988 10470
rect 38936 10406 38988 10412
rect 38580 10084 38700 10112
rect 38384 9716 38436 9722
rect 38384 9658 38436 9664
rect 38292 9648 38344 9654
rect 38292 9590 38344 9596
rect 38580 9382 38608 10084
rect 38658 10024 38714 10033
rect 38658 9959 38660 9968
rect 38712 9959 38714 9968
rect 38660 9930 38712 9936
rect 38568 9376 38620 9382
rect 38568 9318 38620 9324
rect 38200 8492 38252 8498
rect 38200 8434 38252 8440
rect 38672 7478 38700 9930
rect 38764 8974 38792 10406
rect 38844 10260 38896 10266
rect 38844 10202 38896 10208
rect 38856 9926 38884 10202
rect 38844 9920 38896 9926
rect 38844 9862 38896 9868
rect 38844 9580 38896 9586
rect 38844 9522 38896 9528
rect 38856 9178 38884 9522
rect 38844 9172 38896 9178
rect 38844 9114 38896 9120
rect 38752 8968 38804 8974
rect 38752 8910 38804 8916
rect 38660 7472 38712 7478
rect 38660 7414 38712 7420
rect 37924 4752 37976 4758
rect 37924 4694 37976 4700
rect 38844 4480 38896 4486
rect 38844 4422 38896 4428
rect 38108 4004 38160 4010
rect 38108 3946 38160 3952
rect 38120 3602 38148 3946
rect 38108 3596 38160 3602
rect 38108 3538 38160 3544
rect 36832 2746 36952 2774
rect 37660 2746 37872 2774
rect 36360 2508 36412 2514
rect 36360 2450 36412 2456
rect 36832 2446 36860 2746
rect 37660 2446 37688 2746
rect 38856 2632 38884 4422
rect 38948 3058 38976 10406
rect 39040 9874 39068 11086
rect 39132 10742 39160 12854
rect 39316 12424 39344 13262
rect 39396 12436 39448 12442
rect 39316 12396 39396 12424
rect 39868 12434 39896 27406
rect 40696 27130 40724 27406
rect 41248 27334 41276 29200
rect 41984 27470 42012 29294
rect 42522 29294 42656 29322
rect 42522 29200 42578 29294
rect 42628 27606 42656 29294
rect 43166 29294 43300 29322
rect 43166 29200 43222 29294
rect 43272 27606 43300 29294
rect 43810 29200 43866 30000
rect 44454 29322 44510 30000
rect 45098 29322 45154 30000
rect 45742 29322 45798 30000
rect 46386 29322 46442 30000
rect 44454 29294 44588 29322
rect 44454 29200 44510 29294
rect 43824 27606 43852 29200
rect 42616 27600 42668 27606
rect 42616 27542 42668 27548
rect 43260 27600 43312 27606
rect 43260 27542 43312 27548
rect 43812 27600 43864 27606
rect 43812 27542 43864 27548
rect 42524 27532 42576 27538
rect 42524 27474 42576 27480
rect 41604 27464 41656 27470
rect 41604 27406 41656 27412
rect 41972 27464 42024 27470
rect 41972 27406 42024 27412
rect 41052 27328 41104 27334
rect 41052 27270 41104 27276
rect 41236 27328 41288 27334
rect 41236 27270 41288 27276
rect 40684 27124 40736 27130
rect 40684 27066 40736 27072
rect 40682 27024 40738 27033
rect 41064 26994 41092 27270
rect 40682 26959 40738 26968
rect 40776 26988 40828 26994
rect 40696 26518 40724 26959
rect 40776 26930 40828 26936
rect 40960 26988 41012 26994
rect 40960 26930 41012 26936
rect 41052 26988 41104 26994
rect 41052 26930 41104 26936
rect 41420 26988 41472 26994
rect 41420 26930 41472 26936
rect 40684 26512 40736 26518
rect 40684 26454 40736 26460
rect 40684 26376 40736 26382
rect 40682 26344 40684 26353
rect 40736 26344 40738 26353
rect 40682 26279 40738 26288
rect 40788 22094 40816 26930
rect 40972 26518 41000 26930
rect 41432 26790 41460 26930
rect 41052 26784 41104 26790
rect 41052 26726 41104 26732
rect 41420 26784 41472 26790
rect 41420 26726 41472 26732
rect 41064 26518 41092 26726
rect 40960 26512 41012 26518
rect 40960 26454 41012 26460
rect 41052 26512 41104 26518
rect 41052 26454 41104 26460
rect 40868 26376 40920 26382
rect 40868 26318 40920 26324
rect 40880 26246 40908 26318
rect 40868 26240 40920 26246
rect 40868 26182 40920 26188
rect 40788 22066 40908 22094
rect 40682 17912 40738 17921
rect 40682 17847 40738 17856
rect 40500 17808 40552 17814
rect 40500 17750 40552 17756
rect 40224 17536 40276 17542
rect 40224 17478 40276 17484
rect 40132 17196 40184 17202
rect 40132 17138 40184 17144
rect 40144 16726 40172 17138
rect 40132 16720 40184 16726
rect 40132 16662 40184 16668
rect 40236 16590 40264 17478
rect 40512 17241 40540 17750
rect 40696 17746 40724 17847
rect 40684 17740 40736 17746
rect 40684 17682 40736 17688
rect 40498 17232 40554 17241
rect 40498 17167 40554 17176
rect 40316 16992 40368 16998
rect 40316 16934 40368 16940
rect 40328 16726 40356 16934
rect 40316 16720 40368 16726
rect 40316 16662 40368 16668
rect 40224 16584 40276 16590
rect 40224 16526 40276 16532
rect 40684 15972 40736 15978
rect 40684 15914 40736 15920
rect 39948 15020 40000 15026
rect 39948 14962 40000 14968
rect 39960 14521 39988 14962
rect 39946 14512 40002 14521
rect 39946 14447 40002 14456
rect 40592 14408 40644 14414
rect 40592 14350 40644 14356
rect 39948 14340 40000 14346
rect 40224 14340 40276 14346
rect 40000 14300 40224 14328
rect 39948 14282 40000 14288
rect 40224 14282 40276 14288
rect 39948 13864 40000 13870
rect 40130 13832 40186 13841
rect 40000 13812 40080 13818
rect 39948 13806 40080 13812
rect 39960 13790 40080 13806
rect 39948 13456 40000 13462
rect 39948 13398 40000 13404
rect 39960 12646 39988 13398
rect 40052 12918 40080 13790
rect 40130 13767 40186 13776
rect 40314 13832 40370 13841
rect 40314 13767 40316 13776
rect 40144 13326 40172 13767
rect 40368 13767 40370 13776
rect 40316 13738 40368 13744
rect 40408 13388 40460 13394
rect 40408 13330 40460 13336
rect 40132 13320 40184 13326
rect 40132 13262 40184 13268
rect 40040 12912 40092 12918
rect 40040 12854 40092 12860
rect 39948 12640 40000 12646
rect 39948 12582 40000 12588
rect 39396 12378 39448 12384
rect 39776 12406 39896 12434
rect 39672 12164 39724 12170
rect 39672 12106 39724 12112
rect 39394 11792 39450 11801
rect 39684 11762 39712 12106
rect 39394 11727 39450 11736
rect 39672 11756 39724 11762
rect 39408 11694 39436 11727
rect 39672 11698 39724 11704
rect 39396 11688 39448 11694
rect 39396 11630 39448 11636
rect 39212 11144 39264 11150
rect 39212 11086 39264 11092
rect 39120 10736 39172 10742
rect 39120 10678 39172 10684
rect 39132 10033 39160 10678
rect 39224 10266 39252 11086
rect 39408 10674 39436 11630
rect 39486 10840 39542 10849
rect 39486 10775 39542 10784
rect 39500 10674 39528 10775
rect 39396 10668 39448 10674
rect 39396 10610 39448 10616
rect 39488 10668 39540 10674
rect 39488 10610 39540 10616
rect 39304 10600 39356 10606
rect 39304 10542 39356 10548
rect 39212 10260 39264 10266
rect 39212 10202 39264 10208
rect 39316 10130 39344 10542
rect 39776 10470 39804 12406
rect 40040 12232 40092 12238
rect 40038 12200 40040 12209
rect 40092 12200 40094 12209
rect 40144 12170 40172 13262
rect 40420 12850 40448 13330
rect 40604 13161 40632 14350
rect 40590 13152 40646 13161
rect 40590 13087 40646 13096
rect 40408 12844 40460 12850
rect 40408 12786 40460 12792
rect 40224 12640 40276 12646
rect 40224 12582 40276 12588
rect 40236 12238 40264 12582
rect 40224 12232 40276 12238
rect 40224 12174 40276 12180
rect 40038 12135 40094 12144
rect 40132 12164 40184 12170
rect 40132 12106 40184 12112
rect 40420 11762 40448 12786
rect 40500 12232 40552 12238
rect 40500 12174 40552 12180
rect 40224 11756 40276 11762
rect 40224 11698 40276 11704
rect 40408 11756 40460 11762
rect 40408 11698 40460 11704
rect 39856 11688 39908 11694
rect 39856 11630 39908 11636
rect 39868 11354 39896 11630
rect 39856 11348 39908 11354
rect 39856 11290 39908 11296
rect 40132 11348 40184 11354
rect 40132 11290 40184 11296
rect 40040 11144 40092 11150
rect 40040 11086 40092 11092
rect 39764 10464 39816 10470
rect 39764 10406 39816 10412
rect 39304 10124 39356 10130
rect 39304 10066 39356 10072
rect 40052 10062 40080 11086
rect 40144 11014 40172 11290
rect 40236 11150 40264 11698
rect 40316 11552 40368 11558
rect 40316 11494 40368 11500
rect 40224 11144 40276 11150
rect 40224 11086 40276 11092
rect 40132 11008 40184 11014
rect 40132 10950 40184 10956
rect 40144 10062 40172 10950
rect 40236 10810 40264 11086
rect 40328 11014 40356 11494
rect 40316 11008 40368 11014
rect 40316 10950 40368 10956
rect 40224 10804 40276 10810
rect 40224 10746 40276 10752
rect 40040 10056 40092 10062
rect 39118 10024 39174 10033
rect 40040 9998 40092 10004
rect 40132 10056 40184 10062
rect 40132 9998 40184 10004
rect 39118 9959 39174 9968
rect 39304 9920 39356 9926
rect 39040 9868 39304 9874
rect 39040 9862 39356 9868
rect 39040 9846 39344 9862
rect 39028 8560 39080 8566
rect 39028 8502 39080 8508
rect 38936 3052 38988 3058
rect 38936 2994 38988 3000
rect 38847 2604 38884 2632
rect 38752 2576 38804 2582
rect 38847 2564 38875 2604
rect 38804 2536 38875 2564
rect 38936 2576 38988 2582
rect 38752 2518 38804 2524
rect 38936 2518 38988 2524
rect 36820 2440 36872 2446
rect 36820 2382 36872 2388
rect 37648 2440 37700 2446
rect 37648 2382 37700 2388
rect 38752 2440 38804 2446
rect 38948 2428 38976 2518
rect 38804 2400 38976 2428
rect 38752 2382 38804 2388
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 38752 2304 38804 2310
rect 39040 2292 39068 8502
rect 39120 6792 39172 6798
rect 39120 6734 39172 6740
rect 39132 3126 39160 6734
rect 39120 3120 39172 3126
rect 39120 3062 39172 3068
rect 39120 2372 39172 2378
rect 39120 2314 39172 2320
rect 38804 2264 39068 2292
rect 38752 2246 38804 2252
rect 35714 1728 35770 1737
rect 35714 1663 35770 1672
rect 36096 800 36124 2246
rect 36740 800 36768 2246
rect 37384 800 37412 2246
rect 38672 1873 38700 2246
rect 38658 1864 38714 1873
rect 38658 1799 38714 1808
rect 39132 1290 39160 2314
rect 39224 1290 39252 9846
rect 39304 9376 39356 9382
rect 39304 9318 39356 9324
rect 39316 8362 39344 9318
rect 40144 9042 40172 9998
rect 40236 9382 40264 10746
rect 40316 10668 40368 10674
rect 40316 10610 40368 10616
rect 40328 10266 40356 10610
rect 40316 10260 40368 10266
rect 40316 10202 40368 10208
rect 40316 9580 40368 9586
rect 40316 9522 40368 9528
rect 40408 9580 40460 9586
rect 40408 9522 40460 9528
rect 40224 9376 40276 9382
rect 40224 9318 40276 9324
rect 40132 9036 40184 9042
rect 40132 8978 40184 8984
rect 39304 8356 39356 8362
rect 39304 8298 39356 8304
rect 39948 6724 40000 6730
rect 39948 6666 40000 6672
rect 39304 3596 39356 3602
rect 39304 3538 39356 3544
rect 39316 3058 39344 3538
rect 39396 3392 39448 3398
rect 39396 3334 39448 3340
rect 39304 3052 39356 3058
rect 39304 2994 39356 3000
rect 39408 2990 39436 3334
rect 39396 2984 39448 2990
rect 39960 2961 39988 6666
rect 40236 3058 40264 9318
rect 40328 9042 40356 9522
rect 40316 9036 40368 9042
rect 40316 8978 40368 8984
rect 40328 7546 40356 8978
rect 40420 8634 40448 9522
rect 40408 8628 40460 8634
rect 40408 8570 40460 8576
rect 40512 8514 40540 12174
rect 40592 12096 40644 12102
rect 40592 12038 40644 12044
rect 40604 11694 40632 12038
rect 40592 11688 40644 11694
rect 40592 11630 40644 11636
rect 40420 8486 40540 8514
rect 40316 7540 40368 7546
rect 40316 7482 40368 7488
rect 40224 3052 40276 3058
rect 40224 2994 40276 3000
rect 39396 2926 39448 2932
rect 39946 2952 40002 2961
rect 39946 2887 40002 2896
rect 39764 2848 39816 2854
rect 39764 2790 39816 2796
rect 39948 2848 40000 2854
rect 39948 2790 40000 2796
rect 39776 2514 39804 2790
rect 39764 2508 39816 2514
rect 39764 2450 39816 2456
rect 39304 2440 39356 2446
rect 39304 2382 39356 2388
rect 38660 1284 38712 1290
rect 38660 1226 38712 1232
rect 39120 1284 39172 1290
rect 39120 1226 39172 1232
rect 39212 1284 39264 1290
rect 39212 1226 39264 1232
rect 38672 800 38700 1226
rect 39316 800 39344 2382
rect 39960 800 39988 2790
rect 40420 2774 40448 8486
rect 40696 2774 40724 15914
rect 40774 15192 40830 15201
rect 40774 15127 40830 15136
rect 40788 14822 40816 15127
rect 40776 14816 40828 14822
rect 40776 14758 40828 14764
rect 40776 14272 40828 14278
rect 40776 14214 40828 14220
rect 40788 13802 40816 14214
rect 40776 13796 40828 13802
rect 40776 13738 40828 13744
rect 40776 13388 40828 13394
rect 40776 13330 40828 13336
rect 40788 11694 40816 13330
rect 40776 11688 40828 11694
rect 40776 11630 40828 11636
rect 40776 11552 40828 11558
rect 40776 11494 40828 11500
rect 40788 10674 40816 11494
rect 40880 11150 40908 22066
rect 41236 18624 41288 18630
rect 41236 18566 41288 18572
rect 41248 17202 41276 18566
rect 41512 18352 41564 18358
rect 41512 18294 41564 18300
rect 41524 17882 41552 18294
rect 41512 17876 41564 17882
rect 41512 17818 41564 17824
rect 41510 17776 41566 17785
rect 41432 17746 41510 17762
rect 41420 17740 41510 17746
rect 41472 17734 41510 17740
rect 41510 17711 41566 17720
rect 41420 17682 41472 17688
rect 41328 17672 41380 17678
rect 41328 17614 41380 17620
rect 41512 17672 41564 17678
rect 41512 17614 41564 17620
rect 41340 17513 41368 17614
rect 41420 17604 41472 17610
rect 41420 17546 41472 17552
rect 41326 17504 41382 17513
rect 41326 17439 41382 17448
rect 41236 17196 41288 17202
rect 41236 17138 41288 17144
rect 41432 17066 41460 17546
rect 41524 17270 41552 17614
rect 41512 17264 41564 17270
rect 41512 17206 41564 17212
rect 41420 17060 41472 17066
rect 41420 17002 41472 17008
rect 41432 16114 41460 17002
rect 41512 16992 41564 16998
rect 41512 16934 41564 16940
rect 41524 16590 41552 16934
rect 41512 16584 41564 16590
rect 41512 16526 41564 16532
rect 41420 16108 41472 16114
rect 41420 16050 41472 16056
rect 41512 15360 41564 15366
rect 41512 15302 41564 15308
rect 41524 15162 41552 15302
rect 41512 15156 41564 15162
rect 41512 15098 41564 15104
rect 41616 14657 41644 27406
rect 42536 27130 42564 27474
rect 44560 27470 44588 29294
rect 45098 29294 45232 29322
rect 45098 29200 45154 29294
rect 45204 27606 45232 29294
rect 45742 29294 45876 29322
rect 45742 29200 45798 29294
rect 45848 27606 45876 29294
rect 46386 29294 46520 29322
rect 46386 29200 46442 29294
rect 46492 27606 46520 29294
rect 47030 29200 47086 30000
rect 48318 29322 48374 30000
rect 48962 29322 49018 30000
rect 48318 29294 48636 29322
rect 48318 29200 48374 29294
rect 45192 27600 45244 27606
rect 45192 27542 45244 27548
rect 45836 27600 45888 27606
rect 45836 27542 45888 27548
rect 46480 27600 46532 27606
rect 46480 27542 46532 27548
rect 48608 27470 48636 29294
rect 48962 29294 49096 29322
rect 48962 29200 49018 29294
rect 49068 27606 49096 29294
rect 49606 29200 49662 30000
rect 50250 29322 50306 30000
rect 50894 29322 50950 30000
rect 51538 29322 51594 30000
rect 52182 29322 52238 30000
rect 50250 29294 50568 29322
rect 50250 29200 50306 29294
rect 49056 27600 49108 27606
rect 49056 27542 49108 27548
rect 42708 27464 42760 27470
rect 42614 27432 42670 27441
rect 42708 27406 42760 27412
rect 42800 27464 42852 27470
rect 42800 27406 42852 27412
rect 43444 27464 43496 27470
rect 43444 27406 43496 27412
rect 43996 27464 44048 27470
rect 43996 27406 44048 27412
rect 44548 27464 44600 27470
rect 44548 27406 44600 27412
rect 45376 27464 45428 27470
rect 45376 27406 45428 27412
rect 45468 27464 45520 27470
rect 45468 27406 45520 27412
rect 46664 27464 46716 27470
rect 48596 27464 48648 27470
rect 46664 27406 46716 27412
rect 46754 27432 46810 27441
rect 42614 27367 42616 27376
rect 42668 27367 42670 27376
rect 42616 27338 42668 27344
rect 42524 27124 42576 27130
rect 42524 27066 42576 27072
rect 42720 27033 42748 27406
rect 41786 27024 41842 27033
rect 41696 26988 41748 26994
rect 41786 26959 41842 26968
rect 42706 27024 42762 27033
rect 42706 26959 42762 26968
rect 41696 26930 41748 26936
rect 41708 26353 41736 26930
rect 41800 26926 41828 26959
rect 41788 26920 41840 26926
rect 41788 26862 41840 26868
rect 42616 26784 42668 26790
rect 42616 26726 42668 26732
rect 42708 26784 42760 26790
rect 42708 26726 42760 26732
rect 42628 26382 42656 26726
rect 42720 26586 42748 26726
rect 42812 26586 42840 27406
rect 42892 27328 42944 27334
rect 42892 27270 42944 27276
rect 42708 26580 42760 26586
rect 42708 26522 42760 26528
rect 42800 26580 42852 26586
rect 42800 26522 42852 26528
rect 42616 26376 42668 26382
rect 41694 26344 41750 26353
rect 42616 26318 42668 26324
rect 41694 26279 41750 26288
rect 42064 26240 42116 26246
rect 42064 26182 42116 26188
rect 41788 18080 41840 18086
rect 41788 18022 41840 18028
rect 41800 17610 41828 18022
rect 41788 17604 41840 17610
rect 41788 17546 41840 17552
rect 41696 17536 41748 17542
rect 41694 17504 41696 17513
rect 41748 17504 41750 17513
rect 41694 17439 41750 17448
rect 41880 17264 41932 17270
rect 41880 17206 41932 17212
rect 41788 17196 41840 17202
rect 41788 17138 41840 17144
rect 41696 17128 41748 17134
rect 41696 17070 41748 17076
rect 41708 16726 41736 17070
rect 41696 16720 41748 16726
rect 41696 16662 41748 16668
rect 41696 16584 41748 16590
rect 41696 16526 41748 16532
rect 41708 16266 41736 16526
rect 41800 16454 41828 17138
rect 41892 16590 41920 17206
rect 41880 16584 41932 16590
rect 41880 16526 41932 16532
rect 41788 16448 41840 16454
rect 41788 16390 41840 16396
rect 41708 16238 41828 16266
rect 41696 15428 41748 15434
rect 41696 15370 41748 15376
rect 41708 15026 41736 15370
rect 41696 15020 41748 15026
rect 41696 14962 41748 14968
rect 41602 14648 41658 14657
rect 41602 14583 41658 14592
rect 41328 14544 41380 14550
rect 41328 14486 41380 14492
rect 41340 13938 41368 14486
rect 41418 14240 41474 14249
rect 41418 14175 41474 14184
rect 41432 14074 41460 14175
rect 41510 14104 41566 14113
rect 41420 14068 41472 14074
rect 41510 14039 41512 14048
rect 41420 14010 41472 14016
rect 41564 14039 41566 14048
rect 41512 14010 41564 14016
rect 41708 13938 41736 14962
rect 41800 14890 41828 16238
rect 41788 14884 41840 14890
rect 41788 14826 41840 14832
rect 41972 14884 42024 14890
rect 41972 14826 42024 14832
rect 41786 14512 41842 14521
rect 41786 14447 41842 14456
rect 41328 13932 41380 13938
rect 41328 13874 41380 13880
rect 41696 13932 41748 13938
rect 41696 13874 41748 13880
rect 41052 13864 41104 13870
rect 41052 13806 41104 13812
rect 41694 13832 41750 13841
rect 41064 13734 41092 13806
rect 41694 13767 41750 13776
rect 41052 13728 41104 13734
rect 40958 13696 41014 13705
rect 41052 13670 41104 13676
rect 41144 13728 41196 13734
rect 41144 13670 41196 13676
rect 41326 13696 41382 13705
rect 40958 13631 41014 13640
rect 40972 13161 41000 13631
rect 40958 13152 41014 13161
rect 40958 13087 41014 13096
rect 40960 12912 41012 12918
rect 40960 12854 41012 12860
rect 40972 12306 41000 12854
rect 40960 12300 41012 12306
rect 40960 12242 41012 12248
rect 40960 11688 41012 11694
rect 40960 11630 41012 11636
rect 40868 11144 40920 11150
rect 40868 11086 40920 11092
rect 40776 10668 40828 10674
rect 40776 10610 40828 10616
rect 40880 9178 40908 11086
rect 40868 9172 40920 9178
rect 40868 9114 40920 9120
rect 40972 2825 41000 11630
rect 41064 11098 41092 13670
rect 41156 13190 41184 13670
rect 41326 13631 41382 13640
rect 41340 13258 41368 13631
rect 41708 13326 41736 13767
rect 41800 13530 41828 14447
rect 41880 14408 41932 14414
rect 41880 14350 41932 14356
rect 41788 13524 41840 13530
rect 41788 13466 41840 13472
rect 41512 13320 41564 13326
rect 41512 13262 41564 13268
rect 41696 13320 41748 13326
rect 41696 13262 41748 13268
rect 41328 13252 41380 13258
rect 41328 13194 41380 13200
rect 41144 13184 41196 13190
rect 41144 13126 41196 13132
rect 41524 12986 41552 13262
rect 41512 12980 41564 12986
rect 41512 12922 41564 12928
rect 41786 12880 41842 12889
rect 41512 12844 41564 12850
rect 41786 12815 41842 12824
rect 41512 12786 41564 12792
rect 41524 12753 41552 12786
rect 41510 12744 41566 12753
rect 41800 12714 41828 12815
rect 41510 12679 41566 12688
rect 41788 12708 41840 12714
rect 41788 12650 41840 12656
rect 41694 12200 41750 12209
rect 41236 12164 41288 12170
rect 41694 12135 41750 12144
rect 41236 12106 41288 12112
rect 41144 11552 41196 11558
rect 41144 11494 41196 11500
rect 41156 11354 41184 11494
rect 41248 11354 41276 12106
rect 41604 12096 41656 12102
rect 41604 12038 41656 12044
rect 41616 11830 41644 12038
rect 41604 11824 41656 11830
rect 41604 11766 41656 11772
rect 41144 11348 41196 11354
rect 41144 11290 41196 11296
rect 41236 11348 41288 11354
rect 41236 11290 41288 11296
rect 41708 11286 41736 12135
rect 41892 11370 41920 14350
rect 41984 12594 42012 14826
rect 42076 13870 42104 26182
rect 42154 22672 42210 22681
rect 42154 22607 42210 22616
rect 42168 14482 42196 22607
rect 42432 18284 42484 18290
rect 42432 18226 42484 18232
rect 42246 17776 42302 17785
rect 42246 17711 42302 17720
rect 42260 17202 42288 17711
rect 42248 17196 42300 17202
rect 42248 17138 42300 17144
rect 42156 14476 42208 14482
rect 42156 14418 42208 14424
rect 42064 13864 42116 13870
rect 42064 13806 42116 13812
rect 42156 13796 42208 13802
rect 42260 13784 42288 17138
rect 42338 17096 42394 17105
rect 42444 17066 42472 18226
rect 42800 17672 42852 17678
rect 42800 17614 42852 17620
rect 42812 17202 42840 17614
rect 42904 17270 42932 27270
rect 43456 27130 43484 27406
rect 43536 27328 43588 27334
rect 43536 27270 43588 27276
rect 43444 27124 43496 27130
rect 43444 27066 43496 27072
rect 43260 26444 43312 26450
rect 43260 26386 43312 26392
rect 43272 25838 43300 26386
rect 43260 25832 43312 25838
rect 43260 25774 43312 25780
rect 42892 17264 42944 17270
rect 42892 17206 42944 17212
rect 42800 17196 42852 17202
rect 42800 17138 42852 17144
rect 43076 17128 43128 17134
rect 43076 17070 43128 17076
rect 42338 17031 42394 17040
rect 42432 17060 42484 17066
rect 42352 16833 42380 17031
rect 42432 17002 42484 17008
rect 42338 16824 42394 16833
rect 42338 16759 42394 16768
rect 42352 15502 42380 16759
rect 42984 16720 43036 16726
rect 42982 16688 42984 16697
rect 43036 16688 43038 16697
rect 42982 16623 43038 16632
rect 42708 16584 42760 16590
rect 42708 16526 42760 16532
rect 42616 16108 42668 16114
rect 42616 16050 42668 16056
rect 42628 15745 42656 16050
rect 42614 15736 42670 15745
rect 42614 15671 42670 15680
rect 42720 15502 42748 16526
rect 43088 16250 43116 17070
rect 43168 16448 43220 16454
rect 43168 16390 43220 16396
rect 43180 16250 43208 16390
rect 43076 16244 43128 16250
rect 43076 16186 43128 16192
rect 43168 16244 43220 16250
rect 43168 16186 43220 16192
rect 42892 16108 42944 16114
rect 42892 16050 42944 16056
rect 42984 16108 43036 16114
rect 42984 16050 43036 16056
rect 42904 15881 42932 16050
rect 42996 15978 43024 16050
rect 42984 15972 43036 15978
rect 42984 15914 43036 15920
rect 42890 15872 42946 15881
rect 42890 15807 42946 15816
rect 42340 15496 42392 15502
rect 42340 15438 42392 15444
rect 42708 15496 42760 15502
rect 42708 15438 42760 15444
rect 42432 15360 42484 15366
rect 42432 15302 42484 15308
rect 42444 15162 42472 15302
rect 42432 15156 42484 15162
rect 42432 15098 42484 15104
rect 42720 14006 42748 15438
rect 43076 14952 43128 14958
rect 42798 14920 42854 14929
rect 43076 14894 43128 14900
rect 42798 14855 42854 14864
rect 42812 14550 42840 14855
rect 42892 14816 42944 14822
rect 42890 14784 42892 14793
rect 42944 14784 42946 14793
rect 42890 14719 42946 14728
rect 42800 14544 42852 14550
rect 42800 14486 42852 14492
rect 42984 14272 43036 14278
rect 42984 14214 43036 14220
rect 42524 14000 42576 14006
rect 42524 13942 42576 13948
rect 42708 14000 42760 14006
rect 42708 13942 42760 13948
rect 42208 13756 42288 13784
rect 42156 13738 42208 13744
rect 41984 12566 42104 12594
rect 41800 11342 41920 11370
rect 41696 11280 41748 11286
rect 41142 11248 41198 11257
rect 41696 11222 41748 11228
rect 41142 11183 41144 11192
rect 41196 11183 41198 11192
rect 41328 11212 41380 11218
rect 41144 11154 41196 11160
rect 41328 11154 41380 11160
rect 41064 11070 41276 11098
rect 41340 11082 41368 11154
rect 41800 11150 41828 11342
rect 41880 11280 41932 11286
rect 41880 11222 41932 11228
rect 41788 11144 41840 11150
rect 41788 11086 41840 11092
rect 41892 11082 41920 11222
rect 41972 11144 42024 11150
rect 41972 11086 42024 11092
rect 41052 11008 41104 11014
rect 41144 11008 41196 11014
rect 41052 10950 41104 10956
rect 41142 10976 41144 10985
rect 41196 10976 41198 10985
rect 41064 10538 41092 10950
rect 41142 10911 41198 10920
rect 41052 10532 41104 10538
rect 41052 10474 41104 10480
rect 41248 4826 41276 11070
rect 41328 11076 41380 11082
rect 41328 11018 41380 11024
rect 41880 11076 41932 11082
rect 41880 11018 41932 11024
rect 41420 10668 41472 10674
rect 41420 10610 41472 10616
rect 41432 10577 41460 10610
rect 41418 10568 41474 10577
rect 41418 10503 41474 10512
rect 41984 10198 42012 11086
rect 41972 10192 42024 10198
rect 41972 10134 42024 10140
rect 41696 9988 41748 9994
rect 41696 9930 41748 9936
rect 41708 9382 41736 9930
rect 41696 9376 41748 9382
rect 41696 9318 41748 9324
rect 41328 9172 41380 9178
rect 41328 9114 41380 9120
rect 41340 8498 41368 9114
rect 41328 8492 41380 8498
rect 41328 8434 41380 8440
rect 41420 8424 41472 8430
rect 41420 8366 41472 8372
rect 41236 4820 41288 4826
rect 41236 4762 41288 4768
rect 41432 3602 41460 8366
rect 41420 3596 41472 3602
rect 41420 3538 41472 3544
rect 41236 3460 41288 3466
rect 41236 3402 41288 3408
rect 40328 2746 40448 2774
rect 40512 2746 40724 2774
rect 40958 2816 41014 2825
rect 40958 2751 41014 2760
rect 40328 2145 40356 2746
rect 40512 2514 40540 2746
rect 40500 2508 40552 2514
rect 40500 2450 40552 2456
rect 40592 2304 40644 2310
rect 40592 2246 40644 2252
rect 40314 2136 40370 2145
rect 40314 2071 40370 2080
rect 40604 800 40632 2246
rect 41248 800 41276 3402
rect 41604 3120 41656 3126
rect 41604 3062 41656 3068
rect 41616 2922 41644 3062
rect 41604 2916 41656 2922
rect 41604 2858 41656 2864
rect 41708 2378 41736 9318
rect 42076 8430 42104 12566
rect 42168 10305 42196 13738
rect 42432 13524 42484 13530
rect 42432 13466 42484 13472
rect 42248 13320 42300 13326
rect 42248 13262 42300 13268
rect 42260 12918 42288 13262
rect 42340 13184 42392 13190
rect 42340 13126 42392 13132
rect 42248 12912 42300 12918
rect 42248 12854 42300 12860
rect 42248 12640 42300 12646
rect 42248 12582 42300 12588
rect 42260 12442 42288 12582
rect 42248 12436 42300 12442
rect 42248 12378 42300 12384
rect 42248 11212 42300 11218
rect 42248 11154 42300 11160
rect 42154 10296 42210 10305
rect 42260 10266 42288 11154
rect 42352 11150 42380 13126
rect 42444 12850 42472 13466
rect 42432 12844 42484 12850
rect 42536 12832 42564 13942
rect 42720 13258 42748 13942
rect 42996 13938 43024 14214
rect 42984 13932 43036 13938
rect 42984 13874 43036 13880
rect 42892 13864 42944 13870
rect 42892 13806 42944 13812
rect 42904 13569 42932 13806
rect 42890 13560 42946 13569
rect 42890 13495 42946 13504
rect 42984 13524 43036 13530
rect 42800 13320 42852 13326
rect 42800 13262 42852 13268
rect 42708 13252 42760 13258
rect 42708 13194 42760 13200
rect 42812 12889 42840 13262
rect 42904 12918 42932 13495
rect 43088 13512 43116 14894
rect 43168 13796 43220 13802
rect 43168 13738 43220 13744
rect 43036 13484 43116 13512
rect 42984 13466 43036 13472
rect 43088 13258 43116 13484
rect 43076 13252 43128 13258
rect 43076 13194 43128 13200
rect 42892 12912 42944 12918
rect 42798 12880 42854 12889
rect 42616 12844 42668 12850
rect 42536 12804 42616 12832
rect 42432 12786 42484 12792
rect 42892 12854 42944 12860
rect 42798 12815 42854 12824
rect 42616 12786 42668 12792
rect 42984 12776 43036 12782
rect 42984 12718 43036 12724
rect 42996 12238 43024 12718
rect 42984 12232 43036 12238
rect 42984 12174 43036 12180
rect 43180 12170 43208 13738
rect 43168 12164 43220 12170
rect 43168 12106 43220 12112
rect 43076 11212 43128 11218
rect 43076 11154 43128 11160
rect 42340 11144 42392 11150
rect 42340 11086 42392 11092
rect 42628 10662 43024 10690
rect 43088 10674 43116 11154
rect 42628 10606 42656 10662
rect 42616 10600 42668 10606
rect 42616 10542 42668 10548
rect 42996 10538 43024 10662
rect 43076 10668 43128 10674
rect 43076 10610 43128 10616
rect 42892 10532 42944 10538
rect 42892 10474 42944 10480
rect 42984 10532 43036 10538
rect 42984 10474 43036 10480
rect 42432 10464 42484 10470
rect 42432 10406 42484 10412
rect 42154 10231 42210 10240
rect 42248 10260 42300 10266
rect 42248 10202 42300 10208
rect 42444 10146 42472 10406
rect 42904 10266 42932 10474
rect 42892 10260 42944 10266
rect 42892 10202 42944 10208
rect 42444 10118 42840 10146
rect 42812 10062 42840 10118
rect 42800 10056 42852 10062
rect 42800 9998 42852 10004
rect 42708 9988 42760 9994
rect 42708 9930 42760 9936
rect 42720 9042 42748 9930
rect 42904 9586 42932 10202
rect 42984 9920 43036 9926
rect 42984 9862 43036 9868
rect 42892 9580 42944 9586
rect 42892 9522 42944 9528
rect 42996 9518 43024 9862
rect 42984 9512 43036 9518
rect 42984 9454 43036 9460
rect 42708 9036 42760 9042
rect 42708 8978 42760 8984
rect 42800 8968 42852 8974
rect 42800 8910 42852 8916
rect 42812 8634 42840 8910
rect 42800 8628 42852 8634
rect 42800 8570 42852 8576
rect 42064 8424 42116 8430
rect 42064 8366 42116 8372
rect 41880 8288 41932 8294
rect 41880 8230 41932 8236
rect 41892 7886 41920 8230
rect 41880 7880 41932 7886
rect 41880 7822 41932 7828
rect 41972 7744 42024 7750
rect 41972 7686 42024 7692
rect 41880 3664 41932 3670
rect 41880 3606 41932 3612
rect 41892 3398 41920 3606
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 41984 2446 42012 7686
rect 42614 3768 42670 3777
rect 42614 3703 42616 3712
rect 42668 3703 42670 3712
rect 42708 3732 42760 3738
rect 42616 3674 42668 3680
rect 42708 3674 42760 3680
rect 42720 3602 42748 3674
rect 42708 3596 42760 3602
rect 42708 3538 42760 3544
rect 43272 3126 43300 25774
rect 43548 18426 43576 27270
rect 44008 21418 44036 27406
rect 44846 27228 45154 27237
rect 44846 27226 44852 27228
rect 44908 27226 44932 27228
rect 44988 27226 45012 27228
rect 45068 27226 45092 27228
rect 45148 27226 45154 27228
rect 44908 27174 44910 27226
rect 45090 27174 45092 27226
rect 44846 27172 44852 27174
rect 44908 27172 44932 27174
rect 44988 27172 45012 27174
rect 45068 27172 45092 27174
rect 45148 27172 45154 27174
rect 44846 27163 45154 27172
rect 45284 27124 45336 27130
rect 45284 27066 45336 27072
rect 44822 27024 44878 27033
rect 44180 26988 44232 26994
rect 44180 26930 44232 26936
rect 44732 26988 44784 26994
rect 44822 26959 44824 26968
rect 44732 26930 44784 26936
rect 44876 26959 44878 26968
rect 44824 26930 44876 26936
rect 43996 21412 44048 21418
rect 43996 21354 44048 21360
rect 43536 18420 43588 18426
rect 43536 18362 43588 18368
rect 43442 17776 43498 17785
rect 43442 17711 43444 17720
rect 43496 17711 43498 17720
rect 43444 17682 43496 17688
rect 43352 17672 43404 17678
rect 43352 17614 43404 17620
rect 43364 16998 43392 17614
rect 43628 17196 43680 17202
rect 43680 17156 43852 17184
rect 43628 17138 43680 17144
rect 43824 17066 43852 17156
rect 43812 17060 43864 17066
rect 43812 17002 43864 17008
rect 43352 16992 43404 16998
rect 43628 16992 43680 16998
rect 43404 16952 43484 16980
rect 43352 16934 43404 16940
rect 43352 16448 43404 16454
rect 43352 16390 43404 16396
rect 43364 16182 43392 16390
rect 43352 16176 43404 16182
rect 43352 16118 43404 16124
rect 43456 14958 43484 16952
rect 43628 16934 43680 16940
rect 43640 16114 43668 16934
rect 43628 16108 43680 16114
rect 43628 16050 43680 16056
rect 43904 16108 43956 16114
rect 43904 16050 43956 16056
rect 43996 16108 44048 16114
rect 43996 16050 44048 16056
rect 43916 15881 43944 16050
rect 43902 15872 43958 15881
rect 43902 15807 43958 15816
rect 44008 15706 44036 16050
rect 43996 15700 44048 15706
rect 43996 15642 44048 15648
rect 44088 15428 44140 15434
rect 44088 15370 44140 15376
rect 44100 14958 44128 15370
rect 43444 14952 43496 14958
rect 43444 14894 43496 14900
rect 44088 14952 44140 14958
rect 44088 14894 44140 14900
rect 44088 14816 44140 14822
rect 44088 14758 44140 14764
rect 43902 14648 43958 14657
rect 43902 14583 43958 14592
rect 43536 14476 43588 14482
rect 43536 14418 43588 14424
rect 43444 13184 43496 13190
rect 43444 13126 43496 13132
rect 43456 13025 43484 13126
rect 43442 13016 43498 13025
rect 43442 12951 43498 12960
rect 43352 12300 43404 12306
rect 43352 12242 43404 12248
rect 43364 11937 43392 12242
rect 43350 11928 43406 11937
rect 43350 11863 43406 11872
rect 43364 10169 43392 11863
rect 43548 10470 43576 14418
rect 43916 14414 43944 14583
rect 43904 14408 43956 14414
rect 43732 14368 43904 14396
rect 43628 14340 43680 14346
rect 43628 14282 43680 14288
rect 43640 13530 43668 14282
rect 43628 13524 43680 13530
rect 43628 13466 43680 13472
rect 43732 12646 43760 14368
rect 43904 14350 43956 14356
rect 43996 14408 44048 14414
rect 43996 14350 44048 14356
rect 44008 14260 44036 14350
rect 43824 14232 44036 14260
rect 43824 13705 43852 14232
rect 43810 13696 43866 13705
rect 43810 13631 43866 13640
rect 43824 12782 43852 13631
rect 44100 13569 44128 14758
rect 44192 14550 44220 26930
rect 44744 26042 44772 26930
rect 44824 26852 44876 26858
rect 44824 26794 44876 26800
rect 44836 26450 44864 26794
rect 44824 26444 44876 26450
rect 44824 26386 44876 26392
rect 45296 26382 45324 27066
rect 45388 26382 45416 27406
rect 45284 26376 45336 26382
rect 45284 26318 45336 26324
rect 45376 26376 45428 26382
rect 45376 26318 45428 26324
rect 44846 26140 45154 26149
rect 44846 26138 44852 26140
rect 44908 26138 44932 26140
rect 44988 26138 45012 26140
rect 45068 26138 45092 26140
rect 45148 26138 45154 26140
rect 44908 26086 44910 26138
rect 45090 26086 45092 26138
rect 44846 26084 44852 26086
rect 44908 26084 44932 26086
rect 44988 26084 45012 26086
rect 45068 26084 45092 26086
rect 45148 26084 45154 26086
rect 44846 26075 45154 26084
rect 44732 26036 44784 26042
rect 44732 25978 44784 25984
rect 44640 25900 44692 25906
rect 44640 25842 44692 25848
rect 44548 18284 44600 18290
rect 44548 18226 44600 18232
rect 44272 18216 44324 18222
rect 44272 18158 44324 18164
rect 44284 17678 44312 18158
rect 44560 17814 44588 18226
rect 44548 17808 44600 17814
rect 44548 17750 44600 17756
rect 44272 17672 44324 17678
rect 44272 17614 44324 17620
rect 44456 15904 44508 15910
rect 44456 15846 44508 15852
rect 44270 15600 44326 15609
rect 44270 15535 44326 15544
rect 44284 15366 44312 15535
rect 44272 15360 44324 15366
rect 44272 15302 44324 15308
rect 44364 15360 44416 15366
rect 44364 15302 44416 15308
rect 44376 15026 44404 15302
rect 44364 15020 44416 15026
rect 44364 14962 44416 14968
rect 44468 15008 44496 15846
rect 44652 15201 44680 25842
rect 44846 25052 45154 25061
rect 44846 25050 44852 25052
rect 44908 25050 44932 25052
rect 44988 25050 45012 25052
rect 45068 25050 45092 25052
rect 45148 25050 45154 25052
rect 44908 24998 44910 25050
rect 45090 24998 45092 25050
rect 44846 24996 44852 24998
rect 44908 24996 44932 24998
rect 44988 24996 45012 24998
rect 45068 24996 45092 24998
rect 45148 24996 45154 24998
rect 44846 24987 45154 24996
rect 44846 23964 45154 23973
rect 44846 23962 44852 23964
rect 44908 23962 44932 23964
rect 44988 23962 45012 23964
rect 45068 23962 45092 23964
rect 45148 23962 45154 23964
rect 44908 23910 44910 23962
rect 45090 23910 45092 23962
rect 44846 23908 44852 23910
rect 44908 23908 44932 23910
rect 44988 23908 45012 23910
rect 45068 23908 45092 23910
rect 45148 23908 45154 23910
rect 44846 23899 45154 23908
rect 44846 22876 45154 22885
rect 44846 22874 44852 22876
rect 44908 22874 44932 22876
rect 44988 22874 45012 22876
rect 45068 22874 45092 22876
rect 45148 22874 45154 22876
rect 44908 22822 44910 22874
rect 45090 22822 45092 22874
rect 44846 22820 44852 22822
rect 44908 22820 44932 22822
rect 44988 22820 45012 22822
rect 45068 22820 45092 22822
rect 45148 22820 45154 22822
rect 44846 22811 45154 22820
rect 44846 21788 45154 21797
rect 44846 21786 44852 21788
rect 44908 21786 44932 21788
rect 44988 21786 45012 21788
rect 45068 21786 45092 21788
rect 45148 21786 45154 21788
rect 44908 21734 44910 21786
rect 45090 21734 45092 21786
rect 44846 21732 44852 21734
rect 44908 21732 44932 21734
rect 44988 21732 45012 21734
rect 45068 21732 45092 21734
rect 45148 21732 45154 21734
rect 44846 21723 45154 21732
rect 44846 20700 45154 20709
rect 44846 20698 44852 20700
rect 44908 20698 44932 20700
rect 44988 20698 45012 20700
rect 45068 20698 45092 20700
rect 45148 20698 45154 20700
rect 44908 20646 44910 20698
rect 45090 20646 45092 20698
rect 44846 20644 44852 20646
rect 44908 20644 44932 20646
rect 44988 20644 45012 20646
rect 45068 20644 45092 20646
rect 45148 20644 45154 20646
rect 44846 20635 45154 20644
rect 44846 19612 45154 19621
rect 44846 19610 44852 19612
rect 44908 19610 44932 19612
rect 44988 19610 45012 19612
rect 45068 19610 45092 19612
rect 45148 19610 45154 19612
rect 44908 19558 44910 19610
rect 45090 19558 45092 19610
rect 44846 19556 44852 19558
rect 44908 19556 44932 19558
rect 44988 19556 45012 19558
rect 45068 19556 45092 19558
rect 45148 19556 45154 19558
rect 44846 19547 45154 19556
rect 44846 18524 45154 18533
rect 44846 18522 44852 18524
rect 44908 18522 44932 18524
rect 44988 18522 45012 18524
rect 45068 18522 45092 18524
rect 45148 18522 45154 18524
rect 44908 18470 44910 18522
rect 45090 18470 45092 18522
rect 44846 18468 44852 18470
rect 44908 18468 44932 18470
rect 44988 18468 45012 18470
rect 45068 18468 45092 18470
rect 45148 18468 45154 18470
rect 44846 18459 45154 18468
rect 45192 18080 45244 18086
rect 45192 18022 45244 18028
rect 44846 17436 45154 17445
rect 44846 17434 44852 17436
rect 44908 17434 44932 17436
rect 44988 17434 45012 17436
rect 45068 17434 45092 17436
rect 45148 17434 45154 17436
rect 44908 17382 44910 17434
rect 45090 17382 45092 17434
rect 44846 17380 44852 17382
rect 44908 17380 44932 17382
rect 44988 17380 45012 17382
rect 45068 17380 45092 17382
rect 45148 17380 45154 17382
rect 44846 17371 45154 17380
rect 44732 17264 44784 17270
rect 44732 17206 44784 17212
rect 44744 16697 44772 17206
rect 45100 17196 45152 17202
rect 45204 17184 45232 18022
rect 45480 17814 45508 27406
rect 46676 26246 46704 27406
rect 48596 27406 48648 27412
rect 49056 27464 49108 27470
rect 49056 27406 49108 27412
rect 46754 27367 46756 27376
rect 46808 27367 46810 27376
rect 46756 27338 46808 27344
rect 48320 27328 48372 27334
rect 48320 27270 48372 27276
rect 46664 26240 46716 26246
rect 46664 26182 46716 26188
rect 48228 18828 48280 18834
rect 48228 18770 48280 18776
rect 48044 18760 48096 18766
rect 48044 18702 48096 18708
rect 47676 18624 47728 18630
rect 47676 18566 47728 18572
rect 46204 18352 46256 18358
rect 46204 18294 46256 18300
rect 45650 17912 45706 17921
rect 46216 17882 46244 18294
rect 45650 17847 45706 17856
rect 46204 17876 46256 17882
rect 45468 17808 45520 17814
rect 45468 17750 45520 17756
rect 45664 17678 45692 17847
rect 46204 17818 46256 17824
rect 46296 17876 46348 17882
rect 46296 17818 46348 17824
rect 46308 17785 46336 17818
rect 46294 17776 46350 17785
rect 46294 17711 46350 17720
rect 45652 17672 45704 17678
rect 45652 17614 45704 17620
rect 45928 17672 45980 17678
rect 46940 17672 46992 17678
rect 45928 17614 45980 17620
rect 46294 17640 46350 17649
rect 45664 17377 45692 17614
rect 45650 17368 45706 17377
rect 45650 17303 45706 17312
rect 45744 17264 45796 17270
rect 45744 17206 45796 17212
rect 45152 17156 45232 17184
rect 45100 17138 45152 17144
rect 44824 17060 44876 17066
rect 44824 17002 44876 17008
rect 44730 16688 44786 16697
rect 44730 16623 44786 16632
rect 44732 16516 44784 16522
rect 44732 16458 44784 16464
rect 44744 16114 44772 16458
rect 44836 16454 44864 17002
rect 44824 16448 44876 16454
rect 44824 16390 44876 16396
rect 44846 16348 45154 16357
rect 44846 16346 44852 16348
rect 44908 16346 44932 16348
rect 44988 16346 45012 16348
rect 45068 16346 45092 16348
rect 45148 16346 45154 16348
rect 44908 16294 44910 16346
rect 45090 16294 45092 16346
rect 44846 16292 44852 16294
rect 44908 16292 44932 16294
rect 44988 16292 45012 16294
rect 45068 16292 45092 16294
rect 45148 16292 45154 16294
rect 44846 16283 45154 16292
rect 44732 16108 44784 16114
rect 44732 16050 44784 16056
rect 45008 16108 45060 16114
rect 45008 16050 45060 16056
rect 45376 16108 45428 16114
rect 45376 16050 45428 16056
rect 45020 15706 45048 16050
rect 45388 15706 45416 16050
rect 45652 15904 45704 15910
rect 45652 15846 45704 15852
rect 45008 15700 45060 15706
rect 45008 15642 45060 15648
rect 45376 15700 45428 15706
rect 45376 15642 45428 15648
rect 45664 15502 45692 15846
rect 45756 15570 45784 17206
rect 45940 16969 45968 17614
rect 46754 17640 46810 17649
rect 46294 17575 46350 17584
rect 46572 17604 46624 17610
rect 46308 17066 46336 17575
rect 46940 17614 46992 17620
rect 47216 17672 47268 17678
rect 47268 17632 47348 17660
rect 47216 17614 47268 17620
rect 46754 17575 46810 17584
rect 46572 17546 46624 17552
rect 46584 17202 46612 17546
rect 46768 17202 46796 17575
rect 46572 17196 46624 17202
rect 46572 17138 46624 17144
rect 46756 17196 46808 17202
rect 46756 17138 46808 17144
rect 46296 17060 46348 17066
rect 46296 17002 46348 17008
rect 45926 16960 45982 16969
rect 45926 16895 45982 16904
rect 45940 16726 45968 16895
rect 45928 16720 45980 16726
rect 45928 16662 45980 16668
rect 46768 16590 46796 17138
rect 46848 16992 46900 16998
rect 46848 16934 46900 16940
rect 46860 16590 46888 16934
rect 46952 16726 46980 17614
rect 47032 17196 47084 17202
rect 47032 17138 47084 17144
rect 46940 16720 46992 16726
rect 46940 16662 46992 16668
rect 47044 16658 47072 17138
rect 47032 16652 47084 16658
rect 47032 16594 47084 16600
rect 46756 16584 46808 16590
rect 46756 16526 46808 16532
rect 46848 16584 46900 16590
rect 46848 16526 46900 16532
rect 47216 16584 47268 16590
rect 47216 16526 47268 16532
rect 47124 16516 47176 16522
rect 47124 16458 47176 16464
rect 46664 16448 46716 16454
rect 46202 16416 46258 16425
rect 46664 16390 46716 16396
rect 46202 16351 46258 16360
rect 45928 16176 45980 16182
rect 45928 16118 45980 16124
rect 45744 15564 45796 15570
rect 45744 15506 45796 15512
rect 45100 15496 45152 15502
rect 45100 15438 45152 15444
rect 45376 15496 45428 15502
rect 45376 15438 45428 15444
rect 45652 15496 45704 15502
rect 45652 15438 45704 15444
rect 45112 15366 45140 15438
rect 45100 15360 45152 15366
rect 45100 15302 45152 15308
rect 44846 15260 45154 15269
rect 44846 15258 44852 15260
rect 44908 15258 44932 15260
rect 44988 15258 45012 15260
rect 45068 15258 45092 15260
rect 45148 15258 45154 15260
rect 44908 15206 44910 15258
rect 45090 15206 45092 15258
rect 44846 15204 44852 15206
rect 44908 15204 44932 15206
rect 44988 15204 45012 15206
rect 45068 15204 45092 15206
rect 45148 15204 45154 15206
rect 44638 15192 44694 15201
rect 44846 15195 45154 15204
rect 44638 15127 44694 15136
rect 44548 15020 44600 15026
rect 44468 14980 44548 15008
rect 44180 14544 44232 14550
rect 44180 14486 44232 14492
rect 44364 13932 44416 13938
rect 44364 13874 44416 13880
rect 44086 13560 44142 13569
rect 44376 13530 44404 13874
rect 44468 13818 44496 14980
rect 44548 14962 44600 14968
rect 44548 14408 44600 14414
rect 44548 14350 44600 14356
rect 44560 14249 44588 14350
rect 44546 14240 44602 14249
rect 44546 14175 44602 14184
rect 44560 13938 44588 14175
rect 44548 13932 44600 13938
rect 44548 13874 44600 13880
rect 44468 13790 44588 13818
rect 44086 13495 44142 13504
rect 44364 13524 44416 13530
rect 44364 13466 44416 13472
rect 44456 13524 44508 13530
rect 44456 13466 44508 13472
rect 44272 13388 44324 13394
rect 44272 13330 44324 13336
rect 43902 13152 43958 13161
rect 43902 13087 43958 13096
rect 43916 12782 43944 13087
rect 43996 12844 44048 12850
rect 43996 12786 44048 12792
rect 43812 12776 43864 12782
rect 43812 12718 43864 12724
rect 43904 12776 43956 12782
rect 43904 12718 43956 12724
rect 43720 12640 43772 12646
rect 43720 12582 43772 12588
rect 43904 12640 43956 12646
rect 43904 12582 43956 12588
rect 43626 12336 43682 12345
rect 43626 12271 43682 12280
rect 43640 11694 43668 12271
rect 43812 12096 43864 12102
rect 43812 12038 43864 12044
rect 43824 11898 43852 12038
rect 43812 11892 43864 11898
rect 43812 11834 43864 11840
rect 43720 11824 43772 11830
rect 43720 11766 43772 11772
rect 43628 11688 43680 11694
rect 43628 11630 43680 11636
rect 43732 11529 43760 11766
rect 43718 11520 43774 11529
rect 43718 11455 43774 11464
rect 43718 11248 43774 11257
rect 43718 11183 43774 11192
rect 43444 10464 43496 10470
rect 43444 10406 43496 10412
rect 43536 10464 43588 10470
rect 43536 10406 43588 10412
rect 43350 10160 43406 10169
rect 43350 10095 43406 10104
rect 43456 9926 43484 10406
rect 43444 9920 43496 9926
rect 43444 9862 43496 9868
rect 43548 8498 43576 10406
rect 43536 8492 43588 8498
rect 43536 8434 43588 8440
rect 43442 4040 43498 4049
rect 43442 3975 43444 3984
rect 43496 3975 43498 3984
rect 43444 3946 43496 3952
rect 43444 3528 43496 3534
rect 43442 3496 43444 3505
rect 43496 3496 43498 3505
rect 43442 3431 43498 3440
rect 43260 3120 43312 3126
rect 43260 3062 43312 3068
rect 43272 2854 43300 3062
rect 43444 2916 43496 2922
rect 43444 2858 43496 2864
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 43260 2848 43312 2854
rect 43260 2790 43312 2796
rect 42812 2446 42840 2790
rect 43456 2446 43484 2858
rect 43732 2582 43760 11183
rect 43916 3058 43944 12582
rect 44008 12322 44036 12786
rect 44088 12776 44140 12782
rect 44088 12718 44140 12724
rect 44100 12442 44128 12718
rect 44088 12436 44140 12442
rect 44088 12378 44140 12384
rect 44180 12436 44232 12442
rect 44180 12378 44232 12384
rect 44192 12322 44220 12378
rect 44008 12294 44220 12322
rect 44008 12073 44036 12294
rect 43994 12064 44050 12073
rect 43994 11999 44050 12008
rect 44180 11756 44232 11762
rect 44180 11698 44232 11704
rect 44088 11620 44140 11626
rect 44088 11562 44140 11568
rect 44100 11286 44128 11562
rect 44192 11558 44220 11698
rect 44180 11552 44232 11558
rect 44180 11494 44232 11500
rect 44088 11280 44140 11286
rect 44088 11222 44140 11228
rect 44284 11150 44312 13330
rect 44364 12232 44416 12238
rect 44468 12220 44496 13466
rect 44416 12192 44496 12220
rect 44364 12174 44416 12180
rect 44364 11756 44416 11762
rect 44364 11698 44416 11704
rect 44376 11257 44404 11698
rect 44456 11552 44508 11558
rect 44456 11494 44508 11500
rect 44362 11248 44418 11257
rect 44362 11183 44418 11192
rect 44272 11144 44324 11150
rect 44272 11086 44324 11092
rect 44364 11144 44416 11150
rect 44468 11098 44496 11494
rect 44416 11092 44496 11098
rect 44364 11086 44496 11092
rect 44376 11070 44496 11086
rect 43996 10600 44048 10606
rect 43996 10542 44048 10548
rect 44008 9450 44036 10542
rect 44088 9580 44140 9586
rect 44088 9522 44140 9528
rect 43996 9444 44048 9450
rect 43996 9386 44048 9392
rect 44100 9178 44128 9522
rect 44088 9172 44140 9178
rect 44088 9114 44140 9120
rect 44100 8634 44128 9114
rect 44088 8628 44140 8634
rect 44088 8570 44140 8576
rect 44376 4146 44404 11070
rect 44456 10464 44508 10470
rect 44456 10406 44508 10412
rect 44468 10266 44496 10406
rect 44456 10260 44508 10266
rect 44456 10202 44508 10208
rect 44560 5234 44588 13790
rect 44652 13530 44680 15127
rect 45020 14618 45232 14634
rect 45008 14612 45244 14618
rect 45060 14606 45192 14612
rect 45008 14554 45060 14560
rect 45192 14554 45244 14560
rect 45284 14544 45336 14550
rect 44836 14492 45284 14498
rect 44836 14486 45336 14492
rect 44836 14482 45324 14486
rect 44824 14476 45324 14482
rect 44876 14470 45324 14476
rect 44824 14418 44876 14424
rect 45284 14408 45336 14414
rect 45204 14368 45284 14396
rect 44846 14172 45154 14181
rect 44846 14170 44852 14172
rect 44908 14170 44932 14172
rect 44988 14170 45012 14172
rect 45068 14170 45092 14172
rect 45148 14170 45154 14172
rect 44908 14118 44910 14170
rect 45090 14118 45092 14170
rect 44846 14116 44852 14118
rect 44908 14116 44932 14118
rect 44988 14116 45012 14118
rect 45068 14116 45092 14118
rect 45148 14116 45154 14118
rect 44846 14107 45154 14116
rect 45204 13870 45232 14368
rect 45284 14350 45336 14356
rect 45282 14104 45338 14113
rect 45282 14039 45338 14048
rect 45192 13864 45244 13870
rect 45192 13806 45244 13812
rect 45100 13728 45152 13734
rect 45100 13670 45152 13676
rect 44730 13560 44786 13569
rect 44640 13524 44692 13530
rect 45112 13530 45140 13670
rect 44730 13495 44786 13504
rect 45100 13524 45152 13530
rect 44640 13466 44692 13472
rect 44744 12850 44772 13495
rect 45100 13466 45152 13472
rect 45296 13462 45324 14039
rect 45284 13456 45336 13462
rect 45284 13398 45336 13404
rect 44846 13084 45154 13093
rect 44846 13082 44852 13084
rect 44908 13082 44932 13084
rect 44988 13082 45012 13084
rect 45068 13082 45092 13084
rect 45148 13082 45154 13084
rect 44908 13030 44910 13082
rect 45090 13030 45092 13082
rect 44846 13028 44852 13030
rect 44908 13028 44932 13030
rect 44988 13028 45012 13030
rect 45068 13028 45092 13030
rect 45148 13028 45154 13030
rect 44846 13019 45154 13028
rect 45282 12880 45338 12889
rect 44732 12844 44784 12850
rect 44732 12786 44784 12792
rect 44824 12844 44876 12850
rect 45282 12815 45338 12824
rect 44824 12786 44876 12792
rect 44640 12640 44692 12646
rect 44640 12582 44692 12588
rect 44652 11898 44680 12582
rect 44836 12084 44864 12786
rect 45296 12782 45324 12815
rect 45284 12776 45336 12782
rect 45284 12718 45336 12724
rect 45388 12434 45416 15438
rect 45652 14952 45704 14958
rect 45652 14894 45704 14900
rect 45560 14816 45612 14822
rect 45560 14758 45612 14764
rect 45572 14550 45600 14758
rect 45560 14544 45612 14550
rect 45560 14486 45612 14492
rect 45558 13560 45614 13569
rect 45558 13495 45614 13504
rect 45468 13388 45520 13394
rect 45468 13330 45520 13336
rect 45480 13025 45508 13330
rect 45466 13016 45522 13025
rect 45466 12951 45522 12960
rect 45468 12776 45520 12782
rect 45468 12718 45520 12724
rect 44744 12056 44864 12084
rect 45204 12406 45416 12434
rect 44744 11898 44772 12056
rect 44846 11996 45154 12005
rect 44846 11994 44852 11996
rect 44908 11994 44932 11996
rect 44988 11994 45012 11996
rect 45068 11994 45092 11996
rect 45148 11994 45154 11996
rect 44908 11942 44910 11994
rect 45090 11942 45092 11994
rect 44846 11940 44852 11942
rect 44908 11940 44932 11942
rect 44988 11940 45012 11942
rect 45068 11940 45092 11942
rect 45148 11940 45154 11942
rect 44846 11931 45154 11940
rect 44640 11892 44692 11898
rect 44640 11834 44692 11840
rect 44732 11892 44784 11898
rect 44732 11834 44784 11840
rect 44744 11354 44772 11834
rect 44824 11824 44876 11830
rect 44824 11766 44876 11772
rect 45100 11824 45152 11830
rect 45100 11766 45152 11772
rect 44732 11348 44784 11354
rect 44732 11290 44784 11296
rect 44836 11121 44864 11766
rect 45112 11354 45140 11766
rect 45100 11348 45152 11354
rect 45100 11290 45152 11296
rect 44822 11112 44878 11121
rect 44640 11076 44692 11082
rect 44822 11047 44878 11056
rect 44640 11018 44692 11024
rect 44652 10538 44680 11018
rect 44846 10908 45154 10917
rect 44846 10906 44852 10908
rect 44908 10906 44932 10908
rect 44988 10906 45012 10908
rect 45068 10906 45092 10908
rect 45148 10906 45154 10908
rect 44908 10854 44910 10906
rect 45090 10854 45092 10906
rect 44846 10852 44852 10854
rect 44908 10852 44932 10854
rect 44988 10852 45012 10854
rect 45068 10852 45092 10854
rect 45148 10852 45154 10854
rect 44846 10843 45154 10852
rect 45204 10690 45232 12406
rect 45480 12306 45508 12718
rect 45572 12646 45600 13495
rect 45664 13258 45692 14894
rect 45756 14890 45784 15506
rect 45940 15366 45968 16118
rect 46216 16114 46244 16351
rect 46676 16289 46704 16390
rect 46662 16280 46718 16289
rect 46662 16215 46718 16224
rect 46480 16176 46532 16182
rect 46386 16144 46442 16153
rect 46204 16108 46256 16114
rect 46848 16176 46900 16182
rect 46532 16136 46796 16164
rect 46480 16118 46532 16124
rect 46386 16079 46388 16088
rect 46204 16050 46256 16056
rect 46440 16079 46442 16088
rect 46388 16050 46440 16056
rect 46664 15904 46716 15910
rect 46664 15846 46716 15852
rect 46676 15706 46704 15846
rect 46768 15706 46796 16136
rect 46848 16118 46900 16124
rect 46860 15881 46888 16118
rect 47136 16114 47164 16458
rect 47124 16108 47176 16114
rect 47124 16050 47176 16056
rect 47228 15978 47256 16526
rect 47320 16522 47348 17632
rect 47400 17536 47452 17542
rect 47400 17478 47452 17484
rect 47412 16590 47440 17478
rect 47688 17202 47716 18566
rect 48056 18426 48084 18702
rect 48240 18426 48268 18770
rect 48044 18420 48096 18426
rect 48044 18362 48096 18368
rect 48228 18420 48280 18426
rect 48228 18362 48280 18368
rect 48240 18290 48268 18362
rect 47768 18284 47820 18290
rect 47768 18226 47820 18232
rect 48228 18284 48280 18290
rect 48228 18226 48280 18232
rect 47676 17196 47728 17202
rect 47676 17138 47728 17144
rect 47780 16726 47808 18226
rect 48136 17672 48188 17678
rect 48134 17640 48136 17649
rect 48228 17672 48280 17678
rect 48188 17640 48190 17649
rect 47860 17604 47912 17610
rect 48228 17614 48280 17620
rect 48134 17575 48190 17584
rect 47860 17546 47912 17552
rect 47872 17354 47900 17546
rect 47872 17326 47992 17354
rect 47964 17270 47992 17326
rect 47952 17264 48004 17270
rect 47858 17232 47914 17241
rect 47952 17206 48004 17212
rect 47858 17167 47914 17176
rect 47872 16726 47900 17167
rect 48148 16833 48176 17575
rect 48134 16824 48190 16833
rect 48134 16759 48190 16768
rect 47768 16720 47820 16726
rect 47768 16662 47820 16668
rect 47860 16720 47912 16726
rect 47860 16662 47912 16668
rect 48240 16658 48268 17614
rect 48332 17202 48360 27270
rect 48780 26988 48832 26994
rect 48780 26930 48832 26936
rect 48792 17882 48820 26930
rect 48872 18284 48924 18290
rect 48872 18226 48924 18232
rect 48780 17876 48832 17882
rect 48780 17818 48832 17824
rect 48884 17746 48912 18226
rect 48872 17740 48924 17746
rect 48872 17682 48924 17688
rect 48964 17536 49016 17542
rect 48870 17504 48926 17513
rect 48964 17478 49016 17484
rect 48870 17439 48926 17448
rect 48686 17368 48742 17377
rect 48686 17303 48742 17312
rect 48320 17196 48372 17202
rect 48320 17138 48372 17144
rect 48410 16688 48466 16697
rect 48228 16652 48280 16658
rect 48410 16623 48466 16632
rect 48228 16594 48280 16600
rect 47400 16584 47452 16590
rect 47584 16584 47636 16590
rect 47400 16526 47452 16532
rect 47582 16552 47584 16561
rect 47636 16552 47638 16561
rect 47308 16516 47360 16522
rect 47582 16487 47638 16496
rect 48134 16552 48190 16561
rect 48134 16487 48190 16496
rect 47308 16458 47360 16464
rect 47768 16448 47820 16454
rect 47768 16390 47820 16396
rect 48042 16416 48098 16425
rect 47400 16176 47452 16182
rect 47400 16118 47452 16124
rect 47216 15972 47268 15978
rect 47216 15914 47268 15920
rect 46846 15872 46902 15881
rect 46846 15807 46902 15816
rect 46664 15700 46716 15706
rect 46664 15642 46716 15648
rect 46756 15700 46808 15706
rect 46756 15642 46808 15648
rect 45836 15360 45888 15366
rect 45836 15302 45888 15308
rect 45928 15360 45980 15366
rect 45928 15302 45980 15308
rect 45848 14958 45876 15302
rect 46846 15192 46902 15201
rect 46846 15127 46902 15136
rect 46860 14958 46888 15127
rect 45836 14952 45888 14958
rect 45836 14894 45888 14900
rect 46848 14952 46900 14958
rect 46848 14894 46900 14900
rect 46938 14920 46994 14929
rect 45744 14884 45796 14890
rect 45744 14826 45796 14832
rect 46756 14884 46808 14890
rect 46938 14855 46940 14864
rect 46756 14826 46808 14832
rect 46992 14855 46994 14864
rect 46940 14826 46992 14832
rect 45756 13954 45784 14826
rect 46662 14784 46718 14793
rect 46662 14719 46718 14728
rect 46478 14376 46534 14385
rect 46478 14311 46534 14320
rect 45836 14000 45888 14006
rect 45756 13948 45836 13954
rect 45756 13942 45888 13948
rect 45756 13926 45876 13942
rect 46492 13938 46520 14311
rect 46020 13932 46072 13938
rect 45756 13394 45784 13926
rect 46020 13874 46072 13880
rect 46480 13932 46532 13938
rect 46480 13874 46532 13880
rect 45928 13864 45980 13870
rect 45928 13806 45980 13812
rect 45836 13728 45888 13734
rect 45836 13670 45888 13676
rect 45744 13388 45796 13394
rect 45744 13330 45796 13336
rect 45652 13252 45704 13258
rect 45652 13194 45704 13200
rect 45848 13161 45876 13670
rect 45940 13326 45968 13806
rect 46032 13705 46060 13874
rect 46018 13696 46074 13705
rect 46074 13654 46244 13682
rect 46018 13631 46074 13640
rect 45928 13320 45980 13326
rect 45928 13262 45980 13268
rect 45834 13152 45890 13161
rect 45834 13087 45890 13096
rect 45652 12980 45704 12986
rect 45652 12922 45704 12928
rect 45664 12850 45692 12922
rect 45652 12844 45704 12850
rect 45652 12786 45704 12792
rect 46112 12844 46164 12850
rect 46112 12786 46164 12792
rect 45744 12776 45796 12782
rect 46020 12776 46072 12782
rect 45744 12718 45796 12724
rect 45926 12744 45982 12753
rect 45560 12640 45612 12646
rect 45560 12582 45612 12588
rect 45756 12442 45784 12718
rect 46124 12753 46152 12786
rect 46020 12718 46072 12724
rect 46110 12744 46166 12753
rect 45926 12679 45982 12688
rect 45940 12646 45968 12679
rect 45928 12640 45980 12646
rect 45928 12582 45980 12588
rect 45744 12436 45796 12442
rect 45744 12378 45796 12384
rect 46032 12374 46060 12718
rect 46110 12679 46166 12688
rect 46020 12368 46072 12374
rect 46020 12310 46072 12316
rect 46216 12306 46244 13654
rect 46388 13252 46440 13258
rect 46388 13194 46440 13200
rect 46400 12986 46428 13194
rect 46388 12980 46440 12986
rect 46388 12922 46440 12928
rect 46572 12844 46624 12850
rect 46676 12832 46704 14719
rect 46768 13870 46796 14826
rect 46756 13864 46808 13870
rect 46756 13806 46808 13812
rect 47032 13728 47084 13734
rect 47032 13670 47084 13676
rect 47044 13326 47072 13670
rect 47032 13320 47084 13326
rect 47032 13262 47084 13268
rect 46846 13016 46902 13025
rect 46846 12951 46902 12960
rect 46860 12850 46888 12951
rect 46756 12844 46808 12850
rect 46676 12804 46756 12832
rect 46572 12786 46624 12792
rect 46756 12786 46808 12792
rect 46848 12844 46900 12850
rect 46848 12786 46900 12792
rect 47032 12844 47084 12850
rect 47216 12844 47268 12850
rect 47084 12804 47164 12832
rect 47032 12786 47084 12792
rect 46584 12617 46612 12786
rect 46768 12730 46796 12786
rect 46768 12702 46888 12730
rect 46570 12608 46626 12617
rect 46626 12566 46796 12594
rect 46570 12543 46626 12552
rect 46296 12368 46348 12374
rect 46296 12310 46348 12316
rect 45468 12300 45520 12306
rect 45468 12242 45520 12248
rect 46204 12300 46256 12306
rect 46204 12242 46256 12248
rect 45560 12232 45612 12238
rect 45560 12174 45612 12180
rect 45572 11830 45600 12174
rect 46308 12170 46336 12310
rect 46572 12232 46624 12238
rect 46386 12200 46442 12209
rect 46296 12164 46348 12170
rect 46572 12174 46624 12180
rect 46386 12135 46442 12144
rect 46296 12106 46348 12112
rect 46112 11892 46164 11898
rect 46112 11834 46164 11840
rect 45560 11824 45612 11830
rect 45560 11766 45612 11772
rect 46124 11762 46152 11834
rect 46112 11756 46164 11762
rect 46112 11698 46164 11704
rect 46112 11620 46164 11626
rect 46112 11562 46164 11568
rect 45744 11552 45796 11558
rect 45744 11494 45796 11500
rect 45836 11552 45888 11558
rect 45836 11494 45888 11500
rect 45560 11144 45612 11150
rect 45560 11086 45612 11092
rect 45112 10662 45232 10690
rect 45284 10668 45336 10674
rect 44640 10532 44692 10538
rect 44640 10474 44692 10480
rect 45112 10010 45140 10662
rect 45284 10610 45336 10616
rect 45192 10600 45244 10606
rect 45296 10577 45324 10610
rect 45192 10542 45244 10548
rect 45282 10568 45338 10577
rect 45204 10441 45232 10542
rect 45572 10554 45600 11086
rect 45756 10606 45784 11494
rect 45848 11121 45876 11494
rect 46124 11286 46152 11562
rect 46400 11354 46428 12135
rect 46388 11348 46440 11354
rect 46388 11290 46440 11296
rect 46112 11280 46164 11286
rect 46112 11222 46164 11228
rect 46020 11144 46072 11150
rect 45834 11112 45890 11121
rect 46204 11144 46256 11150
rect 46072 11104 46204 11132
rect 46020 11086 46072 11092
rect 46204 11086 46256 11092
rect 45834 11047 45890 11056
rect 46296 10668 46348 10674
rect 46296 10610 46348 10616
rect 45282 10503 45338 10512
rect 45388 10526 45600 10554
rect 45744 10600 45796 10606
rect 45744 10542 45796 10548
rect 45652 10532 45704 10538
rect 45190 10432 45246 10441
rect 45190 10367 45246 10376
rect 45388 10282 45416 10526
rect 45652 10474 45704 10480
rect 45560 10464 45612 10470
rect 45560 10406 45612 10412
rect 45296 10254 45416 10282
rect 45296 10198 45324 10254
rect 45284 10192 45336 10198
rect 45284 10134 45336 10140
rect 45376 10056 45428 10062
rect 45112 9982 45232 10010
rect 45376 9998 45428 10004
rect 44846 9820 45154 9829
rect 44846 9818 44852 9820
rect 44908 9818 44932 9820
rect 44988 9818 45012 9820
rect 45068 9818 45092 9820
rect 45148 9818 45154 9820
rect 44908 9766 44910 9818
rect 45090 9766 45092 9818
rect 44846 9764 44852 9766
rect 44908 9764 44932 9766
rect 44988 9764 45012 9766
rect 45068 9764 45092 9766
rect 45148 9764 45154 9766
rect 44846 9755 45154 9764
rect 44846 8732 45154 8741
rect 44846 8730 44852 8732
rect 44908 8730 44932 8732
rect 44988 8730 45012 8732
rect 45068 8730 45092 8732
rect 45148 8730 45154 8732
rect 44908 8678 44910 8730
rect 45090 8678 45092 8730
rect 44846 8676 44852 8678
rect 44908 8676 44932 8678
rect 44988 8676 45012 8678
rect 45068 8676 45092 8678
rect 45148 8676 45154 8678
rect 44846 8667 45154 8676
rect 44846 7644 45154 7653
rect 44846 7642 44852 7644
rect 44908 7642 44932 7644
rect 44988 7642 45012 7644
rect 45068 7642 45092 7644
rect 45148 7642 45154 7644
rect 44908 7590 44910 7642
rect 45090 7590 45092 7642
rect 44846 7588 44852 7590
rect 44908 7588 44932 7590
rect 44988 7588 45012 7590
rect 45068 7588 45092 7590
rect 45148 7588 45154 7590
rect 44846 7579 45154 7588
rect 44846 6556 45154 6565
rect 44846 6554 44852 6556
rect 44908 6554 44932 6556
rect 44988 6554 45012 6556
rect 45068 6554 45092 6556
rect 45148 6554 45154 6556
rect 44908 6502 44910 6554
rect 45090 6502 45092 6554
rect 44846 6500 44852 6502
rect 44908 6500 44932 6502
rect 44988 6500 45012 6502
rect 45068 6500 45092 6502
rect 45148 6500 45154 6502
rect 44846 6491 45154 6500
rect 44846 5468 45154 5477
rect 44846 5466 44852 5468
rect 44908 5466 44932 5468
rect 44988 5466 45012 5468
rect 45068 5466 45092 5468
rect 45148 5466 45154 5468
rect 44908 5414 44910 5466
rect 45090 5414 45092 5466
rect 44846 5412 44852 5414
rect 44908 5412 44932 5414
rect 44988 5412 45012 5414
rect 45068 5412 45092 5414
rect 45148 5412 45154 5414
rect 44846 5403 45154 5412
rect 44548 5228 44600 5234
rect 44548 5170 44600 5176
rect 44846 4380 45154 4389
rect 44846 4378 44852 4380
rect 44908 4378 44932 4380
rect 44988 4378 45012 4380
rect 45068 4378 45092 4380
rect 45148 4378 45154 4380
rect 44908 4326 44910 4378
rect 45090 4326 45092 4378
rect 44846 4324 44852 4326
rect 44908 4324 44932 4326
rect 44988 4324 45012 4326
rect 45068 4324 45092 4326
rect 45148 4324 45154 4326
rect 44846 4315 45154 4324
rect 44364 4140 44416 4146
rect 44364 4082 44416 4088
rect 45204 3398 45232 9982
rect 45388 9874 45416 9998
rect 45572 9994 45600 10406
rect 45664 9994 45692 10474
rect 45560 9988 45612 9994
rect 45560 9930 45612 9936
rect 45652 9988 45704 9994
rect 45652 9930 45704 9936
rect 45756 9874 45784 10542
rect 45388 9846 45784 9874
rect 45572 9518 45600 9846
rect 45836 9580 45888 9586
rect 45836 9522 45888 9528
rect 45560 9512 45612 9518
rect 45560 9454 45612 9460
rect 45848 9178 45876 9522
rect 45836 9172 45888 9178
rect 45836 9114 45888 9120
rect 46112 8968 46164 8974
rect 46112 8910 46164 8916
rect 46124 8634 46152 8910
rect 46112 8628 46164 8634
rect 46112 8570 46164 8576
rect 45744 8424 45796 8430
rect 45744 8366 45796 8372
rect 45376 4072 45428 4078
rect 45376 4014 45428 4020
rect 45388 3602 45416 4014
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45192 3392 45244 3398
rect 45192 3334 45244 3340
rect 44846 3292 45154 3301
rect 44846 3290 44852 3292
rect 44908 3290 44932 3292
rect 44988 3290 45012 3292
rect 45068 3290 45092 3292
rect 45148 3290 45154 3292
rect 44908 3238 44910 3290
rect 45090 3238 45092 3290
rect 44846 3236 44852 3238
rect 44908 3236 44932 3238
rect 44988 3236 45012 3238
rect 45068 3236 45092 3238
rect 45148 3236 45154 3238
rect 44846 3227 45154 3236
rect 43904 3052 43956 3058
rect 43904 2994 43956 3000
rect 45282 2952 45338 2961
rect 45282 2887 45338 2896
rect 45466 2952 45522 2961
rect 45466 2887 45522 2896
rect 45296 2582 45324 2887
rect 45480 2650 45508 2887
rect 45558 2816 45614 2825
rect 45558 2751 45614 2760
rect 45468 2644 45520 2650
rect 45468 2586 45520 2592
rect 43720 2576 43772 2582
rect 43720 2518 43772 2524
rect 45284 2576 45336 2582
rect 45284 2518 45336 2524
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 42800 2440 42852 2446
rect 42800 2382 42852 2388
rect 43444 2440 43496 2446
rect 43444 2382 43496 2388
rect 44456 2440 44508 2446
rect 44456 2382 44508 2388
rect 45192 2440 45244 2446
rect 45192 2382 45244 2388
rect 41696 2372 41748 2378
rect 41696 2314 41748 2320
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 42524 2304 42576 2310
rect 42524 2246 42576 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 41892 800 41920 2246
rect 42536 800 42564 2246
rect 43180 800 43208 2246
rect 43824 800 43852 2246
rect 44468 800 44496 2382
rect 44846 2204 45154 2213
rect 44846 2202 44852 2204
rect 44908 2202 44932 2204
rect 44988 2202 45012 2204
rect 45068 2202 45092 2204
rect 45148 2202 45154 2204
rect 44908 2150 44910 2202
rect 45090 2150 45092 2202
rect 44846 2148 44852 2150
rect 44908 2148 44932 2150
rect 44988 2148 45012 2150
rect 45068 2148 45092 2150
rect 45148 2148 45154 2150
rect 44846 2139 45154 2148
rect 45204 1306 45232 2382
rect 45572 2310 45600 2751
rect 45560 2304 45612 2310
rect 45560 2246 45612 2252
rect 45560 2032 45612 2038
rect 45558 2000 45560 2009
rect 45652 2032 45704 2038
rect 45612 2000 45614 2009
rect 45652 1974 45704 1980
rect 45558 1935 45614 1944
rect 45558 1728 45614 1737
rect 45558 1663 45560 1672
rect 45612 1663 45614 1672
rect 45560 1634 45612 1640
rect 45376 1624 45428 1630
rect 45376 1566 45428 1572
rect 45388 1358 45416 1566
rect 45664 1442 45692 1974
rect 45572 1426 45692 1442
rect 45756 1426 45784 8366
rect 46308 4486 46336 10610
rect 46388 9376 46440 9382
rect 46388 9318 46440 9324
rect 46400 8974 46428 9318
rect 46388 8968 46440 8974
rect 46388 8910 46440 8916
rect 46296 4480 46348 4486
rect 46296 4422 46348 4428
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3738 46336 3878
rect 46296 3732 46348 3738
rect 46296 3674 46348 3680
rect 46020 3528 46072 3534
rect 46020 3470 46072 3476
rect 46032 3194 46060 3470
rect 46020 3188 46072 3194
rect 46020 3130 46072 3136
rect 46400 2990 46428 8910
rect 46480 8900 46532 8906
rect 46480 8842 46532 8848
rect 46492 8090 46520 8842
rect 46480 8084 46532 8090
rect 46480 8026 46532 8032
rect 46478 4040 46534 4049
rect 46478 3975 46480 3984
rect 46532 3975 46534 3984
rect 46480 3946 46532 3952
rect 46296 2984 46348 2990
rect 46296 2926 46348 2932
rect 46388 2984 46440 2990
rect 46388 2926 46440 2932
rect 46308 2650 46336 2926
rect 46584 2825 46612 12174
rect 46768 12073 46796 12566
rect 46860 12306 46888 12702
rect 47136 12617 47164 12804
rect 47216 12786 47268 12792
rect 47122 12608 47178 12617
rect 47122 12543 47178 12552
rect 46848 12300 46900 12306
rect 46848 12242 46900 12248
rect 46754 12064 46810 12073
rect 46754 11999 46810 12008
rect 46754 11928 46810 11937
rect 46754 11863 46810 11872
rect 46768 11762 46796 11863
rect 46756 11756 46808 11762
rect 46756 11698 46808 11704
rect 47136 11393 47164 12543
rect 47228 11762 47256 12786
rect 47308 12300 47360 12306
rect 47308 12242 47360 12248
rect 47216 11756 47268 11762
rect 47216 11698 47268 11704
rect 47320 11393 47348 12242
rect 47122 11384 47178 11393
rect 47122 11319 47178 11328
rect 47306 11384 47362 11393
rect 47306 11319 47362 11328
rect 46664 11144 46716 11150
rect 46664 11086 46716 11092
rect 46756 11144 46808 11150
rect 46756 11086 46808 11092
rect 47216 11144 47268 11150
rect 47216 11086 47268 11092
rect 46676 10198 46704 11086
rect 46768 10577 46796 11086
rect 47124 10668 47176 10674
rect 47124 10610 47176 10616
rect 46754 10568 46810 10577
rect 46754 10503 46810 10512
rect 46768 10470 46796 10503
rect 46756 10464 46808 10470
rect 46756 10406 46808 10412
rect 46664 10192 46716 10198
rect 46664 10134 46716 10140
rect 46768 9994 46796 10406
rect 47136 10266 47164 10610
rect 47228 10470 47256 11086
rect 47216 10464 47268 10470
rect 47214 10432 47216 10441
rect 47268 10432 47270 10441
rect 47214 10367 47270 10376
rect 47124 10260 47176 10266
rect 47124 10202 47176 10208
rect 46756 9988 46808 9994
rect 46756 9930 46808 9936
rect 47228 9926 47256 10367
rect 47216 9920 47268 9926
rect 47216 9862 47268 9868
rect 47412 9654 47440 16118
rect 47780 16114 47808 16390
rect 48042 16351 48098 16360
rect 47768 16108 47820 16114
rect 47768 16050 47820 16056
rect 48056 16046 48084 16351
rect 47492 16040 47544 16046
rect 47492 15982 47544 15988
rect 47676 16040 47728 16046
rect 47676 15982 47728 15988
rect 48044 16040 48096 16046
rect 48044 15982 48096 15988
rect 47504 15570 47532 15982
rect 47688 15892 47716 15982
rect 48148 15978 48176 16487
rect 48228 16448 48280 16454
rect 48228 16390 48280 16396
rect 48240 16289 48268 16390
rect 48226 16280 48282 16289
rect 48226 16215 48282 16224
rect 48240 16114 48268 16215
rect 48424 16114 48452 16623
rect 48228 16108 48280 16114
rect 48228 16050 48280 16056
rect 48412 16108 48464 16114
rect 48596 16108 48648 16114
rect 48464 16068 48596 16096
rect 48412 16050 48464 16056
rect 48596 16050 48648 16056
rect 48136 15972 48188 15978
rect 48136 15914 48188 15920
rect 47768 15904 47820 15910
rect 47688 15864 47768 15892
rect 47768 15846 47820 15852
rect 48226 15736 48282 15745
rect 48226 15671 48228 15680
rect 48280 15671 48282 15680
rect 48502 15736 48558 15745
rect 48502 15671 48558 15680
rect 48228 15642 48280 15648
rect 48042 15600 48098 15609
rect 47492 15564 47544 15570
rect 48042 15535 48098 15544
rect 47492 15506 47544 15512
rect 47676 15496 47728 15502
rect 47676 15438 47728 15444
rect 47688 14521 47716 15438
rect 48056 15366 48084 15535
rect 48516 15484 48544 15671
rect 48700 15502 48728 17303
rect 48780 17196 48832 17202
rect 48780 17138 48832 17144
rect 48424 15456 48544 15484
rect 48688 15496 48740 15502
rect 48424 15450 48452 15456
rect 48286 15434 48452 15450
rect 48688 15438 48740 15444
rect 48274 15428 48452 15434
rect 48326 15422 48452 15428
rect 48274 15370 48326 15376
rect 48044 15360 48096 15366
rect 48792 15337 48820 17138
rect 48044 15302 48096 15308
rect 48318 15328 48374 15337
rect 48318 15263 48374 15272
rect 48778 15328 48834 15337
rect 48778 15263 48834 15272
rect 48332 15026 48360 15263
rect 48884 15042 48912 17439
rect 48976 17066 49004 17478
rect 48964 17060 49016 17066
rect 48964 17002 49016 17008
rect 48320 15020 48372 15026
rect 48320 14962 48372 14968
rect 48596 15020 48648 15026
rect 48596 14962 48648 14968
rect 48700 15014 48912 15042
rect 48608 14822 48636 14962
rect 48596 14816 48648 14822
rect 48410 14784 48466 14793
rect 48596 14758 48648 14764
rect 48410 14719 48466 14728
rect 47674 14512 47730 14521
rect 47674 14447 47730 14456
rect 47768 14408 47820 14414
rect 47768 14350 47820 14356
rect 47492 14272 47544 14278
rect 47490 14240 47492 14249
rect 47676 14272 47728 14278
rect 47544 14240 47546 14249
rect 47676 14214 47728 14220
rect 47490 14175 47546 14184
rect 47688 13394 47716 14214
rect 47780 14006 47808 14350
rect 48424 14278 48452 14719
rect 48608 14414 48636 14758
rect 48596 14408 48648 14414
rect 48596 14350 48648 14356
rect 48412 14272 48464 14278
rect 48412 14214 48464 14220
rect 48504 14272 48556 14278
rect 48504 14214 48556 14220
rect 47768 14000 47820 14006
rect 47768 13942 47820 13948
rect 47780 13462 47808 13942
rect 48044 13932 48096 13938
rect 48044 13874 48096 13880
rect 47858 13832 47914 13841
rect 47858 13767 47914 13776
rect 47872 13462 47900 13767
rect 47952 13728 48004 13734
rect 47952 13670 48004 13676
rect 47768 13456 47820 13462
rect 47768 13398 47820 13404
rect 47860 13456 47912 13462
rect 47860 13398 47912 13404
rect 47676 13388 47728 13394
rect 47676 13330 47728 13336
rect 47688 12918 47716 13330
rect 47964 13326 47992 13670
rect 47952 13320 48004 13326
rect 47952 13262 48004 13268
rect 47768 13184 47820 13190
rect 48056 13172 48084 13874
rect 48318 13832 48374 13841
rect 48318 13767 48374 13776
rect 48226 13560 48282 13569
rect 48226 13495 48282 13504
rect 48136 13320 48188 13326
rect 48136 13262 48188 13268
rect 47768 13126 47820 13132
rect 47872 13144 48084 13172
rect 47780 12918 47808 13126
rect 47676 12912 47728 12918
rect 47676 12854 47728 12860
rect 47768 12912 47820 12918
rect 47768 12854 47820 12860
rect 47584 12232 47636 12238
rect 47584 12174 47636 12180
rect 47596 11898 47624 12174
rect 47768 12164 47820 12170
rect 47768 12106 47820 12112
rect 47676 12096 47728 12102
rect 47676 12038 47728 12044
rect 47688 11898 47716 12038
rect 47584 11892 47636 11898
rect 47584 11834 47636 11840
rect 47676 11892 47728 11898
rect 47676 11834 47728 11840
rect 47780 11812 47808 12106
rect 47872 12102 47900 13144
rect 48044 12776 48096 12782
rect 48044 12718 48096 12724
rect 48056 12646 48084 12718
rect 48148 12646 48176 13262
rect 48044 12640 48096 12646
rect 48044 12582 48096 12588
rect 48136 12640 48188 12646
rect 48136 12582 48188 12588
rect 48134 12472 48190 12481
rect 48240 12442 48268 13495
rect 48332 13258 48360 13767
rect 48320 13252 48372 13258
rect 48320 13194 48372 13200
rect 48320 12980 48372 12986
rect 48320 12922 48372 12928
rect 48332 12730 48360 12922
rect 48424 12889 48452 14214
rect 48410 12880 48466 12889
rect 48410 12815 48466 12824
rect 48332 12702 48452 12730
rect 48424 12594 48452 12702
rect 48332 12566 48452 12594
rect 48134 12407 48190 12416
rect 48228 12436 48280 12442
rect 48044 12368 48096 12374
rect 48044 12310 48096 12316
rect 47860 12096 47912 12102
rect 48056 12073 48084 12310
rect 47860 12038 47912 12044
rect 48042 12064 48098 12073
rect 48042 11999 48098 12008
rect 48148 11898 48176 12407
rect 48228 12378 48280 12384
rect 48332 12238 48360 12566
rect 48410 12472 48466 12481
rect 48410 12407 48466 12416
rect 48320 12232 48372 12238
rect 48320 12174 48372 12180
rect 48228 12164 48280 12170
rect 48228 12106 48280 12112
rect 48136 11892 48188 11898
rect 48136 11834 48188 11840
rect 48240 11830 48268 12106
rect 48424 12073 48452 12407
rect 48410 12064 48466 12073
rect 48410 11999 48466 12008
rect 47860 11824 47912 11830
rect 47780 11784 47860 11812
rect 47860 11766 47912 11772
rect 48228 11824 48280 11830
rect 48228 11766 48280 11772
rect 47584 11552 47636 11558
rect 48516 11529 48544 14214
rect 48596 14000 48648 14006
rect 48596 13942 48648 13948
rect 48608 12238 48636 13942
rect 48700 13462 48728 15014
rect 48872 14952 48924 14958
rect 48870 14920 48872 14929
rect 48924 14920 48926 14929
rect 48870 14855 48926 14864
rect 49068 14278 49096 27406
rect 49620 26976 49648 29200
rect 50540 27470 50568 29294
rect 50894 29294 51028 29322
rect 50894 29200 50950 29294
rect 51000 27588 51028 29294
rect 51538 29294 51856 29322
rect 51538 29200 51594 29294
rect 51080 27600 51132 27606
rect 51000 27560 51080 27588
rect 51080 27542 51132 27548
rect 51264 27600 51316 27606
rect 51264 27542 51316 27548
rect 50528 27464 50580 27470
rect 50528 27406 50580 27412
rect 51172 27396 51224 27402
rect 51276 27384 51304 27542
rect 51828 27470 51856 29294
rect 52182 29294 52408 29322
rect 52182 29200 52238 29294
rect 52276 27668 52328 27674
rect 52276 27610 52328 27616
rect 51816 27464 51868 27470
rect 51816 27406 51868 27412
rect 51224 27356 51304 27384
rect 51724 27396 51776 27402
rect 51172 27338 51224 27344
rect 51724 27338 51776 27344
rect 50436 27328 50488 27334
rect 50436 27270 50488 27276
rect 49700 26988 49752 26994
rect 49620 26948 49700 26976
rect 49700 26930 49752 26936
rect 49332 26784 49384 26790
rect 49332 26726 49384 26732
rect 50344 26784 50396 26790
rect 50344 26726 50396 26732
rect 49344 18426 49372 26726
rect 50160 18692 50212 18698
rect 50160 18634 50212 18640
rect 49148 18420 49200 18426
rect 49148 18362 49200 18368
rect 49332 18420 49384 18426
rect 49332 18362 49384 18368
rect 49160 17678 49188 18362
rect 49344 18290 49372 18362
rect 49332 18284 49384 18290
rect 49332 18226 49384 18232
rect 49608 18148 49660 18154
rect 49608 18090 49660 18096
rect 49148 17672 49200 17678
rect 49148 17614 49200 17620
rect 49240 17672 49292 17678
rect 49240 17614 49292 17620
rect 49160 17542 49188 17614
rect 49148 17536 49200 17542
rect 49148 17478 49200 17484
rect 49148 14408 49200 14414
rect 49148 14350 49200 14356
rect 49056 14272 49108 14278
rect 49056 14214 49108 14220
rect 48780 14000 48832 14006
rect 48780 13942 48832 13948
rect 48688 13456 48740 13462
rect 48688 13398 48740 13404
rect 48688 13320 48740 13326
rect 48688 13262 48740 13268
rect 48700 13190 48728 13262
rect 48688 13184 48740 13190
rect 48688 13126 48740 13132
rect 48700 12481 48728 13126
rect 48686 12472 48742 12481
rect 48686 12407 48742 12416
rect 48596 12232 48648 12238
rect 48596 12174 48648 12180
rect 48608 11898 48636 12174
rect 48596 11892 48648 11898
rect 48596 11834 48648 11840
rect 47584 11494 47636 11500
rect 48502 11520 48558 11529
rect 47596 11286 47624 11494
rect 48502 11455 48558 11464
rect 47584 11280 47636 11286
rect 47584 11222 47636 11228
rect 48044 10464 48096 10470
rect 48044 10406 48096 10412
rect 47858 10160 47914 10169
rect 47858 10095 47914 10104
rect 47492 9920 47544 9926
rect 47492 9862 47544 9868
rect 47400 9648 47452 9654
rect 47400 9590 47452 9596
rect 47504 9450 47532 9862
rect 47492 9444 47544 9450
rect 47492 9386 47544 9392
rect 46940 8900 46992 8906
rect 46940 8842 46992 8848
rect 46570 2816 46626 2825
rect 46570 2751 46626 2760
rect 46296 2644 46348 2650
rect 46296 2586 46348 2592
rect 46848 2508 46900 2514
rect 46952 2496 46980 8842
rect 47504 8634 47532 9386
rect 47492 8628 47544 8634
rect 47492 8570 47544 8576
rect 47872 3738 47900 10095
rect 47860 3732 47912 3738
rect 47860 3674 47912 3680
rect 47492 3596 47544 3602
rect 47492 3538 47544 3544
rect 47504 3398 47532 3538
rect 47124 3392 47176 3398
rect 47124 3334 47176 3340
rect 47492 3392 47544 3398
rect 47492 3334 47544 3340
rect 47136 3058 47164 3334
rect 47124 3052 47176 3058
rect 47124 2994 47176 3000
rect 47504 2854 47532 3334
rect 47492 2848 47544 2854
rect 47492 2790 47544 2796
rect 48056 2530 48084 10406
rect 48136 9172 48188 9178
rect 48136 9114 48188 9120
rect 48412 9172 48464 9178
rect 48412 9114 48464 9120
rect 48148 7886 48176 9114
rect 48424 8974 48452 9114
rect 48412 8968 48464 8974
rect 48412 8910 48464 8916
rect 48424 8634 48452 8910
rect 48412 8628 48464 8634
rect 48412 8570 48464 8576
rect 48136 7880 48188 7886
rect 48136 7822 48188 7828
rect 48516 6458 48544 11455
rect 48688 10668 48740 10674
rect 48688 10610 48740 10616
rect 48596 9376 48648 9382
rect 48596 9318 48648 9324
rect 48608 9042 48636 9318
rect 48596 9036 48648 9042
rect 48596 8978 48648 8984
rect 48608 8498 48636 8978
rect 48596 8492 48648 8498
rect 48596 8434 48648 8440
rect 48504 6452 48556 6458
rect 48504 6394 48556 6400
rect 48226 3768 48282 3777
rect 48226 3703 48282 3712
rect 48240 3670 48268 3703
rect 48228 3664 48280 3670
rect 48228 3606 48280 3612
rect 48136 3596 48188 3602
rect 48136 3538 48188 3544
rect 48148 3505 48176 3538
rect 48134 3496 48190 3505
rect 48700 3466 48728 10610
rect 48134 3431 48190 3440
rect 48688 3460 48740 3466
rect 48688 3402 48740 3408
rect 48792 2774 48820 13942
rect 48964 13932 49016 13938
rect 48964 13874 49016 13880
rect 48870 13560 48926 13569
rect 48870 13495 48926 13504
rect 48884 13394 48912 13495
rect 48872 13388 48924 13394
rect 48872 13330 48924 13336
rect 48872 12640 48924 12646
rect 48872 12582 48924 12588
rect 48884 12073 48912 12582
rect 48976 12306 49004 13874
rect 49056 13796 49108 13802
rect 49056 13738 49108 13744
rect 49068 13394 49096 13738
rect 49056 13388 49108 13394
rect 49056 13330 49108 13336
rect 49160 12850 49188 14350
rect 49252 14006 49280 17614
rect 49422 17232 49478 17241
rect 49422 17167 49478 17176
rect 49436 17134 49464 17167
rect 49424 17128 49476 17134
rect 49424 17070 49476 17076
rect 49620 17066 49648 18090
rect 50172 17882 50200 18634
rect 50160 17876 50212 17882
rect 50160 17818 50212 17824
rect 49698 17368 49754 17377
rect 49698 17303 49754 17312
rect 50066 17368 50122 17377
rect 50066 17303 50122 17312
rect 49712 17202 49740 17303
rect 49700 17196 49752 17202
rect 49700 17138 49752 17144
rect 49884 17196 49936 17202
rect 49884 17138 49936 17144
rect 49608 17060 49660 17066
rect 49608 17002 49660 17008
rect 49792 16652 49844 16658
rect 49792 16594 49844 16600
rect 49606 16280 49662 16289
rect 49606 16215 49662 16224
rect 49620 16046 49648 16215
rect 49608 16040 49660 16046
rect 49608 15982 49660 15988
rect 49700 16040 49752 16046
rect 49700 15982 49752 15988
rect 49422 15872 49478 15881
rect 49422 15807 49478 15816
rect 49436 15638 49464 15807
rect 49332 15632 49384 15638
rect 49332 15574 49384 15580
rect 49424 15632 49476 15638
rect 49424 15574 49476 15580
rect 49240 14000 49292 14006
rect 49240 13942 49292 13948
rect 49252 13705 49280 13942
rect 49238 13696 49294 13705
rect 49238 13631 49294 13640
rect 49238 13560 49294 13569
rect 49238 13495 49294 13504
rect 49252 13326 49280 13495
rect 49240 13320 49292 13326
rect 49240 13262 49292 13268
rect 49148 12844 49200 12850
rect 49148 12786 49200 12792
rect 48964 12300 49016 12306
rect 48964 12242 49016 12248
rect 48870 12064 48926 12073
rect 48870 11999 48926 12008
rect 49238 11520 49294 11529
rect 49238 11455 49294 11464
rect 49252 11218 49280 11455
rect 49240 11212 49292 11218
rect 49240 11154 49292 11160
rect 48964 10056 49016 10062
rect 48964 9998 49016 10004
rect 48976 8974 49004 9998
rect 48964 8968 49016 8974
rect 48964 8910 49016 8916
rect 49240 4480 49292 4486
rect 49240 4422 49292 4428
rect 49252 4214 49280 4422
rect 49240 4208 49292 4214
rect 49240 4150 49292 4156
rect 48872 3528 48924 3534
rect 48870 3496 48872 3505
rect 48964 3528 49016 3534
rect 48924 3496 48926 3505
rect 48964 3470 49016 3476
rect 48870 3431 48926 3440
rect 46900 2468 46980 2496
rect 47872 2502 48084 2530
rect 48516 2746 48820 2774
rect 46848 2450 46900 2456
rect 46388 2440 46440 2446
rect 46388 2382 46440 2388
rect 46756 2440 46808 2446
rect 46756 2382 46808 2388
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 45834 1864 45890 1873
rect 45834 1799 45890 1808
rect 45848 1698 45876 1799
rect 45836 1692 45888 1698
rect 45836 1634 45888 1640
rect 45560 1420 45692 1426
rect 45612 1414 45692 1420
rect 45744 1420 45796 1426
rect 45560 1362 45612 1368
rect 45744 1362 45796 1368
rect 45112 1278 45232 1306
rect 45376 1352 45428 1358
rect 45376 1294 45428 1300
rect 45112 800 45140 1278
rect 46400 800 46428 2382
rect 46768 1358 46796 2382
rect 46756 1352 46808 1358
rect 46756 1294 46808 1300
rect 47044 800 47072 2382
rect 47872 2378 47900 2502
rect 48228 2440 48280 2446
rect 47964 2400 48228 2428
rect 47860 2372 47912 2378
rect 47860 2314 47912 2320
rect 47124 1624 47176 1630
rect 47124 1566 47176 1572
rect 47136 1426 47164 1566
rect 47124 1420 47176 1426
rect 47124 1362 47176 1368
rect 47688 870 47808 898
rect 47688 800 47716 870
rect 31312 734 31524 762
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 47780 762 47808 870
rect 47964 762 47992 2400
rect 48412 2440 48464 2446
rect 48228 2382 48280 2388
rect 48332 2400 48412 2428
rect 48044 2304 48096 2310
rect 48228 2304 48280 2310
rect 48096 2264 48228 2292
rect 48044 2246 48096 2252
rect 48228 2246 48280 2252
rect 48332 800 48360 2400
rect 48412 2382 48464 2388
rect 48516 1737 48544 2746
rect 48780 2304 48832 2310
rect 48780 2246 48832 2252
rect 48792 2038 48820 2246
rect 48780 2032 48832 2038
rect 48872 2032 48924 2038
rect 48780 1974 48832 1980
rect 48870 2000 48872 2009
rect 48924 2000 48926 2009
rect 48870 1935 48926 1944
rect 48502 1728 48558 1737
rect 48502 1663 48558 1672
rect 48976 800 49004 3470
rect 49240 3392 49292 3398
rect 49240 3334 49292 3340
rect 49252 3233 49280 3334
rect 49238 3224 49294 3233
rect 49238 3159 49294 3168
rect 49344 2774 49372 15574
rect 49712 15366 49740 15982
rect 49700 15360 49752 15366
rect 49700 15302 49752 15308
rect 49804 14822 49832 16594
rect 49896 16046 49924 17138
rect 49974 17096 50030 17105
rect 49974 17031 49976 17040
rect 50028 17031 50030 17040
rect 49976 17002 50028 17008
rect 50080 16726 50108 17303
rect 50160 17128 50212 17134
rect 50160 17070 50212 17076
rect 50068 16720 50120 16726
rect 50068 16662 50120 16668
rect 50172 16114 50200 17070
rect 50250 16824 50306 16833
rect 50250 16759 50306 16768
rect 50264 16590 50292 16759
rect 50252 16584 50304 16590
rect 50252 16526 50304 16532
rect 50356 16454 50384 26726
rect 50252 16448 50304 16454
rect 50252 16390 50304 16396
rect 50344 16448 50396 16454
rect 50344 16390 50396 16396
rect 49976 16108 50028 16114
rect 49976 16050 50028 16056
rect 50160 16108 50212 16114
rect 50160 16050 50212 16056
rect 49884 16040 49936 16046
rect 49884 15982 49936 15988
rect 49884 15904 49936 15910
rect 49884 15846 49936 15852
rect 49792 14816 49844 14822
rect 49792 14758 49844 14764
rect 49516 14272 49568 14278
rect 49516 14214 49568 14220
rect 49528 13802 49556 14214
rect 49804 13870 49832 14758
rect 49792 13864 49844 13870
rect 49792 13806 49844 13812
rect 49516 13796 49568 13802
rect 49516 13738 49568 13744
rect 49804 13462 49832 13806
rect 49792 13456 49844 13462
rect 49792 13398 49844 13404
rect 49424 13320 49476 13326
rect 49424 13262 49476 13268
rect 49516 13320 49568 13326
rect 49516 13262 49568 13268
rect 49436 13161 49464 13262
rect 49422 13152 49478 13161
rect 49422 13087 49478 13096
rect 49528 13025 49556 13262
rect 49606 13152 49662 13161
rect 49606 13087 49662 13096
rect 49514 13016 49570 13025
rect 49514 12951 49570 12960
rect 49620 12850 49648 13087
rect 49608 12844 49660 12850
rect 49608 12786 49660 12792
rect 49896 12764 49924 15846
rect 49988 15609 50016 16050
rect 50160 15972 50212 15978
rect 50160 15914 50212 15920
rect 50172 15881 50200 15914
rect 50158 15872 50214 15881
rect 50158 15807 50214 15816
rect 49974 15600 50030 15609
rect 49974 15535 50030 15544
rect 49988 15366 50016 15535
rect 50172 15434 50200 15807
rect 50264 15706 50292 16390
rect 50356 16114 50384 16390
rect 50344 16108 50396 16114
rect 50344 16050 50396 16056
rect 50252 15700 50304 15706
rect 50252 15642 50304 15648
rect 50252 15496 50304 15502
rect 50448 15450 50476 27270
rect 50804 27124 50856 27130
rect 50804 27066 50856 27072
rect 50526 18184 50582 18193
rect 50526 18119 50582 18128
rect 50540 17678 50568 18119
rect 50528 17672 50580 17678
rect 50528 17614 50580 17620
rect 50816 17202 50844 27066
rect 51172 18216 51224 18222
rect 51172 18158 51224 18164
rect 51080 18148 51132 18154
rect 51080 18090 51132 18096
rect 51092 17882 51120 18090
rect 51080 17876 51132 17882
rect 51080 17818 51132 17824
rect 50528 17196 50580 17202
rect 50528 17138 50580 17144
rect 50804 17196 50856 17202
rect 50804 17138 50856 17144
rect 50540 16046 50568 17138
rect 50816 16998 50844 17138
rect 51080 17128 51132 17134
rect 51184 17082 51212 18158
rect 51132 17076 51304 17082
rect 51080 17070 51304 17076
rect 51092 17054 51304 17070
rect 50804 16992 50856 16998
rect 50724 16952 50804 16980
rect 50618 16688 50674 16697
rect 50618 16623 50674 16632
rect 50632 16114 50660 16623
rect 50620 16108 50672 16114
rect 50620 16050 50672 16056
rect 50528 16040 50580 16046
rect 50528 15982 50580 15988
rect 50252 15438 50304 15444
rect 50160 15428 50212 15434
rect 50160 15370 50212 15376
rect 49976 15360 50028 15366
rect 49976 15302 50028 15308
rect 50264 14006 50292 15438
rect 50356 15422 50476 15450
rect 50356 14113 50384 15422
rect 50436 15360 50488 15366
rect 50436 15302 50488 15308
rect 50448 15094 50476 15302
rect 50436 15088 50488 15094
rect 50436 15030 50488 15036
rect 50434 14376 50490 14385
rect 50434 14311 50436 14320
rect 50488 14311 50490 14320
rect 50436 14282 50488 14288
rect 50342 14104 50398 14113
rect 50540 14090 50568 15982
rect 50724 15910 50752 16952
rect 50988 16992 51040 16998
rect 50804 16934 50856 16940
rect 50986 16960 50988 16969
rect 51040 16960 51042 16969
rect 50986 16895 51042 16904
rect 51276 16726 51304 17054
rect 51356 16992 51408 16998
rect 51356 16934 51408 16940
rect 51264 16720 51316 16726
rect 51264 16662 51316 16668
rect 51172 16652 51224 16658
rect 51092 16612 51172 16640
rect 51092 16522 51120 16612
rect 51172 16594 51224 16600
rect 51368 16590 51396 16934
rect 51356 16584 51408 16590
rect 51356 16526 51408 16532
rect 50896 16516 50948 16522
rect 50896 16458 50948 16464
rect 50988 16516 51040 16522
rect 50988 16458 51040 16464
rect 51080 16516 51132 16522
rect 51080 16458 51132 16464
rect 50908 16182 50936 16458
rect 50804 16176 50856 16182
rect 50804 16118 50856 16124
rect 50896 16176 50948 16182
rect 50896 16118 50948 16124
rect 50712 15904 50764 15910
rect 50712 15846 50764 15852
rect 50816 15434 50844 16118
rect 50804 15428 50856 15434
rect 50804 15370 50856 15376
rect 51000 15201 51028 16458
rect 51448 16448 51500 16454
rect 51354 16416 51410 16425
rect 51632 16448 51684 16454
rect 51500 16396 51632 16402
rect 51448 16390 51684 16396
rect 51460 16374 51672 16390
rect 51354 16351 51410 16360
rect 51368 16250 51396 16351
rect 51356 16244 51408 16250
rect 51356 16186 51408 16192
rect 51172 16176 51224 16182
rect 51172 16118 51224 16124
rect 51184 16017 51212 16118
rect 51540 16108 51592 16114
rect 51540 16050 51592 16056
rect 51170 16008 51226 16017
rect 51170 15943 51226 15952
rect 51448 15700 51500 15706
rect 51448 15642 51500 15648
rect 51460 15502 51488 15642
rect 51080 15496 51132 15502
rect 51264 15496 51316 15502
rect 51132 15456 51212 15484
rect 51080 15438 51132 15444
rect 51078 15328 51134 15337
rect 51078 15263 51134 15272
rect 50986 15192 51042 15201
rect 50986 15127 51042 15136
rect 51092 15094 51120 15263
rect 51080 15088 51132 15094
rect 51080 15030 51132 15036
rect 50988 14884 51040 14890
rect 50988 14826 51040 14832
rect 50618 14648 50674 14657
rect 50618 14583 50674 14592
rect 50894 14648 50950 14657
rect 50894 14583 50896 14592
rect 50632 14362 50660 14583
rect 50948 14583 50950 14592
rect 50896 14554 50948 14560
rect 51000 14550 51028 14826
rect 51080 14816 51132 14822
rect 51080 14758 51132 14764
rect 50988 14544 51040 14550
rect 50988 14486 51040 14492
rect 50896 14408 50948 14414
rect 50632 14334 50752 14362
rect 50896 14350 50948 14356
rect 50620 14272 50672 14278
rect 50618 14240 50620 14249
rect 50672 14240 50674 14249
rect 50724 14226 50752 14334
rect 50802 14240 50858 14249
rect 50724 14198 50802 14226
rect 50618 14175 50674 14184
rect 50802 14175 50858 14184
rect 50908 14090 50936 14350
rect 50540 14062 50752 14090
rect 50342 14039 50398 14048
rect 50160 14000 50212 14006
rect 50160 13942 50212 13948
rect 50252 14000 50304 14006
rect 50252 13942 50304 13948
rect 50172 13734 50200 13942
rect 50160 13728 50212 13734
rect 50160 13670 50212 13676
rect 50158 13560 50214 13569
rect 50158 13495 50214 13504
rect 50172 13394 50200 13495
rect 50160 13388 50212 13394
rect 50160 13330 50212 13336
rect 50172 12782 50200 12813
rect 49804 12736 49924 12764
rect 50160 12776 50212 12782
rect 50158 12744 50160 12753
rect 50212 12744 50214 12753
rect 49700 12232 49752 12238
rect 49700 12174 49752 12180
rect 49424 12164 49476 12170
rect 49424 12106 49476 12112
rect 49436 11150 49464 12106
rect 49608 11892 49660 11898
rect 49608 11834 49660 11840
rect 49516 11688 49568 11694
rect 49516 11630 49568 11636
rect 49424 11144 49476 11150
rect 49424 11086 49476 11092
rect 49528 10849 49556 11630
rect 49620 11121 49648 11834
rect 49606 11112 49662 11121
rect 49606 11047 49662 11056
rect 49514 10840 49570 10849
rect 49514 10775 49570 10784
rect 49712 10266 49740 12174
rect 49804 11506 49832 12736
rect 50158 12679 50214 12688
rect 49974 12336 50030 12345
rect 49974 12271 50030 12280
rect 49988 12238 50016 12271
rect 49976 12232 50028 12238
rect 49976 12174 50028 12180
rect 49884 11892 49936 11898
rect 49884 11834 49936 11840
rect 49896 11626 49924 11834
rect 50172 11778 50200 12679
rect 50264 12238 50292 13942
rect 50436 13728 50488 13734
rect 50436 13670 50488 13676
rect 50448 13530 50476 13670
rect 50436 13524 50488 13530
rect 50436 13466 50488 13472
rect 50344 13456 50396 13462
rect 50344 13398 50396 13404
rect 50528 13456 50580 13462
rect 50528 13398 50580 13404
rect 50356 12238 50384 13398
rect 50436 13320 50488 13326
rect 50436 13262 50488 13268
rect 50448 12986 50476 13262
rect 50436 12980 50488 12986
rect 50436 12922 50488 12928
rect 50448 12782 50476 12922
rect 50436 12776 50488 12782
rect 50436 12718 50488 12724
rect 50434 12336 50490 12345
rect 50434 12271 50436 12280
rect 50488 12271 50490 12280
rect 50436 12242 50488 12248
rect 50252 12232 50304 12238
rect 50252 12174 50304 12180
rect 50344 12232 50396 12238
rect 50344 12174 50396 12180
rect 49976 11756 50028 11762
rect 49976 11698 50028 11704
rect 50080 11750 50200 11778
rect 50356 11762 50384 12174
rect 50344 11756 50396 11762
rect 49884 11620 49936 11626
rect 49884 11562 49936 11568
rect 49804 11478 49924 11506
rect 49792 11144 49844 11150
rect 49792 11086 49844 11092
rect 49700 10260 49752 10266
rect 49700 10202 49752 10208
rect 49804 10198 49832 11086
rect 49792 10192 49844 10198
rect 49792 10134 49844 10140
rect 49608 9988 49660 9994
rect 49608 9930 49660 9936
rect 49620 9738 49648 9930
rect 49700 9920 49752 9926
rect 49700 9862 49752 9868
rect 49436 9722 49648 9738
rect 49712 9722 49740 9862
rect 49424 9716 49648 9722
rect 49476 9710 49648 9716
rect 49700 9716 49752 9722
rect 49424 9658 49476 9664
rect 49700 9658 49752 9664
rect 49792 9716 49844 9722
rect 49792 9658 49844 9664
rect 49608 8424 49660 8430
rect 49608 8366 49660 8372
rect 49424 4276 49476 4282
rect 49424 4218 49476 4224
rect 49436 3126 49464 4218
rect 49620 3738 49648 8366
rect 49700 3936 49752 3942
rect 49700 3878 49752 3884
rect 49712 3738 49740 3878
rect 49608 3732 49660 3738
rect 49608 3674 49660 3680
rect 49700 3732 49752 3738
rect 49700 3674 49752 3680
rect 49700 3596 49752 3602
rect 49700 3538 49752 3544
rect 49514 3496 49570 3505
rect 49514 3431 49516 3440
rect 49568 3431 49570 3440
rect 49516 3402 49568 3408
rect 49424 3120 49476 3126
rect 49712 3074 49740 3538
rect 49424 3062 49476 3068
rect 49620 3058 49740 3074
rect 49608 3052 49740 3058
rect 49660 3046 49740 3052
rect 49608 2994 49660 3000
rect 49804 2961 49832 9658
rect 49896 6866 49924 11478
rect 49988 11286 50016 11698
rect 49976 11280 50028 11286
rect 49976 11222 50028 11228
rect 50080 11098 50108 11750
rect 50344 11698 50396 11704
rect 50252 11620 50304 11626
rect 50252 11562 50304 11568
rect 50160 11212 50212 11218
rect 50160 11154 50212 11160
rect 49988 11082 50108 11098
rect 49976 11076 50108 11082
rect 50028 11070 50108 11076
rect 49976 11018 50028 11024
rect 49976 10464 50028 10470
rect 49976 10406 50028 10412
rect 49988 10130 50016 10406
rect 49976 10124 50028 10130
rect 49976 10066 50028 10072
rect 50068 10056 50120 10062
rect 50068 9998 50120 10004
rect 50080 8838 50108 9998
rect 50172 9654 50200 11154
rect 50264 9674 50292 11562
rect 50356 11218 50384 11698
rect 50344 11212 50396 11218
rect 50344 11154 50396 11160
rect 50540 11150 50568 13398
rect 50620 12640 50672 12646
rect 50620 12582 50672 12588
rect 50632 11150 50660 12582
rect 50528 11144 50580 11150
rect 50528 11086 50580 11092
rect 50620 11144 50672 11150
rect 50620 11086 50672 11092
rect 50540 10674 50568 11086
rect 50528 10668 50580 10674
rect 50528 10610 50580 10616
rect 50528 9920 50580 9926
rect 50528 9862 50580 9868
rect 50160 9648 50212 9654
rect 50264 9646 50384 9674
rect 50540 9654 50568 9862
rect 50160 9590 50212 9596
rect 50172 8974 50200 9590
rect 50160 8968 50212 8974
rect 50160 8910 50212 8916
rect 50252 8968 50304 8974
rect 50252 8910 50304 8916
rect 50068 8832 50120 8838
rect 50068 8774 50120 8780
rect 50080 8634 50108 8774
rect 50068 8628 50120 8634
rect 50068 8570 50120 8576
rect 49884 6860 49936 6866
rect 49884 6802 49936 6808
rect 49976 4140 50028 4146
rect 49976 4082 50028 4088
rect 49790 2952 49846 2961
rect 49790 2887 49846 2896
rect 49344 2746 49464 2774
rect 49436 1358 49464 2746
rect 49988 2650 50016 4082
rect 50172 3602 50200 8910
rect 50264 8634 50292 8910
rect 50252 8628 50304 8634
rect 50252 8570 50304 8576
rect 50160 3596 50212 3602
rect 50160 3538 50212 3544
rect 50252 3528 50304 3534
rect 50252 3470 50304 3476
rect 50264 3369 50292 3470
rect 50250 3360 50306 3369
rect 50250 3295 50306 3304
rect 50264 3058 50292 3295
rect 50356 3194 50384 9646
rect 50528 9648 50580 9654
rect 50528 9590 50580 9596
rect 50632 8786 50660 11086
rect 50448 8758 50660 8786
rect 50344 3188 50396 3194
rect 50344 3130 50396 3136
rect 50252 3052 50304 3058
rect 50252 2994 50304 3000
rect 49976 2644 50028 2650
rect 49976 2586 50028 2592
rect 50252 2644 50304 2650
rect 50252 2586 50304 2592
rect 49608 2440 49660 2446
rect 49608 2382 49660 2388
rect 49424 1352 49476 1358
rect 49424 1294 49476 1300
rect 49620 800 49648 2382
rect 50264 800 50292 2586
rect 50356 2310 50384 3130
rect 50344 2304 50396 2310
rect 50344 2246 50396 2252
rect 50448 2038 50476 8758
rect 50724 7562 50752 14062
rect 50816 14062 50936 14090
rect 51000 14074 51028 14486
rect 51092 14414 51120 14758
rect 51080 14408 51132 14414
rect 51080 14350 51132 14356
rect 50988 14068 51040 14074
rect 50816 14006 50844 14062
rect 50988 14010 51040 14016
rect 50804 14000 50856 14006
rect 51000 13954 51028 14010
rect 50804 13942 50856 13948
rect 50908 13926 51028 13954
rect 50908 13682 50936 13926
rect 51092 13852 51120 14350
rect 50816 13654 50936 13682
rect 51000 13824 51120 13852
rect 50816 12918 50844 13654
rect 51000 13569 51028 13824
rect 51184 13682 51212 15456
rect 51264 15438 51316 15444
rect 51448 15496 51500 15502
rect 51448 15438 51500 15444
rect 51092 13654 51212 13682
rect 50986 13560 51042 13569
rect 50986 13495 51042 13504
rect 50894 13016 50950 13025
rect 50894 12951 50950 12960
rect 50804 12912 50856 12918
rect 50804 12854 50856 12860
rect 50804 12776 50856 12782
rect 50804 12718 50856 12724
rect 50816 10169 50844 12718
rect 50908 12714 50936 12951
rect 50988 12844 51040 12850
rect 50988 12786 51040 12792
rect 50896 12708 50948 12714
rect 50896 12650 50948 12656
rect 51000 12442 51028 12786
rect 50988 12436 51040 12442
rect 50988 12378 51040 12384
rect 51092 11914 51120 13654
rect 51170 13560 51226 13569
rect 51276 13530 51304 15438
rect 51460 15337 51488 15438
rect 51446 15328 51502 15337
rect 51446 15263 51502 15272
rect 51552 15094 51580 16050
rect 51540 15088 51592 15094
rect 51540 15030 51592 15036
rect 51356 14816 51408 14822
rect 51356 14758 51408 14764
rect 51368 14657 51396 14758
rect 51354 14648 51410 14657
rect 51538 14648 51594 14657
rect 51354 14583 51410 14592
rect 51460 14606 51538 14634
rect 51460 13938 51488 14606
rect 51538 14583 51594 14592
rect 51632 14612 51684 14618
rect 51632 14554 51684 14560
rect 51644 14521 51672 14554
rect 51630 14512 51686 14521
rect 51630 14447 51686 14456
rect 51736 13938 51764 27338
rect 52288 27334 52316 27610
rect 52380 27588 52408 29294
rect 52826 29200 52882 30000
rect 53470 29322 53526 30000
rect 54114 29322 54170 30000
rect 53470 29294 53604 29322
rect 53470 29200 53526 29294
rect 52460 27600 52512 27606
rect 52380 27560 52460 27588
rect 52460 27542 52512 27548
rect 52736 27396 52788 27402
rect 52736 27338 52788 27344
rect 52092 27328 52144 27334
rect 52092 27270 52144 27276
rect 52276 27328 52328 27334
rect 52276 27270 52328 27276
rect 51816 18284 51868 18290
rect 51816 18226 51868 18232
rect 51448 13932 51500 13938
rect 51448 13874 51500 13880
rect 51724 13932 51776 13938
rect 51724 13874 51776 13880
rect 51540 13864 51592 13870
rect 51540 13806 51592 13812
rect 51356 13796 51408 13802
rect 51356 13738 51408 13744
rect 51170 13495 51226 13504
rect 51264 13524 51316 13530
rect 51184 13297 51212 13495
rect 51264 13466 51316 13472
rect 51368 13410 51396 13738
rect 51552 13530 51580 13806
rect 51736 13530 51764 13874
rect 51540 13524 51592 13530
rect 51540 13466 51592 13472
rect 51724 13524 51776 13530
rect 51724 13466 51776 13472
rect 51276 13394 51396 13410
rect 51264 13388 51396 13394
rect 51316 13382 51396 13388
rect 51264 13330 51316 13336
rect 51552 13297 51580 13466
rect 51828 13326 51856 18226
rect 51906 16824 51962 16833
rect 51906 16759 51962 16768
rect 51920 16114 51948 16759
rect 52000 16516 52052 16522
rect 52000 16458 52052 16464
rect 52012 16250 52040 16458
rect 52000 16244 52052 16250
rect 52000 16186 52052 16192
rect 51908 16108 51960 16114
rect 51908 16050 51960 16056
rect 51998 15600 52054 15609
rect 51998 15535 52054 15544
rect 51908 15496 51960 15502
rect 51908 15438 51960 15444
rect 51816 13320 51868 13326
rect 51170 13288 51226 13297
rect 51170 13223 51226 13232
rect 51538 13288 51594 13297
rect 51816 13262 51868 13268
rect 51538 13223 51594 13232
rect 51632 13252 51684 13258
rect 51632 13194 51684 13200
rect 51644 13138 51672 13194
rect 51460 13110 51672 13138
rect 51460 12986 51488 13110
rect 51448 12980 51500 12986
rect 51448 12922 51500 12928
rect 51816 12844 51868 12850
rect 51816 12786 51868 12792
rect 51828 12714 51856 12786
rect 51816 12708 51868 12714
rect 51816 12650 51868 12656
rect 51354 12064 51410 12073
rect 51354 11999 51410 12008
rect 51000 11886 51120 11914
rect 51000 11234 51028 11886
rect 51080 11824 51132 11830
rect 51080 11766 51132 11772
rect 51092 11558 51120 11766
rect 51368 11762 51396 11999
rect 51356 11756 51408 11762
rect 51356 11698 51408 11704
rect 51080 11552 51132 11558
rect 51080 11494 51132 11500
rect 51264 11552 51316 11558
rect 51356 11552 51408 11558
rect 51264 11494 51316 11500
rect 51354 11520 51356 11529
rect 51408 11520 51410 11529
rect 51172 11348 51224 11354
rect 51276 11336 51304 11494
rect 51354 11455 51410 11464
rect 51224 11308 51304 11336
rect 51356 11348 51408 11354
rect 51172 11290 51224 11296
rect 51356 11290 51408 11296
rect 51000 11206 51212 11234
rect 50894 10976 50950 10985
rect 50894 10911 50950 10920
rect 50908 10674 50936 10911
rect 50896 10668 50948 10674
rect 50896 10610 50948 10616
rect 50802 10160 50858 10169
rect 50802 10095 50858 10104
rect 50908 10010 50936 10610
rect 50816 9982 50936 10010
rect 50988 10056 51040 10062
rect 50988 9998 51040 10004
rect 50816 9722 50844 9982
rect 51000 9722 51028 9998
rect 50804 9716 50856 9722
rect 50804 9658 50856 9664
rect 50988 9716 51040 9722
rect 50988 9658 51040 9664
rect 51184 9654 51212 11206
rect 51368 10985 51396 11290
rect 51354 10976 51410 10985
rect 51354 10911 51410 10920
rect 51356 10736 51408 10742
rect 51356 10678 51408 10684
rect 51368 10062 51396 10678
rect 51920 10266 51948 15438
rect 52012 15434 52040 15535
rect 52000 15428 52052 15434
rect 52000 15370 52052 15376
rect 52000 14476 52052 14482
rect 52000 14418 52052 14424
rect 52012 14074 52040 14418
rect 52000 14068 52052 14074
rect 52000 14010 52052 14016
rect 52000 13864 52052 13870
rect 52000 13806 52052 13812
rect 52012 11762 52040 13806
rect 52104 13394 52132 27270
rect 52748 27130 52776 27338
rect 52840 27130 52868 29200
rect 53576 27470 53604 29294
rect 54114 29294 54248 29322
rect 54114 29200 54170 29294
rect 52920 27464 52972 27470
rect 52920 27406 52972 27412
rect 53564 27464 53616 27470
rect 53564 27406 53616 27412
rect 54024 27464 54076 27470
rect 54024 27406 54076 27412
rect 52736 27124 52788 27130
rect 52736 27066 52788 27072
rect 52828 27124 52880 27130
rect 52828 27066 52880 27072
rect 52932 18426 52960 27406
rect 53196 27328 53248 27334
rect 53196 27270 53248 27276
rect 53208 27062 53236 27270
rect 53196 27056 53248 27062
rect 53196 26998 53248 27004
rect 53932 26988 53984 26994
rect 53932 26930 53984 26936
rect 53944 24274 53972 26930
rect 53932 24268 53984 24274
rect 53932 24210 53984 24216
rect 52920 18420 52972 18426
rect 52920 18362 52972 18368
rect 53840 18148 53892 18154
rect 53840 18090 53892 18096
rect 53012 17740 53064 17746
rect 53012 17682 53064 17688
rect 53104 17740 53156 17746
rect 53104 17682 53156 17688
rect 52184 17672 52236 17678
rect 53024 17649 53052 17682
rect 52184 17614 52236 17620
rect 53010 17640 53066 17649
rect 52196 14804 52224 17614
rect 53116 17610 53144 17682
rect 53288 17672 53340 17678
rect 53288 17614 53340 17620
rect 53010 17575 53066 17584
rect 53104 17604 53156 17610
rect 53104 17546 53156 17552
rect 52828 16720 52880 16726
rect 52828 16662 52880 16668
rect 52368 16584 52420 16590
rect 52368 16526 52420 16532
rect 52552 16584 52604 16590
rect 52736 16584 52788 16590
rect 52552 16526 52604 16532
rect 52656 16544 52736 16572
rect 52380 15706 52408 16526
rect 52460 16516 52512 16522
rect 52460 16458 52512 16464
rect 52472 16250 52500 16458
rect 52460 16244 52512 16250
rect 52460 16186 52512 16192
rect 52460 16108 52512 16114
rect 52460 16050 52512 16056
rect 52368 15700 52420 15706
rect 52368 15642 52420 15648
rect 52274 15600 52330 15609
rect 52274 15535 52330 15544
rect 52288 15502 52316 15535
rect 52276 15496 52328 15502
rect 52276 15438 52328 15444
rect 52288 14929 52316 15438
rect 52274 14920 52330 14929
rect 52274 14855 52330 14864
rect 52196 14776 52316 14804
rect 52184 14476 52236 14482
rect 52184 14418 52236 14424
rect 52196 14385 52224 14418
rect 52182 14376 52238 14385
rect 52182 14311 52238 14320
rect 52288 14113 52316 14776
rect 52472 14385 52500 16050
rect 52564 15586 52592 16526
rect 52656 16046 52684 16544
rect 52840 16561 52868 16662
rect 52736 16526 52788 16532
rect 52826 16552 52882 16561
rect 52826 16487 52882 16496
rect 53104 16516 53156 16522
rect 53104 16458 53156 16464
rect 53116 16250 53144 16458
rect 53194 16280 53250 16289
rect 53104 16244 53156 16250
rect 53194 16215 53196 16224
rect 53104 16186 53156 16192
rect 53248 16215 53250 16224
rect 53196 16186 53248 16192
rect 52828 16108 52880 16114
rect 52828 16050 52880 16056
rect 52644 16040 52696 16046
rect 52840 16017 52868 16050
rect 52644 15982 52696 15988
rect 52826 16008 52882 16017
rect 52826 15943 52882 15952
rect 53116 15638 53144 16186
rect 53196 16108 53248 16114
rect 53196 16050 53248 16056
rect 53104 15632 53156 15638
rect 52564 15558 52684 15586
rect 53104 15574 53156 15580
rect 52552 15496 52604 15502
rect 52552 15438 52604 15444
rect 52564 15337 52592 15438
rect 52550 15328 52606 15337
rect 52550 15263 52606 15272
rect 52656 14890 52684 15558
rect 53208 15201 53236 16050
rect 53300 15502 53328 17614
rect 53380 17536 53432 17542
rect 53380 17478 53432 17484
rect 53564 17536 53616 17542
rect 53564 17478 53616 17484
rect 53656 17536 53708 17542
rect 53656 17478 53708 17484
rect 53392 17184 53420 17478
rect 53472 17196 53524 17202
rect 53392 17156 53472 17184
rect 53472 17138 53524 17144
rect 53470 16960 53526 16969
rect 53470 16895 53526 16904
rect 53484 16658 53512 16895
rect 53472 16652 53524 16658
rect 53472 16594 53524 16600
rect 53380 16584 53432 16590
rect 53380 16526 53432 16532
rect 53392 15706 53420 16526
rect 53470 15736 53526 15745
rect 53380 15700 53432 15706
rect 53470 15671 53526 15680
rect 53380 15642 53432 15648
rect 53288 15496 53340 15502
rect 53288 15438 53340 15444
rect 53194 15192 53250 15201
rect 53104 15156 53156 15162
rect 53194 15127 53250 15136
rect 53104 15098 53156 15104
rect 52920 15088 52972 15094
rect 52920 15030 52972 15036
rect 52644 14884 52696 14890
rect 52644 14826 52696 14832
rect 52826 14512 52882 14521
rect 52826 14447 52882 14456
rect 52458 14376 52514 14385
rect 52458 14311 52514 14320
rect 52274 14104 52330 14113
rect 52274 14039 52330 14048
rect 52092 13388 52144 13394
rect 52092 13330 52144 13336
rect 52184 13320 52236 13326
rect 52104 13268 52184 13274
rect 52104 13262 52236 13268
rect 52104 13246 52224 13262
rect 52104 12918 52132 13246
rect 52092 12912 52144 12918
rect 52092 12854 52144 12860
rect 52184 12912 52236 12918
rect 52184 12854 52236 12860
rect 52092 12164 52144 12170
rect 52092 12106 52144 12112
rect 52104 11898 52132 12106
rect 52092 11892 52144 11898
rect 52092 11834 52144 11840
rect 52000 11756 52052 11762
rect 52000 11698 52052 11704
rect 52092 10600 52144 10606
rect 52092 10542 52144 10548
rect 52104 10305 52132 10542
rect 52090 10296 52146 10305
rect 51908 10260 51960 10266
rect 52090 10231 52146 10240
rect 51908 10202 51960 10208
rect 52196 10062 52224 12854
rect 52288 12850 52316 14039
rect 52736 14000 52788 14006
rect 52736 13942 52788 13948
rect 52366 13832 52422 13841
rect 52366 13767 52422 13776
rect 52276 12844 52328 12850
rect 52276 12786 52328 12792
rect 52380 12714 52408 13767
rect 52460 13252 52512 13258
rect 52460 13194 52512 13200
rect 52368 12708 52420 12714
rect 52368 12650 52420 12656
rect 52472 11234 52500 13194
rect 52552 13184 52604 13190
rect 52552 13126 52604 13132
rect 52748 13138 52776 13942
rect 52840 13326 52868 14447
rect 52932 14414 52960 15030
rect 53116 14929 53144 15098
rect 53484 15026 53512 15671
rect 53576 15434 53604 17478
rect 53668 17270 53696 17478
rect 53656 17264 53708 17270
rect 53656 17206 53708 17212
rect 53852 17066 53880 18090
rect 53932 17672 53984 17678
rect 53932 17614 53984 17620
rect 53944 17202 53972 17614
rect 53932 17196 53984 17202
rect 53932 17138 53984 17144
rect 53748 17060 53800 17066
rect 53748 17002 53800 17008
rect 53840 17060 53892 17066
rect 53840 17002 53892 17008
rect 53760 16402 53788 17002
rect 53932 16992 53984 16998
rect 53932 16934 53984 16940
rect 53944 16590 53972 16934
rect 53932 16584 53984 16590
rect 53932 16526 53984 16532
rect 53760 16374 53972 16402
rect 53746 16280 53802 16289
rect 53746 16215 53802 16224
rect 53760 16182 53788 16215
rect 53748 16176 53800 16182
rect 53748 16118 53800 16124
rect 53944 16114 53972 16374
rect 53932 16108 53984 16114
rect 53932 16050 53984 16056
rect 53944 16017 53972 16050
rect 53930 16008 53986 16017
rect 53930 15943 53986 15952
rect 53840 15904 53892 15910
rect 53840 15846 53892 15852
rect 53748 15564 53800 15570
rect 53748 15506 53800 15512
rect 53760 15434 53788 15506
rect 53564 15428 53616 15434
rect 53564 15370 53616 15376
rect 53748 15428 53800 15434
rect 53748 15370 53800 15376
rect 53852 15094 53880 15846
rect 53840 15088 53892 15094
rect 53840 15030 53892 15036
rect 53288 15020 53340 15026
rect 53288 14962 53340 14968
rect 53472 15020 53524 15026
rect 53472 14962 53524 14968
rect 53102 14920 53158 14929
rect 53102 14855 53158 14864
rect 53300 14618 53328 14962
rect 53288 14612 53340 14618
rect 53288 14554 53340 14560
rect 52920 14408 52972 14414
rect 52920 14350 52972 14356
rect 53932 14340 53984 14346
rect 53932 14282 53984 14288
rect 52918 13832 52974 13841
rect 52918 13767 52920 13776
rect 52972 13767 52974 13776
rect 52920 13738 52972 13744
rect 53472 13388 53524 13394
rect 53472 13330 53524 13336
rect 52828 13320 52880 13326
rect 52828 13262 52880 13268
rect 52564 12646 52592 13126
rect 52748 13110 53052 13138
rect 53024 13025 53052 13110
rect 52826 13016 52882 13025
rect 52826 12951 52828 12960
rect 52880 12951 52882 12960
rect 53010 13016 53066 13025
rect 53010 12951 53066 12960
rect 52828 12922 52880 12928
rect 52828 12844 52880 12850
rect 52828 12786 52880 12792
rect 53104 12844 53156 12850
rect 53104 12786 53156 12792
rect 53196 12844 53248 12850
rect 53196 12786 53248 12792
rect 52736 12776 52788 12782
rect 52736 12718 52788 12724
rect 52552 12640 52604 12646
rect 52552 12582 52604 12588
rect 52748 11898 52776 12718
rect 52840 12102 52868 12786
rect 53010 12472 53066 12481
rect 53116 12442 53144 12786
rect 53010 12407 53066 12416
rect 53104 12436 53156 12442
rect 52918 12200 52974 12209
rect 52918 12135 52974 12144
rect 52828 12096 52880 12102
rect 52828 12038 52880 12044
rect 52736 11892 52788 11898
rect 52736 11834 52788 11840
rect 52840 11762 52868 12038
rect 52828 11756 52880 11762
rect 52828 11698 52880 11704
rect 52932 11558 52960 12135
rect 52920 11552 52972 11558
rect 52920 11494 52972 11500
rect 52276 11212 52328 11218
rect 52472 11206 52868 11234
rect 52276 11154 52328 11160
rect 52288 11121 52316 11154
rect 52274 11112 52330 11121
rect 52840 11082 52868 11206
rect 52274 11047 52330 11056
rect 52736 11076 52788 11082
rect 52736 11018 52788 11024
rect 52828 11076 52880 11082
rect 52828 11018 52880 11024
rect 52642 10568 52698 10577
rect 52552 10532 52604 10538
rect 52748 10538 52776 11018
rect 52642 10503 52698 10512
rect 52736 10532 52788 10538
rect 52552 10474 52604 10480
rect 52564 10441 52592 10474
rect 52550 10432 52606 10441
rect 52550 10367 52606 10376
rect 51356 10056 51408 10062
rect 51356 9998 51408 10004
rect 52184 10056 52236 10062
rect 52184 9998 52236 10004
rect 51172 9648 51224 9654
rect 51172 9590 51224 9596
rect 52656 9382 52684 10503
rect 52736 10474 52788 10480
rect 52736 9580 52788 9586
rect 52736 9522 52788 9528
rect 52644 9376 52696 9382
rect 52644 9318 52696 9324
rect 52748 9042 52776 9522
rect 52736 9036 52788 9042
rect 52736 8978 52788 8984
rect 52368 8968 52420 8974
rect 52368 8910 52420 8916
rect 50804 8832 50856 8838
rect 50804 8774 50856 8780
rect 50816 8362 50844 8774
rect 52380 8634 52408 8910
rect 52368 8628 52420 8634
rect 52368 8570 52420 8576
rect 50804 8356 50856 8362
rect 50804 8298 50856 8304
rect 50724 7534 50844 7562
rect 50712 4820 50764 4826
rect 50712 4762 50764 4768
rect 50528 3528 50580 3534
rect 50526 3496 50528 3505
rect 50580 3496 50582 3505
rect 50526 3431 50582 3440
rect 50618 2816 50674 2825
rect 50618 2751 50674 2760
rect 50632 2310 50660 2751
rect 50724 2514 50752 4762
rect 50712 2508 50764 2514
rect 50712 2450 50764 2456
rect 50620 2304 50672 2310
rect 50620 2246 50672 2252
rect 50632 2038 50660 2246
rect 50436 2032 50488 2038
rect 50436 1974 50488 1980
rect 50620 2032 50672 2038
rect 50620 1974 50672 1980
rect 50816 1426 50844 7534
rect 51448 4820 51500 4826
rect 51448 4762 51500 4768
rect 51460 4214 51488 4762
rect 51448 4208 51500 4214
rect 51448 4150 51500 4156
rect 51816 4208 51868 4214
rect 51816 4150 51868 4156
rect 51448 4072 51500 4078
rect 51446 4040 51448 4049
rect 51500 4040 51502 4049
rect 51446 3975 51502 3984
rect 51632 3936 51684 3942
rect 51632 3878 51684 3884
rect 51356 3664 51408 3670
rect 51356 3606 51408 3612
rect 51368 3534 51396 3606
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 51448 3460 51500 3466
rect 51448 3402 51500 3408
rect 51460 2922 51488 3402
rect 51644 3058 51672 3878
rect 51828 3505 51856 4150
rect 51908 4072 51960 4078
rect 51908 4014 51960 4020
rect 52550 4040 52606 4049
rect 51814 3496 51870 3505
rect 51814 3431 51870 3440
rect 51632 3052 51684 3058
rect 51632 2994 51684 3000
rect 51724 2984 51776 2990
rect 51724 2926 51776 2932
rect 51448 2916 51500 2922
rect 51448 2858 51500 2864
rect 51736 2774 51764 2926
rect 51920 2922 51948 4014
rect 52550 3975 52606 3984
rect 52564 3602 52592 3975
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 52918 3496 52974 3505
rect 52918 3431 52974 3440
rect 52932 3398 52960 3431
rect 52920 3392 52972 3398
rect 52182 3360 52238 3369
rect 52920 3334 52972 3340
rect 52182 3295 52238 3304
rect 51998 3224 52054 3233
rect 52196 3194 52224 3295
rect 51998 3159 52000 3168
rect 52052 3159 52054 3168
rect 52184 3188 52236 3194
rect 52000 3130 52052 3136
rect 52184 3130 52236 3136
rect 51908 2916 51960 2922
rect 51908 2858 51960 2864
rect 52184 2916 52236 2922
rect 52184 2858 52236 2864
rect 51552 2746 51764 2774
rect 50988 2508 51040 2514
rect 50988 2450 51040 2456
rect 50896 2372 50948 2378
rect 50896 2314 50948 2320
rect 50804 1420 50856 1426
rect 50804 1362 50856 1368
rect 50908 800 50936 2314
rect 51000 2310 51028 2450
rect 50988 2304 51040 2310
rect 50988 2246 51040 2252
rect 51448 2304 51500 2310
rect 51448 2246 51500 2252
rect 51460 1494 51488 2246
rect 51448 1488 51500 1494
rect 51448 1430 51500 1436
rect 51552 800 51580 2746
rect 51632 2032 51684 2038
rect 51632 1974 51684 1980
rect 51644 1426 51672 1974
rect 51632 1420 51684 1426
rect 51632 1362 51684 1368
rect 52196 800 52224 2858
rect 52828 2372 52880 2378
rect 52828 2314 52880 2320
rect 52840 800 52868 2314
rect 52932 2038 52960 3334
rect 53024 2774 53052 12407
rect 53104 12378 53156 12384
rect 53208 11898 53236 12786
rect 53300 12782 53328 12813
rect 53288 12776 53340 12782
rect 53286 12744 53288 12753
rect 53340 12744 53342 12753
rect 53286 12679 53342 12688
rect 53300 12442 53328 12679
rect 53378 12472 53434 12481
rect 53288 12436 53340 12442
rect 53378 12407 53434 12416
rect 53288 12378 53340 12384
rect 53392 12374 53420 12407
rect 53380 12368 53432 12374
rect 53380 12310 53432 12316
rect 53196 11892 53248 11898
rect 53196 11834 53248 11840
rect 53380 11892 53432 11898
rect 53380 11834 53432 11840
rect 53104 11552 53156 11558
rect 53104 11494 53156 11500
rect 53116 11150 53144 11494
rect 53104 11144 53156 11150
rect 53104 11086 53156 11092
rect 53392 10849 53420 11834
rect 53378 10840 53434 10849
rect 53378 10775 53434 10784
rect 53104 10668 53156 10674
rect 53104 10610 53156 10616
rect 53116 10470 53144 10610
rect 53484 10577 53512 13330
rect 53944 13258 53972 14282
rect 53932 13252 53984 13258
rect 53576 13212 53932 13240
rect 53576 12238 53604 13212
rect 53932 13194 53984 13200
rect 53656 12844 53708 12850
rect 53840 12844 53892 12850
rect 53708 12804 53788 12832
rect 53656 12786 53708 12792
rect 53760 12345 53788 12804
rect 53840 12786 53892 12792
rect 53852 12374 53880 12786
rect 53932 12436 53984 12442
rect 53932 12378 53984 12384
rect 53840 12368 53892 12374
rect 53746 12336 53802 12345
rect 53840 12310 53892 12316
rect 53746 12271 53802 12280
rect 53564 12232 53616 12238
rect 53564 12174 53616 12180
rect 53760 12170 53788 12271
rect 53748 12164 53800 12170
rect 53800 12124 53880 12152
rect 53748 12106 53800 12112
rect 53656 12096 53708 12102
rect 53656 12038 53708 12044
rect 53668 11744 53696 12038
rect 53748 11756 53800 11762
rect 53668 11716 53748 11744
rect 53748 11698 53800 11704
rect 53760 10985 53788 11698
rect 53852 11529 53880 12124
rect 53944 12102 53972 12378
rect 53932 12096 53984 12102
rect 53932 12038 53984 12044
rect 53932 11756 53984 11762
rect 53932 11698 53984 11704
rect 53838 11520 53894 11529
rect 53838 11455 53894 11464
rect 53838 11384 53894 11393
rect 53838 11319 53894 11328
rect 53746 10976 53802 10985
rect 53746 10911 53802 10920
rect 53654 10840 53710 10849
rect 53654 10775 53710 10784
rect 53470 10568 53526 10577
rect 53470 10503 53526 10512
rect 53104 10464 53156 10470
rect 53104 10406 53156 10412
rect 53288 10464 53340 10470
rect 53288 10406 53340 10412
rect 53104 10192 53156 10198
rect 53104 10134 53156 10140
rect 53116 10062 53144 10134
rect 53104 10056 53156 10062
rect 53104 9998 53156 10004
rect 53300 9586 53328 10406
rect 53288 9580 53340 9586
rect 53288 9522 53340 9528
rect 53104 9376 53156 9382
rect 53104 9318 53156 9324
rect 53116 8838 53144 9318
rect 53104 8832 53156 8838
rect 53104 8774 53156 8780
rect 53116 8634 53144 8774
rect 53104 8628 53156 8634
rect 53104 8570 53156 8576
rect 53196 6860 53248 6866
rect 53196 6802 53248 6808
rect 53104 4480 53156 4486
rect 53104 4422 53156 4428
rect 53116 4282 53144 4422
rect 53104 4276 53156 4282
rect 53104 4218 53156 4224
rect 53208 3466 53236 6802
rect 53196 3460 53248 3466
rect 53196 3402 53248 3408
rect 53668 3058 53696 10775
rect 53748 10600 53800 10606
rect 53748 10542 53800 10548
rect 53760 10130 53788 10542
rect 53852 10130 53880 11319
rect 53944 11286 53972 11698
rect 53932 11280 53984 11286
rect 53932 11222 53984 11228
rect 53748 10124 53800 10130
rect 53748 10066 53800 10072
rect 53840 10124 53892 10130
rect 53840 10066 53892 10072
rect 53760 9654 53788 10066
rect 53748 9648 53800 9654
rect 53748 9590 53800 9596
rect 54036 4146 54064 27406
rect 54220 26994 54248 29294
rect 54758 29200 54814 30000
rect 56046 29322 56102 30000
rect 56690 29322 56746 30000
rect 56046 29294 56272 29322
rect 56046 29200 56102 29294
rect 55820 27772 56128 27781
rect 55820 27770 55826 27772
rect 55882 27770 55906 27772
rect 55962 27770 55986 27772
rect 56042 27770 56066 27772
rect 56122 27770 56128 27772
rect 55882 27718 55884 27770
rect 56064 27718 56066 27770
rect 55820 27716 55826 27718
rect 55882 27716 55906 27718
rect 55962 27716 55986 27718
rect 56042 27716 56066 27718
rect 56122 27716 56128 27718
rect 55820 27707 56128 27716
rect 56244 27606 56272 29294
rect 56690 29294 56824 29322
rect 56690 29200 56746 29294
rect 56796 27606 56824 29294
rect 57334 29200 57390 30000
rect 57978 29200 58034 30000
rect 58622 29322 58678 30000
rect 58622 29294 58848 29322
rect 58622 29200 58678 29294
rect 57348 27606 57376 29200
rect 55680 27600 55732 27606
rect 55680 27542 55732 27548
rect 56232 27600 56284 27606
rect 56232 27542 56284 27548
rect 56784 27600 56836 27606
rect 56784 27542 56836 27548
rect 57336 27600 57388 27606
rect 57336 27542 57388 27548
rect 54300 27328 54352 27334
rect 54300 27270 54352 27276
rect 54208 26988 54260 26994
rect 54208 26930 54260 26936
rect 54312 26926 54340 27270
rect 55496 26988 55548 26994
rect 55496 26930 55548 26936
rect 54300 26920 54352 26926
rect 54300 26862 54352 26868
rect 54484 26920 54536 26926
rect 54484 26862 54536 26868
rect 54496 22778 54524 26862
rect 54760 26580 54812 26586
rect 54760 26522 54812 26528
rect 54484 22772 54536 22778
rect 54484 22714 54536 22720
rect 54772 18358 54800 26522
rect 54760 18352 54812 18358
rect 54760 18294 54812 18300
rect 55128 18284 55180 18290
rect 55128 18226 55180 18232
rect 55404 18284 55456 18290
rect 55404 18226 55456 18232
rect 55140 18154 55168 18226
rect 55128 18148 55180 18154
rect 55128 18090 55180 18096
rect 54392 18080 54444 18086
rect 54392 18022 54444 18028
rect 54300 17808 54352 17814
rect 54300 17750 54352 17756
rect 54116 17672 54168 17678
rect 54116 17614 54168 17620
rect 54128 16522 54156 17614
rect 54208 17264 54260 17270
rect 54208 17206 54260 17212
rect 54116 16516 54168 16522
rect 54116 16458 54168 16464
rect 54220 16046 54248 17206
rect 54312 16454 54340 17750
rect 54404 17270 54432 18022
rect 55312 17808 55364 17814
rect 55310 17776 55312 17785
rect 55364 17776 55366 17785
rect 55416 17746 55444 18226
rect 55310 17711 55366 17720
rect 55404 17740 55456 17746
rect 55404 17682 55456 17688
rect 54576 17672 54628 17678
rect 54576 17614 54628 17620
rect 54668 17672 54720 17678
rect 54668 17614 54720 17620
rect 55312 17672 55364 17678
rect 55312 17614 55364 17620
rect 54482 17368 54538 17377
rect 54482 17303 54538 17312
rect 54496 17270 54524 17303
rect 54392 17264 54444 17270
rect 54392 17206 54444 17212
rect 54484 17264 54536 17270
rect 54484 17206 54536 17212
rect 54588 16572 54616 17614
rect 54680 16969 54708 17614
rect 55324 17134 55352 17614
rect 55312 17128 55364 17134
rect 55312 17070 55364 17076
rect 55128 17060 55180 17066
rect 55128 17002 55180 17008
rect 54666 16960 54722 16969
rect 54666 16895 54722 16904
rect 55140 16726 55168 17002
rect 55220 16992 55272 16998
rect 55220 16934 55272 16940
rect 55312 16992 55364 16998
rect 55312 16934 55364 16940
rect 55128 16720 55180 16726
rect 55128 16662 55180 16668
rect 55232 16658 55260 16934
rect 55220 16652 55272 16658
rect 55220 16594 55272 16600
rect 54760 16584 54812 16590
rect 54588 16544 54760 16572
rect 54760 16526 54812 16532
rect 54392 16516 54444 16522
rect 54392 16458 54444 16464
rect 54300 16448 54352 16454
rect 54300 16390 54352 16396
rect 54208 16040 54260 16046
rect 54208 15982 54260 15988
rect 54116 15632 54168 15638
rect 54116 15574 54168 15580
rect 54128 14414 54156 15574
rect 54220 15026 54248 15982
rect 54300 15156 54352 15162
rect 54300 15098 54352 15104
rect 54208 15020 54260 15026
rect 54208 14962 54260 14968
rect 54220 14793 54248 14962
rect 54312 14929 54340 15098
rect 54298 14920 54354 14929
rect 54298 14855 54354 14864
rect 54300 14816 54352 14822
rect 54206 14784 54262 14793
rect 54300 14758 54352 14764
rect 54206 14719 54262 14728
rect 54116 14408 54168 14414
rect 54116 14350 54168 14356
rect 54128 13870 54156 14350
rect 54116 13864 54168 13870
rect 54116 13806 54168 13812
rect 54128 13326 54156 13806
rect 54116 13320 54168 13326
rect 54116 13262 54168 13268
rect 54116 13184 54168 13190
rect 54116 13126 54168 13132
rect 54128 13025 54156 13126
rect 54114 13016 54170 13025
rect 54114 12951 54170 12960
rect 54220 11830 54248 14719
rect 54312 12238 54340 14758
rect 54404 14618 54432 16458
rect 54482 16416 54538 16425
rect 54482 16351 54538 16360
rect 54496 15026 54524 16351
rect 54576 16108 54628 16114
rect 54576 16050 54628 16056
rect 54484 15020 54536 15026
rect 54484 14962 54536 14968
rect 54392 14612 54444 14618
rect 54392 14554 54444 14560
rect 54390 14512 54446 14521
rect 54496 14482 54524 14962
rect 54390 14447 54446 14456
rect 54484 14476 54536 14482
rect 54404 13734 54432 14447
rect 54484 14418 54536 14424
rect 54588 14006 54616 16050
rect 54772 15745 54800 16526
rect 54944 16176 54996 16182
rect 54944 16118 54996 16124
rect 54956 15881 54984 16118
rect 55232 16114 55260 16594
rect 55324 16522 55352 16934
rect 55402 16824 55458 16833
rect 55402 16759 55458 16768
rect 55312 16516 55364 16522
rect 55312 16458 55364 16464
rect 55220 16108 55272 16114
rect 55220 16050 55272 16056
rect 55036 15972 55088 15978
rect 55036 15914 55088 15920
rect 54942 15872 54998 15881
rect 54942 15807 54998 15816
rect 54758 15736 54814 15745
rect 54814 15694 54892 15722
rect 54758 15671 54814 15680
rect 54760 15360 54812 15366
rect 54760 15302 54812 15308
rect 54668 14816 54720 14822
rect 54668 14758 54720 14764
rect 54680 14414 54708 14758
rect 54668 14408 54720 14414
rect 54668 14350 54720 14356
rect 54576 14000 54628 14006
rect 54576 13942 54628 13948
rect 54392 13728 54444 13734
rect 54392 13670 54444 13676
rect 54668 13728 54720 13734
rect 54668 13670 54720 13676
rect 54392 13456 54444 13462
rect 54392 13398 54444 13404
rect 54404 13326 54432 13398
rect 54392 13320 54444 13326
rect 54392 13262 54444 13268
rect 54392 13184 54444 13190
rect 54392 13126 54444 13132
rect 54404 12646 54432 13126
rect 54484 12844 54536 12850
rect 54484 12786 54536 12792
rect 54392 12640 54444 12646
rect 54392 12582 54444 12588
rect 54300 12232 54352 12238
rect 54300 12174 54352 12180
rect 54404 11937 54432 12582
rect 54390 11928 54446 11937
rect 54390 11863 54446 11872
rect 54208 11824 54260 11830
rect 54208 11766 54260 11772
rect 54116 11756 54168 11762
rect 54116 11698 54168 11704
rect 54128 11558 54156 11698
rect 54116 11552 54168 11558
rect 54116 11494 54168 11500
rect 54496 10826 54524 12786
rect 54576 12776 54628 12782
rect 54576 12718 54628 12724
rect 54588 11082 54616 12718
rect 54680 12238 54708 13670
rect 54772 13025 54800 15302
rect 54864 14822 54892 15694
rect 54956 15094 54984 15807
rect 54944 15088 54996 15094
rect 54944 15030 54996 15036
rect 55048 14890 55076 15914
rect 55416 15638 55444 16759
rect 55508 16153 55536 26930
rect 55692 26586 55720 27542
rect 57060 27464 57112 27470
rect 57060 27406 57112 27412
rect 56968 27328 57020 27334
rect 56968 27270 57020 27276
rect 56980 26926 57008 27270
rect 57072 27130 57100 27406
rect 57992 27130 58020 29200
rect 58820 27470 58848 29294
rect 59266 29200 59322 30000
rect 59910 29200 59966 30000
rect 60554 29322 60610 30000
rect 61198 29322 61254 30000
rect 61842 29322 61898 30000
rect 60554 29294 60688 29322
rect 60554 29200 60610 29294
rect 59280 27588 59308 29200
rect 59924 27606 59952 29200
rect 59360 27600 59412 27606
rect 59280 27560 59360 27588
rect 59360 27542 59412 27548
rect 59912 27600 59964 27606
rect 59912 27542 59964 27548
rect 60556 27600 60608 27606
rect 60556 27542 60608 27548
rect 58808 27464 58860 27470
rect 58808 27406 58860 27412
rect 59636 27464 59688 27470
rect 59636 27406 59688 27412
rect 58624 27396 58676 27402
rect 58624 27338 58676 27344
rect 57060 27124 57112 27130
rect 57060 27066 57112 27072
rect 57980 27124 58032 27130
rect 57980 27066 58032 27072
rect 58440 26988 58492 26994
rect 58440 26930 58492 26936
rect 56968 26920 57020 26926
rect 56968 26862 57020 26868
rect 55820 26684 56128 26693
rect 55820 26682 55826 26684
rect 55882 26682 55906 26684
rect 55962 26682 55986 26684
rect 56042 26682 56066 26684
rect 56122 26682 56128 26684
rect 55882 26630 55884 26682
rect 56064 26630 56066 26682
rect 55820 26628 55826 26630
rect 55882 26628 55906 26630
rect 55962 26628 55986 26630
rect 56042 26628 56066 26630
rect 56122 26628 56128 26630
rect 55820 26619 56128 26628
rect 55680 26580 55732 26586
rect 55680 26522 55732 26528
rect 55588 26376 55640 26382
rect 55588 26318 55640 26324
rect 55600 17678 55628 26318
rect 58452 26314 58480 26930
rect 58440 26308 58492 26314
rect 58440 26250 58492 26256
rect 58532 25764 58584 25770
rect 58532 25706 58584 25712
rect 55820 25596 56128 25605
rect 55820 25594 55826 25596
rect 55882 25594 55906 25596
rect 55962 25594 55986 25596
rect 56042 25594 56066 25596
rect 56122 25594 56128 25596
rect 55882 25542 55884 25594
rect 56064 25542 56066 25594
rect 55820 25540 55826 25542
rect 55882 25540 55906 25542
rect 55962 25540 55986 25542
rect 56042 25540 56066 25542
rect 56122 25540 56128 25542
rect 55820 25531 56128 25540
rect 55820 24508 56128 24517
rect 55820 24506 55826 24508
rect 55882 24506 55906 24508
rect 55962 24506 55986 24508
rect 56042 24506 56066 24508
rect 56122 24506 56128 24508
rect 55882 24454 55884 24506
rect 56064 24454 56066 24506
rect 55820 24452 55826 24454
rect 55882 24452 55906 24454
rect 55962 24452 55986 24454
rect 56042 24452 56066 24454
rect 56122 24452 56128 24454
rect 55820 24443 56128 24452
rect 56692 24132 56744 24138
rect 56692 24074 56744 24080
rect 55820 23420 56128 23429
rect 55820 23418 55826 23420
rect 55882 23418 55906 23420
rect 55962 23418 55986 23420
rect 56042 23418 56066 23420
rect 56122 23418 56128 23420
rect 55882 23366 55884 23418
rect 56064 23366 56066 23418
rect 55820 23364 55826 23366
rect 55882 23364 55906 23366
rect 55962 23364 55986 23366
rect 56042 23364 56066 23366
rect 56122 23364 56128 23366
rect 55820 23355 56128 23364
rect 56324 22976 56376 22982
rect 56324 22918 56376 22924
rect 55820 22332 56128 22341
rect 55820 22330 55826 22332
rect 55882 22330 55906 22332
rect 55962 22330 55986 22332
rect 56042 22330 56066 22332
rect 56122 22330 56128 22332
rect 55882 22278 55884 22330
rect 56064 22278 56066 22330
rect 55820 22276 55826 22278
rect 55882 22276 55906 22278
rect 55962 22276 55986 22278
rect 56042 22276 56066 22278
rect 56122 22276 56128 22278
rect 55820 22267 56128 22276
rect 55820 21244 56128 21253
rect 55820 21242 55826 21244
rect 55882 21242 55906 21244
rect 55962 21242 55986 21244
rect 56042 21242 56066 21244
rect 56122 21242 56128 21244
rect 55882 21190 55884 21242
rect 56064 21190 56066 21242
rect 55820 21188 55826 21190
rect 55882 21188 55906 21190
rect 55962 21188 55986 21190
rect 56042 21188 56066 21190
rect 56122 21188 56128 21190
rect 55820 21179 56128 21188
rect 55820 20156 56128 20165
rect 55820 20154 55826 20156
rect 55882 20154 55906 20156
rect 55962 20154 55986 20156
rect 56042 20154 56066 20156
rect 56122 20154 56128 20156
rect 55882 20102 55884 20154
rect 56064 20102 56066 20154
rect 55820 20100 55826 20102
rect 55882 20100 55906 20102
rect 55962 20100 55986 20102
rect 56042 20100 56066 20102
rect 56122 20100 56128 20102
rect 55820 20091 56128 20100
rect 56336 19310 56364 22918
rect 56508 19372 56560 19378
rect 56508 19314 56560 19320
rect 56600 19372 56652 19378
rect 56600 19314 56652 19320
rect 56324 19304 56376 19310
rect 56324 19246 56376 19252
rect 55820 19068 56128 19077
rect 55820 19066 55826 19068
rect 55882 19066 55906 19068
rect 55962 19066 55986 19068
rect 56042 19066 56066 19068
rect 56122 19066 56128 19068
rect 55882 19014 55884 19066
rect 56064 19014 56066 19066
rect 55820 19012 55826 19014
rect 55882 19012 55906 19014
rect 55962 19012 55986 19014
rect 56042 19012 56066 19014
rect 56122 19012 56128 19014
rect 55820 19003 56128 19012
rect 56520 18766 56548 19314
rect 55956 18760 56008 18766
rect 55956 18702 56008 18708
rect 56508 18760 56560 18766
rect 56508 18702 56560 18708
rect 55968 18290 55996 18702
rect 56612 18630 56640 19314
rect 56704 18970 56732 24074
rect 57060 21140 57112 21146
rect 57060 21082 57112 21088
rect 56692 18964 56744 18970
rect 56692 18906 56744 18912
rect 56968 18760 57020 18766
rect 56968 18702 57020 18708
rect 56232 18624 56284 18630
rect 56232 18566 56284 18572
rect 56600 18624 56652 18630
rect 56600 18566 56652 18572
rect 56244 18426 56272 18566
rect 56232 18420 56284 18426
rect 56232 18362 56284 18368
rect 55956 18284 56008 18290
rect 55956 18226 56008 18232
rect 55680 18216 55732 18222
rect 55680 18158 55732 18164
rect 55692 17746 55720 18158
rect 55820 17980 56128 17989
rect 55820 17978 55826 17980
rect 55882 17978 55906 17980
rect 55962 17978 55986 17980
rect 56042 17978 56066 17980
rect 56122 17978 56128 17980
rect 55882 17926 55884 17978
rect 56064 17926 56066 17978
rect 55820 17924 55826 17926
rect 55882 17924 55906 17926
rect 55962 17924 55986 17926
rect 56042 17924 56066 17926
rect 56122 17924 56128 17926
rect 55820 17915 56128 17924
rect 55680 17740 55732 17746
rect 55680 17682 55732 17688
rect 55588 17672 55640 17678
rect 55588 17614 55640 17620
rect 56048 17672 56100 17678
rect 56048 17614 56100 17620
rect 56060 17134 56088 17614
rect 56048 17128 56100 17134
rect 56048 17070 56100 17076
rect 55820 16892 56128 16901
rect 55820 16890 55826 16892
rect 55882 16890 55906 16892
rect 55962 16890 55986 16892
rect 56042 16890 56066 16892
rect 56122 16890 56128 16892
rect 55882 16838 55884 16890
rect 56064 16838 56066 16890
rect 55820 16836 55826 16838
rect 55882 16836 55906 16838
rect 55962 16836 55986 16838
rect 56042 16836 56066 16838
rect 56122 16836 56128 16838
rect 55820 16827 56128 16836
rect 55494 16144 55550 16153
rect 55494 16079 55550 16088
rect 55678 16008 55734 16017
rect 55678 15943 55734 15952
rect 55404 15632 55456 15638
rect 55404 15574 55456 15580
rect 55692 15502 55720 15943
rect 55820 15804 56128 15813
rect 55820 15802 55826 15804
rect 55882 15802 55906 15804
rect 55962 15802 55986 15804
rect 56042 15802 56066 15804
rect 56122 15802 56128 15804
rect 55882 15750 55884 15802
rect 56064 15750 56066 15802
rect 55820 15748 55826 15750
rect 55882 15748 55906 15750
rect 55962 15748 55986 15750
rect 56042 15748 56066 15750
rect 56122 15748 56128 15750
rect 55820 15739 56128 15748
rect 56244 15502 56272 18362
rect 56322 18320 56378 18329
rect 56322 18255 56324 18264
rect 56376 18255 56378 18264
rect 56324 18226 56376 18232
rect 56414 18184 56470 18193
rect 56414 18119 56470 18128
rect 56324 18080 56376 18086
rect 56324 18022 56376 18028
rect 56336 17678 56364 18022
rect 56428 17814 56456 18119
rect 56416 17808 56468 17814
rect 56416 17750 56468 17756
rect 56324 17672 56376 17678
rect 56324 17614 56376 17620
rect 56874 17640 56930 17649
rect 56874 17575 56930 17584
rect 56416 17536 56468 17542
rect 56416 17478 56468 17484
rect 56600 17536 56652 17542
rect 56600 17478 56652 17484
rect 56324 17196 56376 17202
rect 56324 17138 56376 17144
rect 56336 17066 56364 17138
rect 56324 17060 56376 17066
rect 56324 17002 56376 17008
rect 56428 16454 56456 17478
rect 56508 16992 56560 16998
rect 56508 16934 56560 16940
rect 56520 16590 56548 16934
rect 56508 16584 56560 16590
rect 56508 16526 56560 16532
rect 56612 16522 56640 17478
rect 56782 17232 56838 17241
rect 56782 17167 56784 17176
rect 56836 17167 56838 17176
rect 56784 17138 56836 17144
rect 56888 16522 56916 17575
rect 56600 16516 56652 16522
rect 56600 16458 56652 16464
rect 56876 16516 56928 16522
rect 56876 16458 56928 16464
rect 56416 16448 56468 16454
rect 56416 16390 56468 16396
rect 56784 16448 56836 16454
rect 56784 16390 56836 16396
rect 56796 16114 56824 16390
rect 56784 16108 56836 16114
rect 56784 16050 56836 16056
rect 56324 16040 56376 16046
rect 56324 15982 56376 15988
rect 56598 16008 56654 16017
rect 56336 15609 56364 15982
rect 56598 15943 56654 15952
rect 56612 15910 56640 15943
rect 56600 15904 56652 15910
rect 56600 15846 56652 15852
rect 56322 15600 56378 15609
rect 56322 15535 56378 15544
rect 55680 15496 55732 15502
rect 55680 15438 55732 15444
rect 56232 15496 56284 15502
rect 56232 15438 56284 15444
rect 56508 15496 56560 15502
rect 56508 15438 56560 15444
rect 55128 15428 55180 15434
rect 55128 15370 55180 15376
rect 55140 15314 55168 15370
rect 55404 15360 55456 15366
rect 55140 15308 55404 15314
rect 55140 15302 55456 15308
rect 55140 15286 55444 15302
rect 55140 15094 55168 15286
rect 55128 15088 55180 15094
rect 55128 15030 55180 15036
rect 56324 15088 56376 15094
rect 56324 15030 56376 15036
rect 55680 15020 55732 15026
rect 55680 14962 55732 14968
rect 55036 14884 55088 14890
rect 55036 14826 55088 14832
rect 54852 14816 54904 14822
rect 54852 14758 54904 14764
rect 54852 14476 54904 14482
rect 54852 14418 54904 14424
rect 54944 14476 54996 14482
rect 54944 14418 54996 14424
rect 54864 13410 54892 14418
rect 54956 14249 54984 14418
rect 55220 14340 55272 14346
rect 55220 14282 55272 14288
rect 54942 14240 54998 14249
rect 54942 14175 54998 14184
rect 55126 14240 55182 14249
rect 55126 14175 55182 14184
rect 55036 13932 55088 13938
rect 55036 13874 55088 13880
rect 54944 13728 54996 13734
rect 54944 13670 54996 13676
rect 54956 13530 54984 13670
rect 55048 13530 55076 13874
rect 54944 13524 54996 13530
rect 54944 13466 54996 13472
rect 55036 13524 55088 13530
rect 55036 13466 55088 13472
rect 54864 13382 55076 13410
rect 54758 13016 54814 13025
rect 54758 12951 54814 12960
rect 55048 12434 55076 13382
rect 55140 13258 55168 14175
rect 55232 13870 55260 14282
rect 55692 14278 55720 14962
rect 55820 14716 56128 14725
rect 55820 14714 55826 14716
rect 55882 14714 55906 14716
rect 55962 14714 55986 14716
rect 56042 14714 56066 14716
rect 56122 14714 56128 14716
rect 55882 14662 55884 14714
rect 56064 14662 56066 14714
rect 55820 14660 55826 14662
rect 55882 14660 55906 14662
rect 55962 14660 55986 14662
rect 56042 14660 56066 14662
rect 56122 14660 56128 14662
rect 55820 14651 56128 14660
rect 55680 14272 55732 14278
rect 55680 14214 55732 14220
rect 55588 14000 55640 14006
rect 55588 13942 55640 13948
rect 55220 13864 55272 13870
rect 55220 13806 55272 13812
rect 55128 13252 55180 13258
rect 55128 13194 55180 13200
rect 55232 12832 55260 13806
rect 55312 13252 55364 13258
rect 55312 13194 55364 13200
rect 55324 12850 55352 13194
rect 55404 13184 55456 13190
rect 55404 13126 55456 13132
rect 54956 12406 55076 12434
rect 55140 12804 55260 12832
rect 55312 12844 55364 12850
rect 54668 12232 54720 12238
rect 54668 12174 54720 12180
rect 54760 12096 54812 12102
rect 54760 12038 54812 12044
rect 54852 12096 54904 12102
rect 54852 12038 54904 12044
rect 54666 11928 54722 11937
rect 54772 11898 54800 12038
rect 54666 11863 54668 11872
rect 54720 11863 54722 11872
rect 54760 11892 54812 11898
rect 54668 11834 54720 11840
rect 54760 11834 54812 11840
rect 54760 11688 54812 11694
rect 54760 11630 54812 11636
rect 54772 11082 54800 11630
rect 54864 11558 54892 12038
rect 54852 11552 54904 11558
rect 54852 11494 54904 11500
rect 54576 11076 54628 11082
rect 54576 11018 54628 11024
rect 54760 11076 54812 11082
rect 54760 11018 54812 11024
rect 54312 10798 54524 10826
rect 54312 10742 54340 10798
rect 54300 10736 54352 10742
rect 54300 10678 54352 10684
rect 54312 9722 54340 10678
rect 54484 10668 54536 10674
rect 54484 10610 54536 10616
rect 54392 9920 54444 9926
rect 54392 9862 54444 9868
rect 54300 9716 54352 9722
rect 54300 9658 54352 9664
rect 54404 9602 54432 9862
rect 54496 9722 54524 10610
rect 54576 9920 54628 9926
rect 54576 9862 54628 9868
rect 54588 9722 54616 9862
rect 54484 9716 54536 9722
rect 54484 9658 54536 9664
rect 54576 9716 54628 9722
rect 54576 9658 54628 9664
rect 54956 9602 54984 12406
rect 55140 12306 55168 12804
rect 55312 12786 55364 12792
rect 55312 12640 55364 12646
rect 55312 12582 55364 12588
rect 55324 12322 55352 12582
rect 55416 12442 55444 13126
rect 55600 12646 55628 13942
rect 55692 13870 55720 14214
rect 56232 14000 56284 14006
rect 56232 13942 56284 13948
rect 55680 13864 55732 13870
rect 55680 13806 55732 13812
rect 55678 13696 55734 13705
rect 55678 13631 55734 13640
rect 55692 13161 55720 13631
rect 55820 13628 56128 13637
rect 55820 13626 55826 13628
rect 55882 13626 55906 13628
rect 55962 13626 55986 13628
rect 56042 13626 56066 13628
rect 56122 13626 56128 13628
rect 55882 13574 55884 13626
rect 56064 13574 56066 13626
rect 55820 13572 55826 13574
rect 55882 13572 55906 13574
rect 55962 13572 55986 13574
rect 56042 13572 56066 13574
rect 56122 13572 56128 13574
rect 55820 13563 56128 13572
rect 56048 13252 56100 13258
rect 56048 13194 56100 13200
rect 55678 13152 55734 13161
rect 55678 13087 55734 13096
rect 56060 13025 56088 13194
rect 56140 13184 56192 13190
rect 56140 13126 56192 13132
rect 56046 13016 56102 13025
rect 55956 12980 56008 12986
rect 56046 12951 56102 12960
rect 55956 12922 56008 12928
rect 55680 12844 55732 12850
rect 55680 12786 55732 12792
rect 55588 12640 55640 12646
rect 55588 12582 55640 12588
rect 55404 12436 55456 12442
rect 55404 12378 55456 12384
rect 55232 12306 55352 12322
rect 55128 12300 55180 12306
rect 55128 12242 55180 12248
rect 55220 12300 55352 12306
rect 55272 12294 55352 12300
rect 55600 12288 55628 12582
rect 55692 12434 55720 12786
rect 55968 12646 55996 12922
rect 56152 12782 56180 13126
rect 56140 12776 56192 12782
rect 56140 12718 56192 12724
rect 55956 12640 56008 12646
rect 55956 12582 56008 12588
rect 55820 12540 56128 12549
rect 55820 12538 55826 12540
rect 55882 12538 55906 12540
rect 55962 12538 55986 12540
rect 56042 12538 56066 12540
rect 56122 12538 56128 12540
rect 55882 12486 55884 12538
rect 56064 12486 56066 12538
rect 55820 12484 55826 12486
rect 55882 12484 55906 12486
rect 55962 12484 55986 12486
rect 56042 12484 56066 12486
rect 56122 12484 56128 12486
rect 55820 12475 56128 12484
rect 55692 12406 55812 12434
rect 55220 12242 55272 12248
rect 55508 12260 55628 12288
rect 55404 12232 55456 12238
rect 55508 12220 55536 12260
rect 55456 12192 55536 12220
rect 55404 12174 55456 12180
rect 55220 11756 55272 11762
rect 55220 11698 55272 11704
rect 55128 11688 55180 11694
rect 55128 11630 55180 11636
rect 55140 11354 55168 11630
rect 55232 11529 55260 11698
rect 55218 11520 55274 11529
rect 55218 11455 55274 11464
rect 55128 11348 55180 11354
rect 55128 11290 55180 11296
rect 55508 11218 55536 12192
rect 55588 12164 55640 12170
rect 55588 12106 55640 12112
rect 55600 11354 55628 12106
rect 55784 11762 55812 12406
rect 55772 11756 55824 11762
rect 55772 11698 55824 11704
rect 55820 11452 56128 11461
rect 55820 11450 55826 11452
rect 55882 11450 55906 11452
rect 55962 11450 55986 11452
rect 56042 11450 56066 11452
rect 56122 11450 56128 11452
rect 55882 11398 55884 11450
rect 56064 11398 56066 11450
rect 55820 11396 55826 11398
rect 55882 11396 55906 11398
rect 55962 11396 55986 11398
rect 56042 11396 56066 11398
rect 56122 11396 56128 11398
rect 55820 11387 56128 11396
rect 55588 11348 55640 11354
rect 55588 11290 55640 11296
rect 55496 11212 55548 11218
rect 55324 11172 55496 11200
rect 55220 11144 55272 11150
rect 55218 11112 55220 11121
rect 55272 11112 55274 11121
rect 55218 11047 55274 11056
rect 55220 10192 55272 10198
rect 55220 10134 55272 10140
rect 55036 10124 55088 10130
rect 55036 10066 55088 10072
rect 55048 9654 55076 10066
rect 54404 9574 54984 9602
rect 55036 9648 55088 9654
rect 55036 9590 55088 9596
rect 54024 4140 54076 4146
rect 54024 4082 54076 4088
rect 53656 3052 53708 3058
rect 53656 2994 53708 3000
rect 54956 2990 54984 9574
rect 55232 8974 55260 10134
rect 55324 10130 55352 11172
rect 55496 11154 55548 11160
rect 56244 11150 56272 13942
rect 56048 11144 56100 11150
rect 56048 11086 56100 11092
rect 56232 11144 56284 11150
rect 56232 11086 56284 11092
rect 56060 10962 56088 11086
rect 56060 10934 56272 10962
rect 55680 10600 55732 10606
rect 55680 10542 55732 10548
rect 55404 10532 55456 10538
rect 55404 10474 55456 10480
rect 55416 10441 55444 10474
rect 55692 10470 55720 10542
rect 55496 10464 55548 10470
rect 55402 10432 55458 10441
rect 55496 10406 55548 10412
rect 55680 10464 55732 10470
rect 55680 10406 55732 10412
rect 55402 10367 55458 10376
rect 55508 10266 55536 10406
rect 55496 10260 55548 10266
rect 55496 10202 55548 10208
rect 55312 10124 55364 10130
rect 55312 10066 55364 10072
rect 55220 8968 55272 8974
rect 55220 8910 55272 8916
rect 55324 6322 55352 10066
rect 55404 9988 55456 9994
rect 55404 9930 55456 9936
rect 55416 9178 55444 9930
rect 55692 9722 55720 10406
rect 55820 10364 56128 10373
rect 55820 10362 55826 10364
rect 55882 10362 55906 10364
rect 55962 10362 55986 10364
rect 56042 10362 56066 10364
rect 56122 10362 56128 10364
rect 55882 10310 55884 10362
rect 56064 10310 56066 10362
rect 55820 10308 55826 10310
rect 55882 10308 55906 10310
rect 55962 10308 55986 10310
rect 56042 10308 56066 10310
rect 56122 10308 56128 10310
rect 55820 10299 56128 10308
rect 56244 9926 56272 10934
rect 56336 10742 56364 15030
rect 56520 15008 56548 15438
rect 56784 15428 56836 15434
rect 56784 15370 56836 15376
rect 56692 15020 56744 15026
rect 56520 14980 56692 15008
rect 56692 14962 56744 14968
rect 56416 14544 56468 14550
rect 56416 14486 56468 14492
rect 56428 12850 56456 14486
rect 56508 14476 56560 14482
rect 56508 14418 56560 14424
rect 56416 12844 56468 12850
rect 56416 12786 56468 12792
rect 56520 11898 56548 14418
rect 56796 14346 56824 15370
rect 56874 15192 56930 15201
rect 56874 15127 56930 15136
rect 56888 15026 56916 15127
rect 56876 15020 56928 15026
rect 56876 14962 56928 14968
rect 56888 14793 56916 14962
rect 56980 14958 57008 18702
rect 56968 14952 57020 14958
rect 56966 14920 56968 14929
rect 57020 14920 57022 14929
rect 56966 14855 57022 14864
rect 56874 14784 56930 14793
rect 56874 14719 56930 14728
rect 57072 14634 57100 21082
rect 57152 20052 57204 20058
rect 57152 19994 57204 20000
rect 57164 19378 57192 19994
rect 57152 19372 57204 19378
rect 57152 19314 57204 19320
rect 57164 19174 57192 19314
rect 57152 19168 57204 19174
rect 57152 19110 57204 19116
rect 57704 18896 57756 18902
rect 57704 18838 57756 18844
rect 57716 17202 57744 18838
rect 57980 18148 58032 18154
rect 57980 18090 58032 18096
rect 57886 17504 57942 17513
rect 57992 17490 58020 18090
rect 57942 17462 58020 17490
rect 57886 17439 57942 17448
rect 57992 17326 58204 17354
rect 57704 17196 57756 17202
rect 57704 17138 57756 17144
rect 57888 17196 57940 17202
rect 57888 17138 57940 17144
rect 57426 16688 57482 16697
rect 57426 16623 57482 16632
rect 57336 16448 57388 16454
rect 57336 16390 57388 16396
rect 57244 15700 57296 15706
rect 57244 15642 57296 15648
rect 57072 14606 57192 14634
rect 56600 14340 56652 14346
rect 56600 14282 56652 14288
rect 56784 14340 56836 14346
rect 56784 14282 56836 14288
rect 56968 14340 57020 14346
rect 56968 14282 57020 14288
rect 56612 12617 56640 14282
rect 56796 13938 56824 14282
rect 56784 13932 56836 13938
rect 56784 13874 56836 13880
rect 56876 13932 56928 13938
rect 56876 13874 56928 13880
rect 56888 13841 56916 13874
rect 56980 13870 57008 14282
rect 57058 14104 57114 14113
rect 57058 14039 57114 14048
rect 56968 13864 57020 13870
rect 56874 13832 56930 13841
rect 56968 13806 57020 13812
rect 56874 13767 56930 13776
rect 56980 13326 57008 13806
rect 57072 13569 57100 14039
rect 57058 13560 57114 13569
rect 57058 13495 57114 13504
rect 57164 13444 57192 14606
rect 57256 14278 57284 15642
rect 57348 15366 57376 16390
rect 57440 15366 57468 16623
rect 57518 16552 57574 16561
rect 57518 16487 57574 16496
rect 57532 15502 57560 16487
rect 57520 15496 57572 15502
rect 57520 15438 57572 15444
rect 57336 15360 57388 15366
rect 57336 15302 57388 15308
rect 57428 15360 57480 15366
rect 57428 15302 57480 15308
rect 57610 14512 57666 14521
rect 57610 14447 57666 14456
rect 57244 14272 57296 14278
rect 57296 14232 57376 14260
rect 57244 14214 57296 14220
rect 57242 14104 57298 14113
rect 57242 14039 57298 14048
rect 57256 13938 57284 14039
rect 57244 13932 57296 13938
rect 57244 13874 57296 13880
rect 57072 13416 57192 13444
rect 56968 13320 57020 13326
rect 56968 13262 57020 13268
rect 57072 13138 57100 13416
rect 56888 13110 57100 13138
rect 56692 12844 56744 12850
rect 56692 12786 56744 12792
rect 56784 12844 56836 12850
rect 56784 12786 56836 12792
rect 56598 12608 56654 12617
rect 56598 12543 56654 12552
rect 56600 12368 56652 12374
rect 56600 12310 56652 12316
rect 56612 12102 56640 12310
rect 56600 12096 56652 12102
rect 56600 12038 56652 12044
rect 56508 11892 56560 11898
rect 56508 11834 56560 11840
rect 56508 11688 56560 11694
rect 56508 11630 56560 11636
rect 56414 11520 56470 11529
rect 56414 11455 56470 11464
rect 56324 10736 56376 10742
rect 56324 10678 56376 10684
rect 56232 9920 56284 9926
rect 56232 9862 56284 9868
rect 55680 9716 55732 9722
rect 55680 9658 55732 9664
rect 55820 9276 56128 9285
rect 55820 9274 55826 9276
rect 55882 9274 55906 9276
rect 55962 9274 55986 9276
rect 56042 9274 56066 9276
rect 56122 9274 56128 9276
rect 55882 9222 55884 9274
rect 56064 9222 56066 9274
rect 55820 9220 55826 9222
rect 55882 9220 55906 9222
rect 55962 9220 55986 9222
rect 56042 9220 56066 9222
rect 56122 9220 56128 9222
rect 55820 9211 56128 9220
rect 55404 9172 55456 9178
rect 55404 9114 55456 9120
rect 55588 8492 55640 8498
rect 55588 8434 55640 8440
rect 55312 6316 55364 6322
rect 55312 6258 55364 6264
rect 54944 2984 54996 2990
rect 54944 2926 54996 2932
rect 54392 2848 54444 2854
rect 54392 2790 54444 2796
rect 53024 2746 53328 2774
rect 53300 2650 53328 2746
rect 53288 2644 53340 2650
rect 53288 2586 53340 2592
rect 54404 2446 54432 2790
rect 55600 2650 55628 8434
rect 55820 8188 56128 8197
rect 55820 8186 55826 8188
rect 55882 8186 55906 8188
rect 55962 8186 55986 8188
rect 56042 8186 56066 8188
rect 56122 8186 56128 8188
rect 55882 8134 55884 8186
rect 56064 8134 56066 8186
rect 55820 8132 55826 8134
rect 55882 8132 55906 8134
rect 55962 8132 55986 8134
rect 56042 8132 56066 8134
rect 56122 8132 56128 8134
rect 55820 8123 56128 8132
rect 55820 7100 56128 7109
rect 55820 7098 55826 7100
rect 55882 7098 55906 7100
rect 55962 7098 55986 7100
rect 56042 7098 56066 7100
rect 56122 7098 56128 7100
rect 55882 7046 55884 7098
rect 56064 7046 56066 7098
rect 55820 7044 55826 7046
rect 55882 7044 55906 7046
rect 55962 7044 55986 7046
rect 56042 7044 56066 7046
rect 56122 7044 56128 7046
rect 55820 7035 56128 7044
rect 56048 6656 56100 6662
rect 56048 6598 56100 6604
rect 56060 6322 56088 6598
rect 56048 6316 56100 6322
rect 56048 6258 56100 6264
rect 55820 6012 56128 6021
rect 55820 6010 55826 6012
rect 55882 6010 55906 6012
rect 55962 6010 55986 6012
rect 56042 6010 56066 6012
rect 56122 6010 56128 6012
rect 55882 5958 55884 6010
rect 56064 5958 56066 6010
rect 55820 5956 55826 5958
rect 55882 5956 55906 5958
rect 55962 5956 55986 5958
rect 56042 5956 56066 5958
rect 56122 5956 56128 5958
rect 55820 5947 56128 5956
rect 55820 4924 56128 4933
rect 55820 4922 55826 4924
rect 55882 4922 55906 4924
rect 55962 4922 55986 4924
rect 56042 4922 56066 4924
rect 56122 4922 56128 4924
rect 55882 4870 55884 4922
rect 56064 4870 56066 4922
rect 55820 4868 55826 4870
rect 55882 4868 55906 4870
rect 55962 4868 55986 4870
rect 56042 4868 56066 4870
rect 56122 4868 56128 4870
rect 55820 4859 56128 4868
rect 55680 4480 55732 4486
rect 55680 4422 55732 4428
rect 55692 3058 55720 4422
rect 55820 3836 56128 3845
rect 55820 3834 55826 3836
rect 55882 3834 55906 3836
rect 55962 3834 55986 3836
rect 56042 3834 56066 3836
rect 56122 3834 56128 3836
rect 55882 3782 55884 3834
rect 56064 3782 56066 3834
rect 55820 3780 55826 3782
rect 55882 3780 55906 3782
rect 55962 3780 55986 3782
rect 56042 3780 56066 3782
rect 56122 3780 56128 3782
rect 55820 3771 56128 3780
rect 55680 3052 55732 3058
rect 55680 2994 55732 3000
rect 56428 2774 56456 11455
rect 56520 10742 56548 11630
rect 56600 11552 56652 11558
rect 56598 11520 56600 11529
rect 56652 11520 56654 11529
rect 56598 11455 56654 11464
rect 56704 11082 56732 12786
rect 56796 12306 56824 12786
rect 56888 12764 56916 13110
rect 57060 12980 57112 12986
rect 57060 12922 57112 12928
rect 56968 12776 57020 12782
rect 56888 12736 56968 12764
rect 56968 12718 57020 12724
rect 57072 12730 57100 12922
rect 57256 12900 57284 13874
rect 57348 13870 57376 14232
rect 57336 13864 57388 13870
rect 57336 13806 57388 13812
rect 57426 13696 57482 13705
rect 57426 13631 57482 13640
rect 57256 12872 57376 12900
rect 57348 12782 57376 12872
rect 57336 12776 57388 12782
rect 56784 12300 56836 12306
rect 56784 12242 56836 12248
rect 56980 11914 57008 12718
rect 57072 12702 57192 12730
rect 57336 12718 57388 12724
rect 57164 12442 57192 12702
rect 57060 12436 57112 12442
rect 57060 12378 57112 12384
rect 57152 12436 57204 12442
rect 57152 12378 57204 12384
rect 57072 12238 57100 12378
rect 57060 12232 57112 12238
rect 57060 12174 57112 12180
rect 56980 11886 57100 11914
rect 57072 11830 57100 11886
rect 56968 11824 57020 11830
rect 56968 11766 57020 11772
rect 57060 11824 57112 11830
rect 57060 11766 57112 11772
rect 56692 11076 56744 11082
rect 56692 11018 56744 11024
rect 56508 10736 56560 10742
rect 56980 10713 57008 11766
rect 57152 11756 57204 11762
rect 57152 11698 57204 11704
rect 57164 11626 57192 11698
rect 57152 11620 57204 11626
rect 57152 11562 57204 11568
rect 57060 11076 57112 11082
rect 57060 11018 57112 11024
rect 56508 10678 56560 10684
rect 56966 10704 57022 10713
rect 56600 10668 56652 10674
rect 56966 10639 57022 10648
rect 56600 10610 56652 10616
rect 56612 10470 56640 10610
rect 56600 10464 56652 10470
rect 56600 10406 56652 10412
rect 57072 9450 57100 11018
rect 57440 10826 57468 13631
rect 57520 13184 57572 13190
rect 57520 13126 57572 13132
rect 57532 12986 57560 13126
rect 57624 12986 57652 14447
rect 57520 12980 57572 12986
rect 57520 12922 57572 12928
rect 57612 12980 57664 12986
rect 57612 12922 57664 12928
rect 57624 12850 57652 12922
rect 57520 12844 57572 12850
rect 57520 12786 57572 12792
rect 57612 12844 57664 12850
rect 57612 12786 57664 12792
rect 57532 12442 57560 12786
rect 57520 12436 57572 12442
rect 57520 12378 57572 12384
rect 57612 12232 57664 12238
rect 57612 12174 57664 12180
rect 57520 11824 57572 11830
rect 57520 11766 57572 11772
rect 57532 11529 57560 11766
rect 57518 11520 57574 11529
rect 57518 11455 57574 11464
rect 57164 10798 57468 10826
rect 57060 9444 57112 9450
rect 57060 9386 57112 9392
rect 56968 6792 57020 6798
rect 56968 6734 57020 6740
rect 56980 5914 57008 6734
rect 56968 5908 57020 5914
rect 56968 5850 57020 5856
rect 56600 2848 56652 2854
rect 56600 2790 56652 2796
rect 55820 2748 56128 2757
rect 55820 2746 55826 2748
rect 55882 2746 55906 2748
rect 55962 2746 55986 2748
rect 56042 2746 56066 2748
rect 56122 2746 56128 2748
rect 56428 2746 56548 2774
rect 55882 2694 55884 2746
rect 56064 2694 56066 2746
rect 55820 2692 55826 2694
rect 55882 2692 55906 2694
rect 55962 2692 55986 2694
rect 56042 2692 56066 2694
rect 56122 2692 56128 2694
rect 55820 2683 56128 2692
rect 55588 2644 55640 2650
rect 55588 2586 55640 2592
rect 54392 2440 54444 2446
rect 54392 2382 54444 2388
rect 54760 2440 54812 2446
rect 56520 2417 56548 2746
rect 56612 2446 56640 2790
rect 57164 2446 57192 10798
rect 57428 10668 57480 10674
rect 57428 10610 57480 10616
rect 57440 10266 57468 10610
rect 57428 10260 57480 10266
rect 57428 10202 57480 10208
rect 57624 10169 57652 12174
rect 57610 10160 57666 10169
rect 57610 10095 57666 10104
rect 57244 9920 57296 9926
rect 57244 9862 57296 9868
rect 57256 9586 57284 9862
rect 57244 9580 57296 9586
rect 57244 9522 57296 9528
rect 57336 6452 57388 6458
rect 57336 6394 57388 6400
rect 57348 5710 57376 6394
rect 57716 5778 57744 17138
rect 57900 16522 57928 17138
rect 57888 16516 57940 16522
rect 57888 16458 57940 16464
rect 57900 16114 57928 16458
rect 57992 16153 58020 17326
rect 58176 17202 58204 17326
rect 58544 17270 58572 25706
rect 58636 17785 58664 27338
rect 58716 27328 58768 27334
rect 58716 27270 58768 27276
rect 59268 27328 59320 27334
rect 59268 27270 59320 27276
rect 58728 18154 58756 27270
rect 58992 26988 59044 26994
rect 58992 26930 59044 26936
rect 59004 26450 59032 26930
rect 58992 26444 59044 26450
rect 58992 26386 59044 26392
rect 59280 21457 59308 27270
rect 59648 26790 59676 27406
rect 60004 27396 60056 27402
rect 60004 27338 60056 27344
rect 59636 26784 59688 26790
rect 59636 26726 59688 26732
rect 59266 21448 59322 21457
rect 59266 21383 59322 21392
rect 59268 20052 59320 20058
rect 59268 19994 59320 20000
rect 59176 18692 59228 18698
rect 59176 18634 59228 18640
rect 58716 18148 58768 18154
rect 58716 18090 58768 18096
rect 58622 17776 58678 17785
rect 58622 17711 58678 17720
rect 58716 17672 58768 17678
rect 58716 17614 58768 17620
rect 58992 17672 59044 17678
rect 58992 17614 59044 17620
rect 58532 17264 58584 17270
rect 58532 17206 58584 17212
rect 58622 17232 58678 17241
rect 58072 17196 58124 17202
rect 58072 17138 58124 17144
rect 58164 17196 58216 17202
rect 58622 17167 58678 17176
rect 58164 17138 58216 17144
rect 57978 16144 58034 16153
rect 57888 16108 57940 16114
rect 58084 16130 58112 17138
rect 58636 17134 58664 17167
rect 58624 17128 58676 17134
rect 58624 17070 58676 17076
rect 58728 16726 58756 17614
rect 58808 17196 58860 17202
rect 58808 17138 58860 17144
rect 58900 17196 58952 17202
rect 58900 17138 58952 17144
rect 58820 17105 58848 17138
rect 58806 17096 58862 17105
rect 58806 17031 58862 17040
rect 58912 16833 58940 17138
rect 58898 16824 58954 16833
rect 58820 16782 58898 16810
rect 58716 16720 58768 16726
rect 58716 16662 58768 16668
rect 58440 16516 58492 16522
rect 58440 16458 58492 16464
rect 58452 16182 58480 16458
rect 58532 16448 58584 16454
rect 58532 16390 58584 16396
rect 58440 16176 58492 16182
rect 58254 16144 58310 16153
rect 58084 16102 58254 16130
rect 58440 16118 58492 16124
rect 58544 16114 58572 16390
rect 58622 16280 58678 16289
rect 58622 16215 58678 16224
rect 58636 16182 58664 16215
rect 58624 16176 58676 16182
rect 58624 16118 58676 16124
rect 57978 16079 58034 16088
rect 58254 16079 58256 16088
rect 57888 16050 57940 16056
rect 58308 16079 58310 16088
rect 58348 16108 58400 16114
rect 58256 16050 58308 16056
rect 58348 16050 58400 16056
rect 58532 16108 58584 16114
rect 58532 16050 58584 16056
rect 57794 14376 57850 14385
rect 57794 14311 57796 14320
rect 57848 14311 57850 14320
rect 57796 14282 57848 14288
rect 57900 13954 57928 16050
rect 57980 16040 58032 16046
rect 57978 16008 57980 16017
rect 58032 16008 58034 16017
rect 58034 15966 58112 15994
rect 57978 15943 58034 15952
rect 57980 15428 58032 15434
rect 57980 15370 58032 15376
rect 57992 14890 58020 15370
rect 58084 14958 58112 15966
rect 58164 15972 58216 15978
rect 58164 15914 58216 15920
rect 58176 15570 58204 15914
rect 58268 15706 58296 16050
rect 58256 15700 58308 15706
rect 58256 15642 58308 15648
rect 58360 15638 58388 16050
rect 58636 15994 58664 16118
rect 58452 15966 58664 15994
rect 58348 15632 58400 15638
rect 58348 15574 58400 15580
rect 58164 15564 58216 15570
rect 58164 15506 58216 15512
rect 58256 15564 58308 15570
rect 58256 15506 58308 15512
rect 58268 15094 58296 15506
rect 58164 15088 58216 15094
rect 58164 15030 58216 15036
rect 58256 15088 58308 15094
rect 58256 15030 58308 15036
rect 58072 14952 58124 14958
rect 58176 14940 58204 15030
rect 58176 14912 58296 14940
rect 58072 14894 58124 14900
rect 57980 14884 58032 14890
rect 57980 14826 58032 14832
rect 57978 14648 58034 14657
rect 57978 14583 58034 14592
rect 57992 14414 58020 14583
rect 58164 14476 58216 14482
rect 58164 14418 58216 14424
rect 57980 14408 58032 14414
rect 57980 14350 58032 14356
rect 58072 14408 58124 14414
rect 58072 14350 58124 14356
rect 58084 14090 58112 14350
rect 58176 14346 58204 14418
rect 58164 14340 58216 14346
rect 58164 14282 58216 14288
rect 58084 14062 58204 14090
rect 57900 13938 58020 13954
rect 57888 13932 58020 13938
rect 57940 13926 58020 13932
rect 57888 13874 57940 13880
rect 57888 13320 57940 13326
rect 57888 13262 57940 13268
rect 57900 12434 57928 13262
rect 57992 12850 58020 13926
rect 58176 13326 58204 14062
rect 58164 13320 58216 13326
rect 58070 13288 58126 13297
rect 58164 13262 58216 13268
rect 58070 13223 58126 13232
rect 57980 12844 58032 12850
rect 57980 12786 58032 12792
rect 58084 12782 58112 13223
rect 58176 13025 58204 13262
rect 58162 13016 58218 13025
rect 58162 12951 58218 12960
rect 58072 12776 58124 12782
rect 58072 12718 58124 12724
rect 58084 12434 58112 12718
rect 57808 12406 58020 12434
rect 58084 12406 58204 12434
rect 57808 12374 57836 12406
rect 57796 12368 57848 12374
rect 57796 12310 57848 12316
rect 57888 12368 57940 12374
rect 57888 12310 57940 12316
rect 57796 12232 57848 12238
rect 57796 12174 57848 12180
rect 57808 12102 57836 12174
rect 57796 12096 57848 12102
rect 57796 12038 57848 12044
rect 57900 11762 57928 12310
rect 57992 12238 58020 12406
rect 57980 12232 58032 12238
rect 57980 12174 58032 12180
rect 57888 11756 57940 11762
rect 57888 11698 57940 11704
rect 58072 11620 58124 11626
rect 58072 11562 58124 11568
rect 57796 11280 57848 11286
rect 58084 11257 58112 11562
rect 57796 11222 57848 11228
rect 58070 11248 58126 11257
rect 57808 10470 57836 11222
rect 58070 11183 58126 11192
rect 58072 11076 58124 11082
rect 58072 11018 58124 11024
rect 58084 10538 58112 11018
rect 58072 10532 58124 10538
rect 58072 10474 58124 10480
rect 57796 10464 57848 10470
rect 57796 10406 57848 10412
rect 57808 10062 57836 10406
rect 57796 10056 57848 10062
rect 57796 9998 57848 10004
rect 58176 9994 58204 12406
rect 58164 9988 58216 9994
rect 58164 9930 58216 9936
rect 57704 5772 57756 5778
rect 57704 5714 57756 5720
rect 57336 5704 57388 5710
rect 57336 5646 57388 5652
rect 57348 4622 57376 5646
rect 57336 4616 57388 4622
rect 57336 4558 57388 4564
rect 58268 2774 58296 14912
rect 58348 14816 58400 14822
rect 58348 14758 58400 14764
rect 58360 14550 58388 14758
rect 58348 14544 58400 14550
rect 58348 14486 58400 14492
rect 58452 14482 58480 15966
rect 58716 15904 58768 15910
rect 58716 15846 58768 15852
rect 58622 15600 58678 15609
rect 58622 15535 58624 15544
rect 58676 15535 58678 15544
rect 58624 15506 58676 15512
rect 58530 14512 58586 14521
rect 58440 14476 58492 14482
rect 58636 14482 58664 15506
rect 58728 15502 58756 15846
rect 58716 15496 58768 15502
rect 58716 15438 58768 15444
rect 58716 14952 58768 14958
rect 58716 14894 58768 14900
rect 58530 14447 58586 14456
rect 58624 14476 58676 14482
rect 58440 14418 58492 14424
rect 58348 13932 58400 13938
rect 58348 13874 58400 13880
rect 58360 13530 58388 13874
rect 58544 13870 58572 14447
rect 58624 14418 58676 14424
rect 58532 13864 58584 13870
rect 58532 13806 58584 13812
rect 58348 13524 58400 13530
rect 58348 13466 58400 13472
rect 58348 13320 58400 13326
rect 58346 13288 58348 13297
rect 58400 13288 58402 13297
rect 58346 13223 58402 13232
rect 58346 13016 58402 13025
rect 58346 12951 58402 12960
rect 58360 12170 58388 12951
rect 58636 12186 58664 14418
rect 58728 12850 58756 14894
rect 58716 12844 58768 12850
rect 58716 12786 58768 12792
rect 58714 12472 58770 12481
rect 58714 12407 58770 12416
rect 58348 12164 58400 12170
rect 58348 12106 58400 12112
rect 58452 12158 58664 12186
rect 58348 11756 58400 11762
rect 58348 11698 58400 11704
rect 58360 11529 58388 11698
rect 58346 11520 58402 11529
rect 58346 11455 58402 11464
rect 58360 3602 58388 11455
rect 58452 11150 58480 12158
rect 58624 12096 58676 12102
rect 58728 12084 58756 12407
rect 58676 12056 58756 12084
rect 58624 12038 58676 12044
rect 58532 11688 58584 11694
rect 58532 11630 58584 11636
rect 58440 11144 58492 11150
rect 58440 11086 58492 11092
rect 58544 10742 58572 11630
rect 58820 11257 58848 16782
rect 58898 16759 58954 16768
rect 58900 16652 58952 16658
rect 58900 16594 58952 16600
rect 58912 16561 58940 16594
rect 58898 16552 58954 16561
rect 58898 16487 58954 16496
rect 59004 16114 59032 17614
rect 59084 17536 59136 17542
rect 59082 17504 59084 17513
rect 59136 17504 59138 17513
rect 59082 17439 59138 17448
rect 59084 16516 59136 16522
rect 59084 16458 59136 16464
rect 58992 16108 59044 16114
rect 58992 16050 59044 16056
rect 58992 15904 59044 15910
rect 58992 15846 59044 15852
rect 59004 15706 59032 15846
rect 58992 15700 59044 15706
rect 58992 15642 59044 15648
rect 58900 13184 58952 13190
rect 58900 13126 58952 13132
rect 58912 11830 58940 13126
rect 58900 11824 58952 11830
rect 58900 11766 58952 11772
rect 58900 11552 58952 11558
rect 58900 11494 58952 11500
rect 58806 11248 58862 11257
rect 58806 11183 58862 11192
rect 58532 10736 58584 10742
rect 58532 10678 58584 10684
rect 58716 10668 58768 10674
rect 58820 10656 58848 11183
rect 58912 11082 58940 11494
rect 58900 11076 58952 11082
rect 58900 11018 58952 11024
rect 58768 10628 58848 10656
rect 58900 10668 58952 10674
rect 58716 10610 58768 10616
rect 58900 10610 58952 10616
rect 58912 10470 58940 10610
rect 58440 10464 58492 10470
rect 58440 10406 58492 10412
rect 58900 10464 58952 10470
rect 58900 10406 58952 10412
rect 58452 7818 58480 10406
rect 58624 9920 58676 9926
rect 58624 9862 58676 9868
rect 58440 7812 58492 7818
rect 58440 7754 58492 7760
rect 58636 3602 58664 9862
rect 58348 3596 58400 3602
rect 58348 3538 58400 3544
rect 58624 3596 58676 3602
rect 58624 3538 58676 3544
rect 58636 3058 58664 3538
rect 58624 3052 58676 3058
rect 58624 2994 58676 3000
rect 58348 2848 58400 2854
rect 58348 2790 58400 2796
rect 57992 2746 58296 2774
rect 57992 2446 58020 2746
rect 58360 2446 58388 2790
rect 56600 2440 56652 2446
rect 54760 2382 54812 2388
rect 56506 2408 56562 2417
rect 53196 2304 53248 2310
rect 53196 2246 53248 2252
rect 54116 2304 54168 2310
rect 54116 2246 54168 2252
rect 52920 2032 52972 2038
rect 52920 1974 52972 1980
rect 53208 1902 53236 2246
rect 53196 1896 53248 1902
rect 53196 1838 53248 1844
rect 54128 800 54156 2246
rect 54772 800 54800 2382
rect 55404 2372 55456 2378
rect 56600 2382 56652 2388
rect 57152 2440 57204 2446
rect 57152 2382 57204 2388
rect 57980 2440 58032 2446
rect 57980 2382 58032 2388
rect 58348 2440 58400 2446
rect 58348 2382 58400 2388
rect 56506 2343 56562 2352
rect 55404 2314 55456 2320
rect 55416 800 55444 2314
rect 56048 2304 56100 2310
rect 56048 2246 56100 2252
rect 56692 2304 56744 2310
rect 56692 2246 56744 2252
rect 57336 2304 57388 2310
rect 57336 2246 57388 2252
rect 57980 2304 58032 2310
rect 57980 2246 58032 2252
rect 58624 2304 58676 2310
rect 58624 2246 58676 2252
rect 56060 800 56088 2246
rect 56704 800 56732 2246
rect 57348 800 57376 2246
rect 57992 800 58020 2246
rect 58636 800 58664 2246
rect 59004 1902 59032 15642
rect 59096 14346 59124 16458
rect 59188 16114 59216 18634
rect 59280 17678 59308 19994
rect 59268 17672 59320 17678
rect 59268 17614 59320 17620
rect 59912 17672 59964 17678
rect 59912 17614 59964 17620
rect 59360 17604 59412 17610
rect 59360 17546 59412 17552
rect 59372 17354 59400 17546
rect 59728 17536 59780 17542
rect 59728 17478 59780 17484
rect 59280 17326 59400 17354
rect 59280 17134 59308 17326
rect 59740 17202 59768 17478
rect 59924 17270 59952 17614
rect 59912 17264 59964 17270
rect 59912 17206 59964 17212
rect 59728 17196 59780 17202
rect 59728 17138 59780 17144
rect 60016 17134 60044 27338
rect 60568 27334 60596 27542
rect 60556 27328 60608 27334
rect 60556 27270 60608 27276
rect 60660 27130 60688 29294
rect 61198 29294 61332 29322
rect 61198 29200 61254 29294
rect 61304 27470 61332 29294
rect 61842 29294 61976 29322
rect 61842 29200 61898 29294
rect 61948 27606 61976 29294
rect 62486 29200 62542 30000
rect 63774 29322 63830 30000
rect 64418 29322 64474 30000
rect 63774 29294 63908 29322
rect 63774 29200 63830 29294
rect 62500 27606 62528 29200
rect 61936 27600 61988 27606
rect 61936 27542 61988 27548
rect 62488 27600 62540 27606
rect 62488 27542 62540 27548
rect 63880 27470 63908 29294
rect 64418 29294 64828 29322
rect 64418 29200 64474 29294
rect 64800 27554 64828 29294
rect 65062 29200 65118 30000
rect 65706 29200 65762 30000
rect 66350 29200 66406 30000
rect 66994 29200 67050 30000
rect 67638 29200 67694 30000
rect 68282 29322 68338 30000
rect 68282 29294 68692 29322
rect 68282 29200 68338 29294
rect 65076 27606 65104 29200
rect 65720 27606 65748 29200
rect 66364 27606 66392 29200
rect 65064 27600 65116 27606
rect 64800 27526 64920 27554
rect 65064 27542 65116 27548
rect 65708 27600 65760 27606
rect 65708 27542 65760 27548
rect 66352 27600 66404 27606
rect 66352 27542 66404 27548
rect 61292 27464 61344 27470
rect 61292 27406 61344 27412
rect 61384 27464 61436 27470
rect 61384 27406 61436 27412
rect 63868 27464 63920 27470
rect 63868 27406 63920 27412
rect 64420 27464 64472 27470
rect 64420 27406 64472 27412
rect 60648 27124 60700 27130
rect 60648 27066 60700 27072
rect 61396 18222 61424 27406
rect 61568 27396 61620 27402
rect 61568 27338 61620 27344
rect 61580 22094 61608 27338
rect 63408 24268 63460 24274
rect 63408 24210 63460 24216
rect 61488 22066 61608 22094
rect 60372 18216 60424 18222
rect 60372 18158 60424 18164
rect 60556 18216 60608 18222
rect 60556 18158 60608 18164
rect 61384 18216 61436 18222
rect 61384 18158 61436 18164
rect 60384 17626 60412 18158
rect 60568 17882 60596 18158
rect 60556 17876 60608 17882
rect 60556 17818 60608 17824
rect 60464 17808 60516 17814
rect 60462 17776 60464 17785
rect 60648 17808 60700 17814
rect 60516 17776 60518 17785
rect 61016 17808 61068 17814
rect 60648 17750 60700 17756
rect 60830 17776 60886 17785
rect 60462 17711 60518 17720
rect 60384 17598 60596 17626
rect 60660 17610 60688 17750
rect 61016 17750 61068 17756
rect 61108 17808 61160 17814
rect 61108 17750 61160 17756
rect 60830 17711 60832 17720
rect 60884 17711 60886 17720
rect 60832 17682 60884 17688
rect 60372 17536 60424 17542
rect 60372 17478 60424 17484
rect 60278 17368 60334 17377
rect 60278 17303 60334 17312
rect 59268 17128 59320 17134
rect 59268 17070 59320 17076
rect 59544 17128 59596 17134
rect 59544 17070 59596 17076
rect 59820 17128 59872 17134
rect 59820 17070 59872 17076
rect 60004 17128 60056 17134
rect 60004 17070 60056 17076
rect 59268 16992 59320 16998
rect 59268 16934 59320 16940
rect 59280 16726 59308 16934
rect 59268 16720 59320 16726
rect 59556 16697 59584 17070
rect 59542 16688 59598 16697
rect 59268 16662 59320 16668
rect 59372 16646 59542 16674
rect 59268 16516 59320 16522
rect 59268 16458 59320 16464
rect 59176 16108 59228 16114
rect 59176 16050 59228 16056
rect 59280 16017 59308 16458
rect 59266 16008 59322 16017
rect 59266 15943 59322 15952
rect 59372 15094 59400 16646
rect 59542 16623 59598 16632
rect 59360 15088 59412 15094
rect 59412 15036 59492 15042
rect 59360 15030 59492 15036
rect 59372 15014 59492 15030
rect 59360 14952 59412 14958
rect 59360 14894 59412 14900
rect 59372 14770 59400 14894
rect 59280 14742 59400 14770
rect 59084 14340 59136 14346
rect 59084 14282 59136 14288
rect 59280 13870 59308 14742
rect 59464 13938 59492 15014
rect 59544 15020 59596 15026
rect 59544 14962 59596 14968
rect 59556 14498 59584 14962
rect 59636 14544 59688 14550
rect 59556 14492 59636 14498
rect 59556 14486 59688 14492
rect 59556 14470 59676 14486
rect 59452 13932 59504 13938
rect 59452 13874 59504 13880
rect 59176 13864 59228 13870
rect 59176 13806 59228 13812
rect 59268 13864 59320 13870
rect 59268 13806 59320 13812
rect 59188 12986 59216 13806
rect 59280 13258 59308 13806
rect 59452 13456 59504 13462
rect 59452 13398 59504 13404
rect 59360 13320 59412 13326
rect 59464 13297 59492 13398
rect 59360 13262 59412 13268
rect 59450 13288 59506 13297
rect 59268 13252 59320 13258
rect 59268 13194 59320 13200
rect 59372 13002 59400 13262
rect 59450 13223 59506 13232
rect 59372 12986 59492 13002
rect 59084 12980 59136 12986
rect 59084 12922 59136 12928
rect 59176 12980 59228 12986
rect 59372 12980 59504 12986
rect 59372 12974 59452 12980
rect 59176 12922 59228 12928
rect 59452 12922 59504 12928
rect 59096 12288 59124 12922
rect 59452 12776 59504 12782
rect 59452 12718 59504 12724
rect 59176 12300 59228 12306
rect 59096 12260 59176 12288
rect 59176 12242 59228 12248
rect 59176 12164 59228 12170
rect 59176 12106 59228 12112
rect 59188 11830 59216 12106
rect 59266 11928 59322 11937
rect 59266 11863 59322 11872
rect 59176 11824 59228 11830
rect 59176 11766 59228 11772
rect 59084 11756 59136 11762
rect 59084 11698 59136 11704
rect 59096 10674 59124 11698
rect 59280 11558 59308 11863
rect 59360 11756 59412 11762
rect 59464 11744 59492 12718
rect 59412 11716 59492 11744
rect 59360 11698 59412 11704
rect 59176 11552 59228 11558
rect 59176 11494 59228 11500
rect 59268 11552 59320 11558
rect 59268 11494 59320 11500
rect 59084 10668 59136 10674
rect 59084 10610 59136 10616
rect 59188 10538 59216 11494
rect 59372 10985 59400 11698
rect 59452 11144 59504 11150
rect 59452 11086 59504 11092
rect 59358 10976 59414 10985
rect 59358 10911 59414 10920
rect 59176 10532 59228 10538
rect 59176 10474 59228 10480
rect 59188 10062 59216 10474
rect 59176 10056 59228 10062
rect 59176 9998 59228 10004
rect 59268 9716 59320 9722
rect 59268 9658 59320 9664
rect 59176 2848 59228 2854
rect 59176 2790 59228 2796
rect 59188 2446 59216 2790
rect 59280 2650 59308 9658
rect 59464 9586 59492 11086
rect 59452 9580 59504 9586
rect 59452 9522 59504 9528
rect 59452 4548 59504 4554
rect 59452 4490 59504 4496
rect 59464 4214 59492 4490
rect 59452 4208 59504 4214
rect 59452 4150 59504 4156
rect 59556 2774 59584 14470
rect 59832 13326 59860 17070
rect 60292 17066 60320 17303
rect 60384 17202 60412 17478
rect 60372 17196 60424 17202
rect 60372 17138 60424 17144
rect 60280 17060 60332 17066
rect 60280 17002 60332 17008
rect 59912 16652 59964 16658
rect 59912 16594 59964 16600
rect 59924 15201 59952 16594
rect 60096 16516 60148 16522
rect 60096 16458 60148 16464
rect 60004 16108 60056 16114
rect 60004 16050 60056 16056
rect 60016 15706 60044 16050
rect 60004 15700 60056 15706
rect 60004 15642 60056 15648
rect 59910 15192 59966 15201
rect 59910 15127 59966 15136
rect 59924 14482 59952 15127
rect 60002 14784 60058 14793
rect 60002 14719 60058 14728
rect 59912 14476 59964 14482
rect 59912 14418 59964 14424
rect 60016 13841 60044 14719
rect 60002 13832 60058 13841
rect 60002 13767 60058 13776
rect 59820 13320 59872 13326
rect 59820 13262 59872 13268
rect 59636 13252 59688 13258
rect 59636 13194 59688 13200
rect 59648 12442 59676 13194
rect 59820 12912 59872 12918
rect 59820 12854 59872 12860
rect 59636 12436 59688 12442
rect 59636 12378 59688 12384
rect 59636 11076 59688 11082
rect 59636 11018 59688 11024
rect 59648 10577 59676 11018
rect 59832 10742 59860 12854
rect 60108 12646 60136 16458
rect 60188 16448 60240 16454
rect 60568 16436 60596 17598
rect 60648 17604 60700 17610
rect 60648 17546 60700 17552
rect 60832 17604 60884 17610
rect 60832 17546 60884 17552
rect 60646 17096 60702 17105
rect 60646 17031 60702 17040
rect 60660 16998 60688 17031
rect 60648 16992 60700 16998
rect 60648 16934 60700 16940
rect 60844 16590 60872 17546
rect 61028 17542 61056 17750
rect 60924 17536 60976 17542
rect 60924 17478 60976 17484
rect 61016 17536 61068 17542
rect 61016 17478 61068 17484
rect 60832 16584 60884 16590
rect 60832 16526 60884 16532
rect 60740 16516 60792 16522
rect 60740 16458 60792 16464
rect 60648 16448 60700 16454
rect 60568 16408 60648 16436
rect 60188 16390 60240 16396
rect 60752 16425 60780 16458
rect 60648 16390 60700 16396
rect 60738 16416 60794 16425
rect 60004 12640 60056 12646
rect 60004 12582 60056 12588
rect 60096 12640 60148 12646
rect 60096 12582 60148 12588
rect 59912 12436 59964 12442
rect 59912 12378 59964 12384
rect 59924 12345 59952 12378
rect 59910 12336 59966 12345
rect 59910 12271 59966 12280
rect 60016 12238 60044 12582
rect 60004 12232 60056 12238
rect 60004 12174 60056 12180
rect 60004 11756 60056 11762
rect 60004 11698 60056 11704
rect 60016 11354 60044 11698
rect 60004 11348 60056 11354
rect 60004 11290 60056 11296
rect 59820 10736 59872 10742
rect 59820 10678 59872 10684
rect 60200 10674 60228 16390
rect 60738 16351 60794 16360
rect 60740 16244 60792 16250
rect 60740 16186 60792 16192
rect 60464 16108 60516 16114
rect 60464 16050 60516 16056
rect 60280 16040 60332 16046
rect 60280 15982 60332 15988
rect 60372 16040 60424 16046
rect 60372 15982 60424 15988
rect 60292 15706 60320 15982
rect 60280 15700 60332 15706
rect 60280 15642 60332 15648
rect 60280 15564 60332 15570
rect 60280 15506 60332 15512
rect 60292 14249 60320 15506
rect 60384 15502 60412 15982
rect 60372 15496 60424 15502
rect 60372 15438 60424 15444
rect 60476 15314 60504 16050
rect 60752 15688 60780 16186
rect 60832 15700 60884 15706
rect 60752 15660 60832 15688
rect 60832 15642 60884 15648
rect 60936 15450 60964 17478
rect 61120 16590 61148 17750
rect 61384 17128 61436 17134
rect 61384 17070 61436 17076
rect 61396 16794 61424 17070
rect 61384 16788 61436 16794
rect 61384 16730 61436 16736
rect 61016 16584 61068 16590
rect 61016 16526 61068 16532
rect 61108 16584 61160 16590
rect 61108 16526 61160 16532
rect 61488 16538 61516 22066
rect 63224 21412 63276 21418
rect 63224 21354 63276 21360
rect 62764 18080 62816 18086
rect 62764 18022 62816 18028
rect 62776 17882 62804 18022
rect 62764 17876 62816 17882
rect 62132 17836 62344 17864
rect 61568 17672 61620 17678
rect 61568 17614 61620 17620
rect 61580 16794 61608 17614
rect 62132 17610 62160 17836
rect 62120 17604 62172 17610
rect 62120 17546 62172 17552
rect 62120 17196 62172 17202
rect 62120 17138 62172 17144
rect 61660 16992 61712 16998
rect 61660 16934 61712 16940
rect 61568 16788 61620 16794
rect 61568 16730 61620 16736
rect 61028 16402 61056 16526
rect 61200 16516 61252 16522
rect 61488 16510 61608 16538
rect 61672 16522 61700 16934
rect 62028 16720 62080 16726
rect 62028 16662 62080 16668
rect 61200 16458 61252 16464
rect 61212 16402 61240 16458
rect 61028 16374 61240 16402
rect 60844 15422 60964 15450
rect 60556 15360 60608 15366
rect 60384 15286 60504 15314
rect 60554 15328 60556 15337
rect 60608 15328 60610 15337
rect 60384 14346 60412 15286
rect 60554 15263 60610 15272
rect 60844 14958 60872 15422
rect 60924 15360 60976 15366
rect 60924 15302 60976 15308
rect 60832 14952 60884 14958
rect 60830 14920 60832 14929
rect 60884 14920 60886 14929
rect 60830 14855 60886 14864
rect 60844 14829 60872 14855
rect 60936 14414 60964 15302
rect 60464 14408 60516 14414
rect 60464 14350 60516 14356
rect 60924 14408 60976 14414
rect 60924 14350 60976 14356
rect 61292 14408 61344 14414
rect 61580 14396 61608 16510
rect 61660 16516 61712 16522
rect 61660 16458 61712 16464
rect 61842 15464 61898 15473
rect 61842 15399 61844 15408
rect 61896 15399 61898 15408
rect 61844 15370 61896 15376
rect 62040 15026 62068 16662
rect 62132 16114 62160 17138
rect 62316 17082 62344 17836
rect 62764 17818 62816 17824
rect 62764 17740 62816 17746
rect 62684 17700 62764 17728
rect 62396 17672 62448 17678
rect 62396 17614 62448 17620
rect 62488 17672 62540 17678
rect 62488 17614 62540 17620
rect 62408 17202 62436 17614
rect 62396 17196 62448 17202
rect 62396 17138 62448 17144
rect 62316 17054 62436 17082
rect 62408 16794 62436 17054
rect 62396 16788 62448 16794
rect 62396 16730 62448 16736
rect 62408 16114 62436 16730
rect 62120 16108 62172 16114
rect 62120 16050 62172 16056
rect 62396 16108 62448 16114
rect 62396 16050 62448 16056
rect 62212 16040 62264 16046
rect 62212 15982 62264 15988
rect 62224 15688 62252 15982
rect 62132 15660 62252 15688
rect 62132 15366 62160 15660
rect 62408 15638 62436 16050
rect 62396 15632 62448 15638
rect 62210 15600 62266 15609
rect 62396 15574 62448 15580
rect 62210 15535 62266 15544
rect 62120 15360 62172 15366
rect 62120 15302 62172 15308
rect 61752 15020 61804 15026
rect 61752 14962 61804 14968
rect 62028 15020 62080 15026
rect 62028 14962 62080 14968
rect 61764 14414 61792 14962
rect 61844 14952 61896 14958
rect 61844 14894 61896 14900
rect 61856 14550 61884 14894
rect 61844 14544 61896 14550
rect 61844 14486 61896 14492
rect 62028 14544 62080 14550
rect 62028 14486 62080 14492
rect 62118 14512 62174 14521
rect 62040 14414 62068 14486
rect 62118 14447 62120 14456
rect 62172 14447 62174 14456
rect 62120 14418 62172 14424
rect 61752 14408 61804 14414
rect 61580 14368 61700 14396
rect 61292 14350 61344 14356
rect 60372 14340 60424 14346
rect 60372 14282 60424 14288
rect 60278 14240 60334 14249
rect 60278 14175 60334 14184
rect 60292 14056 60320 14175
rect 60292 14028 60412 14056
rect 60278 13560 60334 13569
rect 60278 13495 60334 13504
rect 60292 13462 60320 13495
rect 60280 13456 60332 13462
rect 60280 13398 60332 13404
rect 60384 12481 60412 14028
rect 60476 12714 60504 14350
rect 60554 14240 60610 14249
rect 60554 14175 60610 14184
rect 60568 14074 60596 14175
rect 60556 14068 60608 14074
rect 60556 14010 60608 14016
rect 60648 13864 60700 13870
rect 60646 13832 60648 13841
rect 61016 13864 61068 13870
rect 60700 13832 60702 13841
rect 60646 13767 60702 13776
rect 60830 13832 60886 13841
rect 60830 13767 60886 13776
rect 61014 13832 61016 13841
rect 61068 13832 61070 13841
rect 61014 13767 61070 13776
rect 60554 13560 60610 13569
rect 60554 13495 60610 13504
rect 60568 13326 60596 13495
rect 60844 13462 60872 13767
rect 60740 13456 60792 13462
rect 60740 13398 60792 13404
rect 60832 13456 60884 13462
rect 60832 13398 60884 13404
rect 61108 13456 61160 13462
rect 61108 13398 61160 13404
rect 60556 13320 60608 13326
rect 60554 13288 60556 13297
rect 60752 13297 60780 13398
rect 60832 13320 60884 13326
rect 60608 13288 60610 13297
rect 60738 13288 60794 13297
rect 60554 13223 60610 13232
rect 60648 13252 60700 13258
rect 60832 13262 60884 13268
rect 61016 13320 61068 13326
rect 61016 13262 61068 13268
rect 60738 13223 60794 13232
rect 60648 13194 60700 13200
rect 60556 12912 60608 12918
rect 60556 12854 60608 12860
rect 60464 12708 60516 12714
rect 60464 12650 60516 12656
rect 60370 12472 60426 12481
rect 60370 12407 60426 12416
rect 60278 12336 60334 12345
rect 60278 12271 60334 12280
rect 60464 12300 60516 12306
rect 60292 11529 60320 12271
rect 60568 12288 60596 12854
rect 60660 12850 60688 13194
rect 60844 13161 60872 13262
rect 60830 13152 60886 13161
rect 60830 13087 60886 13096
rect 61028 12986 61056 13262
rect 61016 12980 61068 12986
rect 61016 12922 61068 12928
rect 60648 12844 60700 12850
rect 60648 12786 60700 12792
rect 60648 12708 60700 12714
rect 60648 12650 60700 12656
rect 60516 12260 60596 12288
rect 60464 12242 60516 12248
rect 60660 12186 60688 12650
rect 61016 12640 61068 12646
rect 61016 12582 61068 12588
rect 60384 12158 60688 12186
rect 60740 12164 60792 12170
rect 60384 12102 60412 12158
rect 60740 12106 60792 12112
rect 60372 12096 60424 12102
rect 60648 12096 60700 12102
rect 60372 12038 60424 12044
rect 60462 12064 60518 12073
rect 60646 12064 60648 12073
rect 60700 12064 60702 12073
rect 60518 12022 60596 12050
rect 60462 11999 60518 12008
rect 60568 11898 60596 12022
rect 60646 11999 60702 12008
rect 60556 11892 60608 11898
rect 60556 11834 60608 11840
rect 60568 11626 60688 11642
rect 60556 11620 60688 11626
rect 60608 11614 60688 11620
rect 60556 11562 60608 11568
rect 60278 11520 60334 11529
rect 60278 11455 60334 11464
rect 60554 11520 60610 11529
rect 60554 11455 60610 11464
rect 60568 11218 60596 11455
rect 60556 11212 60608 11218
rect 60556 11154 60608 11160
rect 60660 11150 60688 11614
rect 60752 11354 60780 12106
rect 60832 11688 60884 11694
rect 60832 11630 60884 11636
rect 60740 11348 60792 11354
rect 60740 11290 60792 11296
rect 60648 11144 60700 11150
rect 60648 11086 60700 11092
rect 60646 10976 60702 10985
rect 60646 10911 60702 10920
rect 60660 10742 60688 10911
rect 60844 10742 60872 11630
rect 61028 11064 61056 12582
rect 61120 12345 61148 13398
rect 61106 12336 61162 12345
rect 61106 12271 61162 12280
rect 61108 11892 61160 11898
rect 61108 11834 61160 11840
rect 61200 11892 61252 11898
rect 61200 11834 61252 11840
rect 61120 11801 61148 11834
rect 61106 11792 61162 11801
rect 61106 11727 61162 11736
rect 61212 11558 61240 11834
rect 61200 11552 61252 11558
rect 61200 11494 61252 11500
rect 61200 11076 61252 11082
rect 61028 11036 61200 11064
rect 61200 11018 61252 11024
rect 60648 10736 60700 10742
rect 60648 10678 60700 10684
rect 60832 10736 60884 10742
rect 60832 10678 60884 10684
rect 60188 10668 60240 10674
rect 60188 10610 60240 10616
rect 60740 10668 60792 10674
rect 60740 10610 60792 10616
rect 59634 10568 59690 10577
rect 59634 10503 59690 10512
rect 60752 10266 60780 10610
rect 60740 10260 60792 10266
rect 60740 10202 60792 10208
rect 60832 10056 60884 10062
rect 60832 9998 60884 10004
rect 59820 9920 59872 9926
rect 59820 9862 59872 9868
rect 59832 9654 59860 9862
rect 60844 9722 60872 9998
rect 60924 9920 60976 9926
rect 60924 9862 60976 9868
rect 60832 9716 60884 9722
rect 60832 9658 60884 9664
rect 59820 9648 59872 9654
rect 59820 9590 59872 9596
rect 60936 9110 60964 9862
rect 60924 9104 60976 9110
rect 60924 9046 60976 9052
rect 59636 3936 59688 3942
rect 59636 3878 59688 3884
rect 59648 3194 59676 3878
rect 59636 3188 59688 3194
rect 59636 3130 59688 3136
rect 59372 2746 59584 2774
rect 59268 2644 59320 2650
rect 59268 2586 59320 2592
rect 59176 2440 59228 2446
rect 59176 2382 59228 2388
rect 59268 2440 59320 2446
rect 59268 2382 59320 2388
rect 58992 1896 59044 1902
rect 58992 1838 59044 1844
rect 59280 800 59308 2382
rect 59372 1970 59400 2746
rect 61304 2650 61332 14350
rect 61384 14272 61436 14278
rect 61384 14214 61436 14220
rect 61396 13705 61424 14214
rect 61566 14104 61622 14113
rect 61566 14039 61568 14048
rect 61620 14039 61622 14048
rect 61568 14010 61620 14016
rect 61382 13696 61438 13705
rect 61382 13631 61438 13640
rect 61672 13530 61700 14368
rect 61752 14350 61804 14356
rect 62028 14408 62080 14414
rect 62028 14350 62080 14356
rect 61842 14104 61898 14113
rect 61842 14039 61898 14048
rect 61752 14000 61804 14006
rect 61752 13942 61804 13948
rect 61660 13524 61712 13530
rect 61660 13466 61712 13472
rect 61672 13326 61700 13466
rect 61660 13320 61712 13326
rect 61660 13262 61712 13268
rect 61476 11552 61528 11558
rect 61396 11512 61476 11540
rect 61396 11150 61424 11512
rect 61476 11494 61528 11500
rect 61764 11234 61792 13942
rect 61856 13938 61884 14039
rect 61844 13932 61896 13938
rect 61844 13874 61896 13880
rect 62028 13932 62080 13938
rect 62028 13874 62080 13880
rect 61844 12912 61896 12918
rect 61844 12854 61896 12860
rect 61856 12442 61884 12854
rect 61844 12436 61896 12442
rect 61844 12378 61896 12384
rect 61936 11620 61988 11626
rect 61936 11562 61988 11568
rect 61948 11354 61976 11562
rect 61936 11348 61988 11354
rect 61936 11290 61988 11296
rect 61764 11206 61976 11234
rect 61384 11144 61436 11150
rect 61384 11086 61436 11092
rect 61948 11014 61976 11206
rect 61844 11008 61896 11014
rect 61844 10950 61896 10956
rect 61936 11008 61988 11014
rect 61936 10950 61988 10956
rect 61856 10441 61884 10950
rect 61936 10532 61988 10538
rect 61936 10474 61988 10480
rect 61842 10432 61898 10441
rect 61842 10367 61898 10376
rect 61948 10198 61976 10474
rect 61936 10192 61988 10198
rect 61936 10134 61988 10140
rect 61292 2644 61344 2650
rect 61292 2586 61344 2592
rect 59912 2440 59964 2446
rect 59912 2382 59964 2388
rect 61200 2440 61252 2446
rect 61200 2382 61252 2388
rect 59360 1964 59412 1970
rect 59360 1906 59412 1912
rect 59924 800 59952 2382
rect 61212 800 61240 2382
rect 61844 2304 61896 2310
rect 61844 2246 61896 2252
rect 61856 800 61884 2246
rect 62040 2106 62068 13874
rect 62120 13728 62172 13734
rect 62118 13696 62120 13705
rect 62172 13696 62174 13705
rect 62118 13631 62174 13640
rect 62224 13326 62252 15535
rect 62396 15428 62448 15434
rect 62396 15370 62448 15376
rect 62302 15192 62358 15201
rect 62302 15127 62358 15136
rect 62316 15026 62344 15127
rect 62408 15065 62436 15370
rect 62394 15056 62450 15065
rect 62304 15020 62356 15026
rect 62394 14991 62396 15000
rect 62304 14962 62356 14968
rect 62448 14991 62450 15000
rect 62396 14962 62448 14968
rect 62500 14940 62528 17614
rect 62580 17536 62632 17542
rect 62578 17504 62580 17513
rect 62632 17504 62634 17513
rect 62578 17439 62634 17448
rect 62592 16998 62620 17439
rect 62684 17270 62712 17700
rect 62764 17682 62816 17688
rect 62672 17264 62724 17270
rect 62672 17206 62724 17212
rect 62580 16992 62632 16998
rect 62580 16934 62632 16940
rect 62580 16584 62632 16590
rect 62580 16526 62632 16532
rect 62592 15570 62620 16526
rect 62684 15609 62712 17206
rect 63052 16726 63080 16757
rect 63040 16720 63092 16726
rect 63038 16688 63040 16697
rect 63092 16688 63094 16697
rect 63038 16623 63094 16632
rect 62764 16584 62816 16590
rect 62764 16526 62816 16532
rect 62776 16114 62804 16526
rect 63052 16114 63080 16623
rect 63132 16516 63184 16522
rect 63132 16458 63184 16464
rect 62764 16108 62816 16114
rect 62764 16050 62816 16056
rect 63040 16108 63092 16114
rect 63040 16050 63092 16056
rect 62670 15600 62726 15609
rect 62580 15564 62632 15570
rect 62670 15535 62672 15544
rect 62580 15506 62632 15512
rect 62724 15535 62726 15544
rect 62672 15506 62724 15512
rect 62592 15065 62620 15506
rect 62684 15475 62712 15506
rect 62672 15360 62724 15366
rect 62672 15302 62724 15308
rect 62578 15056 62634 15065
rect 62578 14991 62634 15000
rect 62500 14912 62620 14940
rect 62592 14396 62620 14912
rect 62684 14414 62712 15302
rect 62776 14958 62804 16050
rect 62856 15632 62908 15638
rect 62856 15574 62908 15580
rect 62764 14952 62816 14958
rect 62764 14894 62816 14900
rect 62500 14368 62620 14396
rect 62672 14408 62724 14414
rect 62304 14000 62356 14006
rect 62304 13942 62356 13948
rect 62316 13569 62344 13942
rect 62500 13938 62528 14368
rect 62672 14350 62724 14356
rect 62488 13932 62540 13938
rect 62488 13874 62540 13880
rect 62580 13864 62632 13870
rect 62580 13806 62632 13812
rect 62396 13728 62448 13734
rect 62396 13670 62448 13676
rect 62302 13560 62358 13569
rect 62302 13495 62358 13504
rect 62212 13320 62264 13326
rect 62212 13262 62264 13268
rect 62224 12986 62252 13262
rect 62212 12980 62264 12986
rect 62212 12922 62264 12928
rect 62304 12232 62356 12238
rect 62304 12174 62356 12180
rect 62316 12073 62344 12174
rect 62408 12170 62436 13670
rect 62486 12336 62542 12345
rect 62486 12271 62542 12280
rect 62396 12164 62448 12170
rect 62396 12106 62448 12112
rect 62302 12064 62358 12073
rect 62302 11999 62358 12008
rect 62120 11688 62172 11694
rect 62120 11630 62172 11636
rect 62132 10538 62160 11630
rect 62304 11552 62356 11558
rect 62304 11494 62356 11500
rect 62212 11280 62264 11286
rect 62212 11222 62264 11228
rect 62224 10674 62252 11222
rect 62212 10668 62264 10674
rect 62212 10610 62264 10616
rect 62120 10532 62172 10538
rect 62120 10474 62172 10480
rect 62316 10062 62344 11494
rect 62304 10056 62356 10062
rect 62304 9998 62356 10004
rect 62408 3534 62436 12106
rect 62500 11150 62528 12271
rect 62592 11354 62620 13806
rect 62672 13184 62724 13190
rect 62672 13126 62724 13132
rect 62684 12850 62712 13126
rect 62672 12844 62724 12850
rect 62672 12786 62724 12792
rect 62762 12608 62818 12617
rect 62762 12543 62818 12552
rect 62670 12472 62726 12481
rect 62670 12407 62726 12416
rect 62684 12238 62712 12407
rect 62672 12232 62724 12238
rect 62672 12174 62724 12180
rect 62776 12102 62804 12543
rect 62764 12096 62816 12102
rect 62764 12038 62816 12044
rect 62670 11792 62726 11801
rect 62670 11727 62726 11736
rect 62684 11354 62712 11727
rect 62580 11348 62632 11354
rect 62580 11290 62632 11296
rect 62672 11348 62724 11354
rect 62672 11290 62724 11296
rect 62488 11144 62540 11150
rect 62488 11086 62540 11092
rect 62776 11014 62804 12038
rect 62868 11150 62896 15574
rect 63040 15496 63092 15502
rect 63144 15484 63172 16458
rect 63236 16114 63264 21354
rect 63314 16824 63370 16833
rect 63314 16759 63370 16768
rect 63328 16454 63356 16759
rect 63316 16448 63368 16454
rect 63316 16390 63368 16396
rect 63224 16108 63276 16114
rect 63224 16050 63276 16056
rect 63092 15456 63172 15484
rect 63040 15438 63092 15444
rect 63130 15328 63186 15337
rect 63130 15263 63186 15272
rect 62948 15156 63000 15162
rect 62948 15098 63000 15104
rect 62960 14929 62988 15098
rect 62946 14920 63002 14929
rect 62946 14855 63002 14864
rect 63038 14104 63094 14113
rect 63038 14039 63094 14048
rect 63052 14006 63080 14039
rect 63040 14000 63092 14006
rect 63040 13942 63092 13948
rect 63040 12776 63092 12782
rect 63040 12718 63092 12724
rect 63052 12617 63080 12718
rect 63038 12608 63094 12617
rect 63038 12543 63094 12552
rect 63038 11928 63094 11937
rect 63038 11863 63094 11872
rect 62948 11824 63000 11830
rect 62948 11766 63000 11772
rect 62960 11529 62988 11766
rect 62946 11520 63002 11529
rect 62946 11455 63002 11464
rect 63052 11218 63080 11863
rect 63040 11212 63092 11218
rect 63040 11154 63092 11160
rect 62856 11144 62908 11150
rect 62856 11086 62908 11092
rect 62764 11008 62816 11014
rect 62868 10985 62896 11086
rect 62764 10950 62816 10956
rect 62854 10976 62910 10985
rect 62854 10911 62910 10920
rect 63038 10704 63094 10713
rect 63038 10639 63094 10648
rect 63052 10606 63080 10639
rect 63040 10600 63092 10606
rect 63040 10542 63092 10548
rect 62396 3528 62448 3534
rect 62396 3470 62448 3476
rect 63144 3058 63172 15263
rect 63236 14822 63264 16050
rect 63328 15609 63356 16390
rect 63314 15600 63370 15609
rect 63314 15535 63370 15544
rect 63224 14816 63276 14822
rect 63224 14758 63276 14764
rect 63222 14512 63278 14521
rect 63222 14447 63278 14456
rect 63236 13938 63264 14447
rect 63224 13932 63276 13938
rect 63224 13874 63276 13880
rect 63236 13025 63264 13874
rect 63316 13184 63368 13190
rect 63316 13126 63368 13132
rect 63222 13016 63278 13025
rect 63222 12951 63278 12960
rect 63236 12238 63264 12951
rect 63224 12232 63276 12238
rect 63328 12209 63356 13126
rect 63224 12174 63276 12180
rect 63314 12200 63370 12209
rect 63314 12135 63370 12144
rect 63420 11880 63448 24210
rect 64328 24200 64380 24206
rect 64328 24142 64380 24148
rect 63868 19508 63920 19514
rect 63868 19450 63920 19456
rect 63500 17196 63552 17202
rect 63500 17138 63552 17144
rect 63684 17196 63736 17202
rect 63684 17138 63736 17144
rect 63512 16794 63540 17138
rect 63500 16788 63552 16794
rect 63500 16730 63552 16736
rect 63590 15056 63646 15065
rect 63590 14991 63592 15000
rect 63644 14991 63646 15000
rect 63592 14962 63644 14968
rect 63592 14816 63644 14822
rect 63592 14758 63644 14764
rect 63604 14278 63632 14758
rect 63592 14272 63644 14278
rect 63592 14214 63644 14220
rect 63592 14000 63644 14006
rect 63592 13942 63644 13948
rect 63500 13932 63552 13938
rect 63500 13874 63552 13880
rect 63512 13841 63540 13874
rect 63498 13832 63554 13841
rect 63498 13767 63554 13776
rect 63512 12986 63540 13767
rect 63604 13530 63632 13942
rect 63592 13524 63644 13530
rect 63592 13466 63644 13472
rect 63500 12980 63552 12986
rect 63500 12922 63552 12928
rect 63590 12608 63646 12617
rect 63590 12543 63646 12552
rect 63500 12436 63552 12442
rect 63500 12378 63552 12384
rect 63328 11852 63448 11880
rect 63224 11552 63276 11558
rect 63224 11494 63276 11500
rect 63236 10674 63264 11494
rect 63328 11082 63356 11852
rect 63406 11792 63462 11801
rect 63406 11727 63408 11736
rect 63460 11727 63462 11736
rect 63408 11698 63460 11704
rect 63512 11642 63540 12378
rect 63604 12356 63632 12543
rect 63696 12481 63724 17138
rect 63776 15904 63828 15910
rect 63776 15846 63828 15852
rect 63788 15502 63816 15846
rect 63776 15496 63828 15502
rect 63776 15438 63828 15444
rect 63774 15328 63830 15337
rect 63774 15263 63830 15272
rect 63788 14414 63816 15263
rect 63880 14822 63908 19450
rect 64236 16992 64288 16998
rect 64236 16934 64288 16940
rect 64144 16720 64196 16726
rect 64144 16662 64196 16668
rect 64156 16572 64184 16662
rect 64248 16640 64276 16934
rect 64340 16794 64368 24142
rect 64432 17270 64460 27406
rect 64892 27130 64920 27526
rect 67008 27470 67036 29200
rect 67652 27470 67680 29200
rect 68664 27470 68692 29294
rect 68926 29200 68982 30000
rect 69570 29322 69626 30000
rect 70214 29322 70270 30000
rect 69570 29294 69888 29322
rect 69570 29200 69626 29294
rect 68940 27588 68968 29200
rect 69020 27600 69072 27606
rect 68940 27560 69020 27588
rect 69020 27542 69072 27548
rect 66260 27464 66312 27470
rect 66260 27406 66312 27412
rect 66444 27464 66496 27470
rect 66444 27406 66496 27412
rect 66996 27464 67048 27470
rect 66996 27406 67048 27412
rect 67640 27464 67692 27470
rect 67640 27406 67692 27412
rect 68652 27464 68704 27470
rect 68652 27406 68704 27412
rect 69388 27464 69440 27470
rect 69388 27406 69440 27412
rect 64880 27124 64932 27130
rect 64880 27066 64932 27072
rect 64512 26988 64564 26994
rect 64512 26930 64564 26936
rect 65616 26988 65668 26994
rect 65616 26930 65668 26936
rect 64524 17814 64552 26930
rect 65628 26586 65656 26930
rect 65064 26580 65116 26586
rect 65064 26522 65116 26528
rect 65616 26580 65668 26586
rect 65616 26522 65668 26528
rect 64972 19372 65024 19378
rect 64972 19314 65024 19320
rect 64880 18284 64932 18290
rect 64880 18226 64932 18232
rect 64512 17808 64564 17814
rect 64512 17750 64564 17756
rect 64524 17649 64552 17750
rect 64510 17640 64566 17649
rect 64510 17575 64566 17584
rect 64420 17264 64472 17270
rect 64420 17206 64472 17212
rect 64788 17196 64840 17202
rect 64788 17138 64840 17144
rect 64696 17128 64748 17134
rect 64696 17070 64748 17076
rect 64708 16969 64736 17070
rect 64694 16960 64750 16969
rect 64694 16895 64750 16904
rect 64328 16788 64380 16794
rect 64328 16730 64380 16736
rect 64800 16726 64828 17138
rect 64788 16720 64840 16726
rect 64788 16662 64840 16668
rect 64248 16612 64552 16640
rect 64156 16544 64276 16572
rect 64144 15564 64196 15570
rect 64144 15506 64196 15512
rect 64156 15366 64184 15506
rect 64144 15360 64196 15366
rect 64144 15302 64196 15308
rect 63960 14884 64012 14890
rect 63960 14826 64012 14832
rect 63868 14816 63920 14822
rect 63868 14758 63920 14764
rect 63972 14414 64000 14826
rect 63776 14408 63828 14414
rect 63776 14350 63828 14356
rect 63960 14408 64012 14414
rect 64052 14408 64104 14414
rect 63960 14350 64012 14356
rect 64050 14376 64052 14385
rect 64104 14376 64106 14385
rect 63788 12617 63816 14350
rect 64248 14362 64276 16544
rect 64328 15360 64380 15366
rect 64328 15302 64380 15308
rect 64340 15162 64368 15302
rect 64328 15156 64380 15162
rect 64328 15098 64380 15104
rect 64420 14408 64472 14414
rect 64248 14334 64368 14362
rect 64420 14350 64472 14356
rect 64050 14311 64106 14320
rect 64144 14272 64196 14278
rect 64144 14214 64196 14220
rect 64050 14104 64106 14113
rect 64050 14039 64106 14048
rect 64064 13938 64092 14039
rect 64052 13932 64104 13938
rect 64052 13874 64104 13880
rect 63960 13864 64012 13870
rect 63960 13806 64012 13812
rect 63868 13728 63920 13734
rect 63868 13670 63920 13676
rect 63774 12608 63830 12617
rect 63774 12543 63830 12552
rect 63682 12472 63738 12481
rect 63682 12407 63738 12416
rect 63604 12328 63724 12356
rect 63590 12200 63646 12209
rect 63590 12135 63646 12144
rect 63604 11830 63632 12135
rect 63592 11824 63644 11830
rect 63592 11766 63644 11772
rect 63592 11688 63644 11694
rect 63420 11614 63540 11642
rect 63590 11656 63592 11665
rect 63644 11656 63646 11665
rect 63316 11076 63368 11082
rect 63316 11018 63368 11024
rect 63224 10668 63276 10674
rect 63224 10610 63276 10616
rect 63328 9674 63356 11018
rect 63420 10849 63448 11614
rect 63590 11591 63646 11600
rect 63590 11520 63646 11529
rect 63590 11455 63646 11464
rect 63406 10840 63462 10849
rect 63406 10775 63462 10784
rect 63406 10704 63462 10713
rect 63406 10639 63408 10648
rect 63460 10639 63462 10648
rect 63408 10610 63460 10616
rect 63236 9646 63356 9674
rect 63236 4826 63264 9646
rect 63420 9518 63448 10610
rect 63498 10296 63554 10305
rect 63498 10231 63554 10240
rect 63408 9512 63460 9518
rect 63408 9454 63460 9460
rect 63408 9376 63460 9382
rect 63408 9318 63460 9324
rect 63224 4820 63276 4826
rect 63224 4762 63276 4768
rect 63132 3052 63184 3058
rect 63132 2994 63184 3000
rect 62488 2848 62540 2854
rect 62488 2790 62540 2796
rect 62212 2508 62264 2514
rect 62212 2450 62264 2456
rect 62028 2100 62080 2106
rect 62028 2042 62080 2048
rect 62224 1494 62252 2450
rect 62304 1896 62356 1902
rect 62304 1838 62356 1844
rect 62316 1494 62344 1838
rect 62212 1488 62264 1494
rect 62212 1430 62264 1436
rect 62304 1488 62356 1494
rect 62304 1430 62356 1436
rect 62500 800 62528 2790
rect 63132 2440 63184 2446
rect 63132 2382 63184 2388
rect 63144 800 63172 2382
rect 63420 1970 63448 9318
rect 63512 3194 63540 10231
rect 63604 4146 63632 11455
rect 63696 10742 63724 12328
rect 63774 11928 63830 11937
rect 63774 11863 63830 11872
rect 63684 10736 63736 10742
rect 63684 10678 63736 10684
rect 63788 10577 63816 11863
rect 63774 10568 63830 10577
rect 63774 10503 63830 10512
rect 63592 4140 63644 4146
rect 63592 4082 63644 4088
rect 63500 3188 63552 3194
rect 63500 3130 63552 3136
rect 63788 2774 63816 10503
rect 63880 4010 63908 13670
rect 63972 12986 64000 13806
rect 64050 13152 64106 13161
rect 64050 13087 64106 13096
rect 63960 12980 64012 12986
rect 63960 12922 64012 12928
rect 63972 6186 64000 12922
rect 64064 12782 64092 13087
rect 64052 12776 64104 12782
rect 64052 12718 64104 12724
rect 64052 12232 64104 12238
rect 64052 12174 64104 12180
rect 64064 11801 64092 12174
rect 64050 11792 64106 11801
rect 64050 11727 64052 11736
rect 64104 11727 64106 11736
rect 64052 11698 64104 11704
rect 64064 11150 64092 11698
rect 64052 11144 64104 11150
rect 64052 11086 64104 11092
rect 63960 6180 64012 6186
rect 63960 6122 64012 6128
rect 64052 4140 64104 4146
rect 64052 4082 64104 4088
rect 63868 4004 63920 4010
rect 63868 3946 63920 3952
rect 63696 2746 63816 2774
rect 63696 2650 63724 2746
rect 63684 2644 63736 2650
rect 63684 2586 63736 2592
rect 63500 2440 63552 2446
rect 63500 2382 63552 2388
rect 63408 1964 63460 1970
rect 63408 1906 63460 1912
rect 63512 1426 63540 2382
rect 64064 1426 64092 4082
rect 64156 3738 64184 14214
rect 64340 14090 64368 14334
rect 64432 14249 64460 14350
rect 64418 14240 64474 14249
rect 64418 14175 64474 14184
rect 64340 14062 64460 14090
rect 64524 14074 64552 16612
rect 64892 16114 64920 18226
rect 64984 17202 65012 19314
rect 64972 17196 65024 17202
rect 64972 17138 65024 17144
rect 64604 16108 64656 16114
rect 64880 16108 64932 16114
rect 64656 16068 64736 16096
rect 64604 16050 64656 16056
rect 64604 15360 64656 15366
rect 64604 15302 64656 15308
rect 64616 15026 64644 15302
rect 64708 15201 64736 16068
rect 64880 16050 64932 16056
rect 64984 15910 65012 17138
rect 64972 15904 65024 15910
rect 64972 15846 65024 15852
rect 64880 15496 64932 15502
rect 64880 15438 64932 15444
rect 64694 15192 64750 15201
rect 64694 15127 64750 15136
rect 64604 15020 64656 15026
rect 64604 14962 64656 14968
rect 64604 14816 64656 14822
rect 64604 14758 64656 14764
rect 64616 14482 64644 14758
rect 64604 14476 64656 14482
rect 64604 14418 64656 14424
rect 64892 14074 64920 15438
rect 64970 15192 65026 15201
rect 64970 15127 65026 15136
rect 64984 14482 65012 15127
rect 64972 14476 65024 14482
rect 64972 14418 65024 14424
rect 64972 14272 65024 14278
rect 64972 14214 65024 14220
rect 64432 13818 64460 14062
rect 64512 14068 64564 14074
rect 64512 14010 64564 14016
rect 64880 14068 64932 14074
rect 64880 14010 64932 14016
rect 64984 13938 65012 14214
rect 64604 13932 64656 13938
rect 64604 13874 64656 13880
rect 64972 13932 65024 13938
rect 64972 13874 65024 13880
rect 64616 13818 64644 13874
rect 64432 13790 64644 13818
rect 64512 13524 64564 13530
rect 64512 13466 64564 13472
rect 64420 13456 64472 13462
rect 64420 13398 64472 13404
rect 64328 13184 64380 13190
rect 64328 13126 64380 13132
rect 64340 11642 64368 13126
rect 64432 12170 64460 13398
rect 64524 13297 64552 13466
rect 64510 13288 64566 13297
rect 64510 13223 64566 13232
rect 64604 13184 64656 13190
rect 64604 13126 64656 13132
rect 64616 12918 64644 13126
rect 64604 12912 64656 12918
rect 64604 12854 64656 12860
rect 64512 12708 64564 12714
rect 64512 12650 64564 12656
rect 64524 12238 64552 12650
rect 64788 12436 64840 12442
rect 64788 12378 64840 12384
rect 64512 12232 64564 12238
rect 64696 12232 64748 12238
rect 64512 12174 64564 12180
rect 64616 12192 64696 12220
rect 64420 12164 64472 12170
rect 64420 12106 64472 12112
rect 64340 11614 64460 11642
rect 64326 11248 64382 11257
rect 64326 11183 64382 11192
rect 64340 11150 64368 11183
rect 64236 11144 64288 11150
rect 64236 11086 64288 11092
rect 64328 11144 64380 11150
rect 64328 11086 64380 11092
rect 64248 10146 64276 11086
rect 64248 10118 64368 10146
rect 64236 10056 64288 10062
rect 64236 9998 64288 10004
rect 64248 9654 64276 9998
rect 64236 9648 64288 9654
rect 64236 9590 64288 9596
rect 64340 7886 64368 10118
rect 64328 7880 64380 7886
rect 64328 7822 64380 7828
rect 64432 7698 64460 11614
rect 64512 11144 64564 11150
rect 64510 11112 64512 11121
rect 64564 11112 64566 11121
rect 64510 11047 64566 11056
rect 64340 7670 64460 7698
rect 64144 3732 64196 3738
rect 64144 3674 64196 3680
rect 64340 2774 64368 7670
rect 64420 2984 64472 2990
rect 64420 2926 64472 2932
rect 64156 2746 64368 2774
rect 64156 1902 64184 2746
rect 64144 1896 64196 1902
rect 64144 1838 64196 1844
rect 63500 1420 63552 1426
rect 63500 1362 63552 1368
rect 64052 1420 64104 1426
rect 64052 1362 64104 1368
rect 64432 800 64460 2926
rect 64524 2774 64552 11047
rect 64616 10266 64644 12192
rect 64696 12174 64748 12180
rect 64800 12050 64828 12378
rect 64878 12336 64934 12345
rect 64878 12271 64934 12280
rect 64892 12170 64920 12271
rect 64880 12164 64932 12170
rect 64880 12106 64932 12112
rect 64800 12022 64920 12050
rect 64892 11898 64920 12022
rect 64788 11892 64840 11898
rect 64788 11834 64840 11840
rect 64880 11892 64932 11898
rect 64880 11834 64932 11840
rect 64696 11756 64748 11762
rect 64696 11698 64748 11704
rect 64708 11558 64736 11698
rect 64696 11552 64748 11558
rect 64696 11494 64748 11500
rect 64604 10260 64656 10266
rect 64604 10202 64656 10208
rect 64708 10130 64736 11494
rect 64800 10538 64828 11834
rect 64878 11112 64934 11121
rect 64878 11047 64934 11056
rect 64788 10532 64840 10538
rect 64788 10474 64840 10480
rect 64696 10124 64748 10130
rect 64696 10066 64748 10072
rect 64708 9722 64736 10066
rect 64800 10062 64828 10474
rect 64892 10470 64920 11047
rect 64880 10464 64932 10470
rect 64880 10406 64932 10412
rect 64788 10056 64840 10062
rect 64788 9998 64840 10004
rect 64696 9716 64748 9722
rect 64696 9658 64748 9664
rect 64524 2746 64736 2774
rect 64708 2106 64736 2746
rect 64984 2514 65012 13874
rect 65076 12986 65104 26522
rect 65524 17808 65576 17814
rect 65524 17750 65576 17756
rect 65156 17672 65208 17678
rect 65156 17614 65208 17620
rect 65168 17066 65196 17614
rect 65536 17610 65564 17750
rect 65524 17604 65576 17610
rect 65524 17546 65576 17552
rect 65156 17060 65208 17066
rect 65156 17002 65208 17008
rect 65340 16992 65392 16998
rect 66272 16969 66300 27406
rect 66456 27130 66484 27406
rect 68192 27396 68244 27402
rect 68192 27338 68244 27344
rect 67456 27328 67508 27334
rect 67456 27270 67508 27276
rect 66794 27228 67102 27237
rect 66794 27226 66800 27228
rect 66856 27226 66880 27228
rect 66936 27226 66960 27228
rect 67016 27226 67040 27228
rect 67096 27226 67102 27228
rect 66856 27174 66858 27226
rect 67038 27174 67040 27226
rect 66794 27172 66800 27174
rect 66856 27172 66880 27174
rect 66936 27172 66960 27174
rect 67016 27172 67040 27174
rect 67096 27172 67102 27174
rect 66794 27163 67102 27172
rect 66444 27124 66496 27130
rect 66444 27066 66496 27072
rect 66794 26140 67102 26149
rect 66794 26138 66800 26140
rect 66856 26138 66880 26140
rect 66936 26138 66960 26140
rect 67016 26138 67040 26140
rect 67096 26138 67102 26140
rect 66856 26086 66858 26138
rect 67038 26086 67040 26138
rect 66794 26084 66800 26086
rect 66856 26084 66880 26086
rect 66936 26084 66960 26086
rect 67016 26084 67040 26086
rect 67096 26084 67102 26086
rect 66794 26075 67102 26084
rect 66794 25052 67102 25061
rect 66794 25050 66800 25052
rect 66856 25050 66880 25052
rect 66936 25050 66960 25052
rect 67016 25050 67040 25052
rect 67096 25050 67102 25052
rect 66856 24998 66858 25050
rect 67038 24998 67040 25050
rect 66794 24996 66800 24998
rect 66856 24996 66880 24998
rect 66936 24996 66960 24998
rect 67016 24996 67040 24998
rect 67096 24996 67102 24998
rect 66794 24987 67102 24996
rect 66794 23964 67102 23973
rect 66794 23962 66800 23964
rect 66856 23962 66880 23964
rect 66936 23962 66960 23964
rect 67016 23962 67040 23964
rect 67096 23962 67102 23964
rect 66856 23910 66858 23962
rect 67038 23910 67040 23962
rect 66794 23908 66800 23910
rect 66856 23908 66880 23910
rect 66936 23908 66960 23910
rect 67016 23908 67040 23910
rect 67096 23908 67102 23910
rect 66794 23899 67102 23908
rect 66794 22876 67102 22885
rect 66794 22874 66800 22876
rect 66856 22874 66880 22876
rect 66936 22874 66960 22876
rect 67016 22874 67040 22876
rect 67096 22874 67102 22876
rect 66856 22822 66858 22874
rect 67038 22822 67040 22874
rect 66794 22820 66800 22822
rect 66856 22820 66880 22822
rect 66936 22820 66960 22822
rect 67016 22820 67040 22822
rect 67096 22820 67102 22822
rect 66794 22811 67102 22820
rect 66794 21788 67102 21797
rect 66794 21786 66800 21788
rect 66856 21786 66880 21788
rect 66936 21786 66960 21788
rect 67016 21786 67040 21788
rect 67096 21786 67102 21788
rect 66856 21734 66858 21786
rect 67038 21734 67040 21786
rect 66794 21732 66800 21734
rect 66856 21732 66880 21734
rect 66936 21732 66960 21734
rect 67016 21732 67040 21734
rect 67096 21732 67102 21734
rect 66794 21723 67102 21732
rect 66794 20700 67102 20709
rect 66794 20698 66800 20700
rect 66856 20698 66880 20700
rect 66936 20698 66960 20700
rect 67016 20698 67040 20700
rect 67096 20698 67102 20700
rect 66856 20646 66858 20698
rect 67038 20646 67040 20698
rect 66794 20644 66800 20646
rect 66856 20644 66880 20646
rect 66936 20644 66960 20646
rect 67016 20644 67040 20646
rect 67096 20644 67102 20646
rect 66794 20635 67102 20644
rect 66794 19612 67102 19621
rect 66794 19610 66800 19612
rect 66856 19610 66880 19612
rect 66936 19610 66960 19612
rect 67016 19610 67040 19612
rect 67096 19610 67102 19612
rect 66856 19558 66858 19610
rect 67038 19558 67040 19610
rect 66794 19556 66800 19558
rect 66856 19556 66880 19558
rect 66936 19556 66960 19558
rect 67016 19556 67040 19558
rect 67096 19556 67102 19558
rect 66794 19547 67102 19556
rect 66794 18524 67102 18533
rect 66794 18522 66800 18524
rect 66856 18522 66880 18524
rect 66936 18522 66960 18524
rect 67016 18522 67040 18524
rect 67096 18522 67102 18524
rect 66856 18470 66858 18522
rect 67038 18470 67040 18522
rect 66794 18468 66800 18470
rect 66856 18468 66880 18470
rect 66936 18468 66960 18470
rect 67016 18468 67040 18470
rect 67096 18468 67102 18470
rect 66794 18459 67102 18468
rect 67468 18426 67496 27270
rect 68008 18692 68060 18698
rect 68008 18634 68060 18640
rect 67456 18420 67508 18426
rect 67456 18362 67508 18368
rect 67364 18148 67416 18154
rect 67364 18090 67416 18096
rect 66720 17536 66772 17542
rect 66720 17478 66772 17484
rect 66534 17368 66590 17377
rect 66534 17303 66590 17312
rect 66548 17134 66576 17303
rect 66732 17202 66760 17478
rect 66794 17436 67102 17445
rect 66794 17434 66800 17436
rect 66856 17434 66880 17436
rect 66936 17434 66960 17436
rect 67016 17434 67040 17436
rect 67096 17434 67102 17436
rect 66856 17382 66858 17434
rect 67038 17382 67040 17434
rect 66794 17380 66800 17382
rect 66856 17380 66880 17382
rect 66936 17380 66960 17382
rect 67016 17380 67040 17382
rect 67096 17380 67102 17382
rect 66794 17371 67102 17380
rect 66994 17232 67050 17241
rect 66720 17196 66772 17202
rect 66994 17167 66996 17176
rect 66720 17138 66772 17144
rect 67048 17167 67050 17176
rect 66996 17138 67048 17144
rect 66444 17128 66496 17134
rect 66442 17096 66444 17105
rect 66536 17128 66588 17134
rect 66496 17096 66498 17105
rect 66536 17070 66588 17076
rect 66442 17031 66498 17040
rect 65340 16934 65392 16940
rect 66258 16960 66314 16969
rect 65248 16652 65300 16658
rect 65248 16594 65300 16600
rect 65260 15502 65288 16594
rect 65352 16590 65380 16934
rect 66258 16895 66314 16904
rect 65524 16652 65576 16658
rect 65524 16594 65576 16600
rect 65340 16584 65392 16590
rect 65340 16526 65392 16532
rect 65340 16448 65392 16454
rect 65340 16390 65392 16396
rect 65352 15570 65380 16390
rect 65340 15564 65392 15570
rect 65340 15506 65392 15512
rect 65248 15496 65300 15502
rect 65248 15438 65300 15444
rect 65536 15162 65564 16594
rect 66456 16561 66484 17031
rect 66442 16552 66498 16561
rect 66442 16487 66498 16496
rect 65984 16448 66036 16454
rect 65984 16390 66036 16396
rect 65996 16250 66024 16390
rect 66794 16348 67102 16357
rect 66794 16346 66800 16348
rect 66856 16346 66880 16348
rect 66936 16346 66960 16348
rect 67016 16346 67040 16348
rect 67096 16346 67102 16348
rect 66856 16294 66858 16346
rect 67038 16294 67040 16346
rect 66794 16292 66800 16294
rect 66856 16292 66880 16294
rect 66936 16292 66960 16294
rect 67016 16292 67040 16294
rect 67096 16292 67102 16294
rect 66794 16283 67102 16292
rect 65984 16244 66036 16250
rect 65984 16186 66036 16192
rect 66076 16244 66128 16250
rect 66076 16186 66128 16192
rect 66088 16153 66116 16186
rect 66074 16144 66130 16153
rect 65708 16108 65760 16114
rect 66074 16079 66130 16088
rect 65708 16050 65760 16056
rect 65616 15904 65668 15910
rect 65616 15846 65668 15852
rect 65628 15706 65656 15846
rect 65616 15700 65668 15706
rect 65616 15642 65668 15648
rect 65524 15156 65576 15162
rect 65524 15098 65576 15104
rect 65248 15088 65300 15094
rect 65720 15065 65748 16050
rect 66444 16040 66496 16046
rect 66444 15982 66496 15988
rect 65800 15496 65852 15502
rect 65800 15438 65852 15444
rect 65248 15030 65300 15036
rect 65706 15056 65762 15065
rect 65260 14929 65288 15030
rect 65706 14991 65708 15000
rect 65760 14991 65762 15000
rect 65708 14962 65760 14968
rect 65720 14931 65748 14962
rect 65812 14958 65840 15438
rect 66456 15026 66484 15982
rect 67272 15564 67324 15570
rect 67272 15506 67324 15512
rect 66794 15260 67102 15269
rect 66794 15258 66800 15260
rect 66856 15258 66880 15260
rect 66936 15258 66960 15260
rect 67016 15258 67040 15260
rect 67096 15258 67102 15260
rect 66856 15206 66858 15258
rect 67038 15206 67040 15258
rect 66794 15204 66800 15206
rect 66856 15204 66880 15206
rect 66936 15204 66960 15206
rect 67016 15204 67040 15206
rect 67096 15204 67102 15206
rect 66794 15195 67102 15204
rect 67284 15162 67312 15506
rect 67272 15156 67324 15162
rect 67272 15098 67324 15104
rect 66444 15020 66496 15026
rect 66444 14962 66496 14968
rect 65800 14952 65852 14958
rect 65246 14920 65302 14929
rect 65800 14894 65852 14900
rect 65246 14855 65302 14864
rect 65340 14884 65392 14890
rect 65340 14826 65392 14832
rect 65352 14482 65380 14826
rect 65340 14476 65392 14482
rect 65340 14418 65392 14424
rect 65812 14113 65840 14894
rect 66718 14784 66774 14793
rect 66718 14719 66774 14728
rect 66732 14414 66760 14719
rect 66536 14408 66588 14414
rect 66536 14350 66588 14356
rect 66720 14408 66772 14414
rect 66720 14350 66772 14356
rect 65798 14104 65854 14113
rect 65798 14039 65854 14048
rect 65156 13932 65208 13938
rect 65156 13874 65208 13880
rect 65168 13705 65196 13874
rect 65154 13696 65210 13705
rect 65154 13631 65210 13640
rect 66350 13560 66406 13569
rect 66350 13495 66406 13504
rect 66260 13456 66312 13462
rect 66260 13398 66312 13404
rect 65064 12980 65116 12986
rect 65064 12922 65116 12928
rect 66272 12850 66300 13398
rect 66364 12986 66392 13495
rect 66352 12980 66404 12986
rect 66352 12922 66404 12928
rect 66364 12850 66392 12922
rect 65156 12844 65208 12850
rect 65156 12786 65208 12792
rect 65340 12844 65392 12850
rect 65340 12786 65392 12792
rect 66260 12844 66312 12850
rect 66260 12786 66312 12792
rect 66352 12844 66404 12850
rect 66352 12786 66404 12792
rect 65168 12442 65196 12786
rect 65156 12436 65208 12442
rect 65156 12378 65208 12384
rect 65352 12238 65380 12786
rect 66260 12640 66312 12646
rect 66260 12582 66312 12588
rect 65984 12436 66036 12442
rect 65984 12378 66036 12384
rect 65996 12345 66024 12378
rect 65982 12336 66038 12345
rect 65982 12271 66038 12280
rect 65340 12232 65392 12238
rect 65340 12174 65392 12180
rect 66166 12064 66222 12073
rect 66166 11999 66222 12008
rect 65156 11824 65208 11830
rect 65156 11766 65208 11772
rect 65168 11218 65196 11766
rect 66180 11762 66208 11999
rect 66272 11762 66300 12582
rect 66548 12238 66576 14350
rect 66794 14172 67102 14181
rect 66794 14170 66800 14172
rect 66856 14170 66880 14172
rect 66936 14170 66960 14172
rect 67016 14170 67040 14172
rect 67096 14170 67102 14172
rect 66856 14118 66858 14170
rect 67038 14118 67040 14170
rect 66794 14116 66800 14118
rect 66856 14116 66880 14118
rect 66936 14116 66960 14118
rect 67016 14116 67040 14118
rect 67096 14116 67102 14118
rect 66794 14107 67102 14116
rect 66794 13084 67102 13093
rect 66794 13082 66800 13084
rect 66856 13082 66880 13084
rect 66936 13082 66960 13084
rect 67016 13082 67040 13084
rect 67096 13082 67102 13084
rect 66856 13030 66858 13082
rect 67038 13030 67040 13082
rect 66794 13028 66800 13030
rect 66856 13028 66880 13030
rect 66936 13028 66960 13030
rect 67016 13028 67040 13030
rect 67096 13028 67102 13030
rect 66626 13016 66682 13025
rect 66794 13019 67102 13028
rect 66626 12951 66682 12960
rect 66640 12832 66668 12951
rect 66720 12844 66772 12850
rect 66640 12804 66720 12832
rect 66720 12786 66772 12792
rect 67376 12434 67404 18090
rect 67824 15360 67876 15366
rect 67824 15302 67876 15308
rect 67456 14476 67508 14482
rect 67456 14418 67508 14424
rect 67468 14385 67496 14418
rect 67836 14385 67864 15302
rect 68020 15094 68048 18634
rect 68100 18080 68152 18086
rect 68100 18022 68152 18028
rect 68112 17678 68140 18022
rect 68100 17672 68152 17678
rect 68100 17614 68152 17620
rect 68100 16040 68152 16046
rect 68100 15982 68152 15988
rect 68008 15088 68060 15094
rect 68008 15030 68060 15036
rect 67454 14376 67510 14385
rect 67454 14311 67510 14320
rect 67822 14376 67878 14385
rect 67822 14311 67878 14320
rect 67454 14240 67510 14249
rect 67454 14175 67510 14184
rect 67468 14006 67496 14175
rect 67730 14104 67786 14113
rect 67730 14039 67732 14048
rect 67784 14039 67786 14048
rect 68008 14068 68060 14074
rect 67732 14010 67784 14016
rect 68008 14010 68060 14016
rect 67456 14000 67508 14006
rect 67456 13942 67508 13948
rect 67732 13932 67784 13938
rect 67732 13874 67784 13880
rect 67454 13832 67510 13841
rect 67454 13767 67510 13776
rect 67468 12850 67496 13767
rect 67640 13252 67692 13258
rect 67640 13194 67692 13200
rect 67456 12844 67508 12850
rect 67456 12786 67508 12792
rect 67652 12481 67680 13194
rect 67744 13161 67772 13874
rect 68020 13870 68048 14010
rect 68008 13864 68060 13870
rect 68008 13806 68060 13812
rect 68112 13274 68140 15982
rect 68204 13802 68232 27338
rect 68652 27328 68704 27334
rect 68652 27270 68704 27276
rect 68468 27056 68520 27062
rect 68468 26998 68520 27004
rect 68480 22094 68508 26998
rect 68560 26784 68612 26790
rect 68560 26726 68612 26732
rect 68572 26518 68600 26726
rect 68560 26512 68612 26518
rect 68560 26454 68612 26460
rect 68388 22066 68508 22094
rect 68284 17604 68336 17610
rect 68284 17546 68336 17552
rect 68192 13796 68244 13802
rect 68192 13738 68244 13744
rect 68112 13258 68232 13274
rect 68112 13252 68244 13258
rect 68112 13246 68192 13252
rect 68192 13194 68244 13200
rect 68100 13184 68152 13190
rect 67730 13152 67786 13161
rect 68100 13126 68152 13132
rect 67730 13087 67786 13096
rect 67916 12912 67968 12918
rect 67916 12854 67968 12860
rect 67638 12472 67694 12481
rect 67548 12436 67600 12442
rect 67376 12406 67496 12434
rect 66536 12232 66588 12238
rect 66536 12174 66588 12180
rect 66168 11756 66220 11762
rect 66168 11698 66220 11704
rect 66260 11756 66312 11762
rect 66260 11698 66312 11704
rect 65156 11212 65208 11218
rect 65156 11154 65208 11160
rect 65168 10470 65196 11154
rect 65616 10668 65668 10674
rect 65616 10610 65668 10616
rect 65156 10464 65208 10470
rect 65156 10406 65208 10412
rect 65168 9382 65196 10406
rect 65628 10266 65656 10610
rect 65616 10260 65668 10266
rect 65616 10202 65668 10208
rect 65156 9376 65208 9382
rect 65156 9318 65208 9324
rect 64972 2508 65024 2514
rect 64972 2450 65024 2456
rect 66272 2446 66300 11698
rect 66548 11257 66576 12174
rect 67180 12164 67232 12170
rect 67180 12106 67232 12112
rect 67272 12164 67324 12170
rect 67272 12106 67324 12112
rect 66794 11996 67102 12005
rect 66794 11994 66800 11996
rect 66856 11994 66880 11996
rect 66936 11994 66960 11996
rect 67016 11994 67040 11996
rect 67096 11994 67102 11996
rect 66856 11942 66858 11994
rect 67038 11942 67040 11994
rect 66794 11940 66800 11942
rect 66856 11940 66880 11942
rect 66936 11940 66960 11942
rect 67016 11940 67040 11942
rect 67096 11940 67102 11942
rect 66794 11931 67102 11940
rect 67192 11898 67220 12106
rect 67284 11898 67312 12106
rect 66812 11892 66864 11898
rect 66812 11834 66864 11840
rect 67180 11892 67232 11898
rect 67180 11834 67232 11840
rect 67272 11892 67324 11898
rect 67272 11834 67324 11840
rect 66824 11665 66852 11834
rect 66996 11824 67048 11830
rect 66994 11792 66996 11801
rect 67048 11792 67050 11801
rect 67364 11756 67416 11762
rect 66994 11727 67050 11736
rect 67192 11716 67364 11744
rect 66810 11656 66866 11665
rect 67192 11626 67220 11716
rect 67364 11698 67416 11704
rect 67468 11642 67496 12406
rect 67928 12442 67956 12854
rect 67638 12407 67694 12416
rect 67916 12436 67968 12442
rect 67548 12378 67600 12384
rect 67916 12378 67968 12384
rect 67560 11898 67588 12378
rect 68112 12102 68140 13126
rect 68100 12096 68152 12102
rect 68100 12038 68152 12044
rect 67548 11892 67600 11898
rect 67548 11834 67600 11840
rect 67560 11694 67588 11834
rect 66810 11591 66866 11600
rect 67180 11620 67232 11626
rect 67180 11562 67232 11568
rect 67272 11620 67324 11626
rect 67272 11562 67324 11568
rect 67376 11614 67496 11642
rect 67548 11688 67600 11694
rect 67548 11630 67600 11636
rect 67088 11552 67140 11558
rect 67088 11494 67140 11500
rect 66534 11248 66590 11257
rect 67100 11218 67128 11494
rect 66534 11183 66590 11192
rect 67088 11212 67140 11218
rect 66548 10674 66576 11183
rect 67088 11154 67140 11160
rect 67284 11150 67312 11562
rect 67272 11144 67324 11150
rect 67272 11086 67324 11092
rect 66794 10908 67102 10917
rect 66794 10906 66800 10908
rect 66856 10906 66880 10908
rect 66936 10906 66960 10908
rect 67016 10906 67040 10908
rect 67096 10906 67102 10908
rect 66856 10854 66858 10906
rect 67038 10854 67040 10906
rect 66794 10852 66800 10854
rect 66856 10852 66880 10854
rect 66936 10852 66960 10854
rect 67016 10852 67040 10854
rect 67096 10852 67102 10854
rect 66794 10843 67102 10852
rect 66536 10668 66588 10674
rect 66536 10610 66588 10616
rect 66794 9820 67102 9829
rect 66794 9818 66800 9820
rect 66856 9818 66880 9820
rect 66936 9818 66960 9820
rect 67016 9818 67040 9820
rect 67096 9818 67102 9820
rect 66856 9766 66858 9818
rect 67038 9766 67040 9818
rect 66794 9764 66800 9766
rect 66856 9764 66880 9766
rect 66936 9764 66960 9766
rect 67016 9764 67040 9766
rect 67096 9764 67102 9766
rect 66794 9755 67102 9764
rect 67376 9330 67404 11614
rect 67822 11384 67878 11393
rect 67732 11348 67784 11354
rect 67822 11319 67878 11328
rect 67732 11290 67784 11296
rect 67456 11280 67508 11286
rect 67548 11280 67600 11286
rect 67456 11222 67508 11228
rect 67546 11248 67548 11257
rect 67744 11257 67772 11290
rect 67600 11248 67602 11257
rect 67468 11132 67496 11222
rect 67546 11183 67602 11192
rect 67730 11248 67786 11257
rect 67836 11218 67864 11319
rect 67730 11183 67786 11192
rect 67824 11212 67876 11218
rect 67824 11154 67876 11160
rect 67468 11104 67588 11132
rect 67560 11064 67588 11104
rect 67640 11076 67692 11082
rect 67560 11036 67640 11064
rect 67640 11018 67692 11024
rect 67456 11008 67508 11014
rect 67456 10950 67508 10956
rect 67468 10441 67496 10950
rect 67548 10668 67600 10674
rect 67548 10610 67600 10616
rect 67454 10432 67510 10441
rect 67454 10367 67510 10376
rect 67560 9518 67588 10610
rect 68192 9580 68244 9586
rect 68192 9522 68244 9528
rect 67548 9512 67600 9518
rect 67548 9454 67600 9460
rect 67376 9302 67588 9330
rect 67560 9042 67588 9302
rect 68204 9178 68232 9522
rect 68296 9382 68324 17546
rect 68388 16454 68416 22066
rect 68468 17808 68520 17814
rect 68468 17750 68520 17756
rect 68480 17678 68508 17750
rect 68468 17672 68520 17678
rect 68468 17614 68520 17620
rect 68572 17610 68600 26454
rect 68664 19334 68692 27270
rect 69400 27130 69428 27406
rect 69480 27396 69532 27402
rect 69480 27338 69532 27344
rect 69388 27124 69440 27130
rect 69388 27066 69440 27072
rect 69204 26920 69256 26926
rect 69204 26862 69256 26868
rect 68928 26444 68980 26450
rect 68928 26386 68980 26392
rect 68940 25809 68968 26386
rect 68926 25800 68982 25809
rect 68926 25735 68982 25744
rect 68664 19306 68876 19334
rect 68560 17604 68612 17610
rect 68560 17546 68612 17552
rect 68560 17060 68612 17066
rect 68560 17002 68612 17008
rect 68652 17060 68704 17066
rect 68652 17002 68704 17008
rect 68572 16794 68600 17002
rect 68560 16788 68612 16794
rect 68560 16730 68612 16736
rect 68664 16522 68692 17002
rect 68652 16516 68704 16522
rect 68652 16458 68704 16464
rect 68376 16448 68428 16454
rect 68376 16390 68428 16396
rect 68560 16448 68612 16454
rect 68560 16390 68612 16396
rect 68376 14272 68428 14278
rect 68376 14214 68428 14220
rect 68468 14272 68520 14278
rect 68468 14214 68520 14220
rect 68388 13938 68416 14214
rect 68376 13932 68428 13938
rect 68376 13874 68428 13880
rect 68480 13326 68508 14214
rect 68468 13320 68520 13326
rect 68468 13262 68520 13268
rect 68376 13252 68428 13258
rect 68376 13194 68428 13200
rect 68388 12986 68416 13194
rect 68572 13190 68600 16390
rect 68744 15904 68796 15910
rect 68744 15846 68796 15852
rect 68650 15192 68706 15201
rect 68650 15127 68706 15136
rect 68664 14958 68692 15127
rect 68756 15026 68784 15846
rect 68744 15020 68796 15026
rect 68744 14962 68796 14968
rect 68652 14952 68704 14958
rect 68652 14894 68704 14900
rect 68744 14816 68796 14822
rect 68744 14758 68796 14764
rect 68650 14512 68706 14521
rect 68650 14447 68706 14456
rect 68664 14346 68692 14447
rect 68652 14340 68704 14346
rect 68652 14282 68704 14288
rect 68756 14226 68784 14758
rect 68664 14198 68784 14226
rect 68664 13938 68692 14198
rect 68848 14090 68876 19306
rect 69216 18290 69244 26862
rect 69204 18284 69256 18290
rect 69204 18226 69256 18232
rect 69020 18080 69072 18086
rect 69020 18022 69072 18028
rect 69032 17202 69060 18022
rect 69216 17746 69244 18226
rect 69296 18216 69348 18222
rect 69296 18158 69348 18164
rect 69204 17740 69256 17746
rect 69204 17682 69256 17688
rect 69110 17640 69166 17649
rect 69110 17575 69166 17584
rect 69124 17202 69152 17575
rect 69020 17196 69072 17202
rect 69020 17138 69072 17144
rect 69112 17196 69164 17202
rect 69112 17138 69164 17144
rect 69308 17105 69336 18158
rect 69388 17264 69440 17270
rect 69388 17206 69440 17212
rect 69294 17096 69350 17105
rect 69294 17031 69350 17040
rect 69400 16726 69428 17206
rect 69388 16720 69440 16726
rect 69388 16662 69440 16668
rect 68928 16584 68980 16590
rect 68928 16526 68980 16532
rect 68940 16046 68968 16526
rect 68928 16040 68980 16046
rect 68928 15982 68980 15988
rect 68940 15502 68968 15982
rect 69492 15978 69520 27338
rect 69860 27334 69888 29294
rect 70214 29294 70348 29322
rect 70214 29200 70270 29294
rect 70320 27588 70348 29294
rect 71502 29200 71558 30000
rect 72146 29322 72202 30000
rect 72790 29322 72846 30000
rect 73434 29322 73490 30000
rect 74078 29322 74134 30000
rect 74722 29322 74778 30000
rect 75366 29322 75422 30000
rect 76010 29322 76066 30000
rect 76654 29322 76710 30000
rect 77298 29322 77354 30000
rect 77942 29322 77998 30000
rect 79230 29322 79286 30000
rect 72146 29294 72464 29322
rect 72146 29200 72202 29294
rect 71516 27606 71544 29200
rect 72436 27606 72464 29294
rect 72790 29294 73108 29322
rect 72790 29200 72846 29294
rect 70400 27600 70452 27606
rect 70320 27560 70400 27588
rect 70400 27542 70452 27548
rect 71504 27600 71556 27606
rect 71504 27542 71556 27548
rect 72424 27600 72476 27606
rect 72424 27542 72476 27548
rect 70860 27464 70912 27470
rect 70860 27406 70912 27412
rect 71504 27464 71556 27470
rect 71504 27406 71556 27412
rect 72056 27464 72108 27470
rect 72056 27406 72108 27412
rect 69848 27328 69900 27334
rect 69848 27270 69900 27276
rect 70124 26988 70176 26994
rect 70124 26930 70176 26936
rect 70136 26382 70164 26930
rect 70124 26376 70176 26382
rect 70124 26318 70176 26324
rect 70136 22094 70164 26318
rect 69860 22066 70164 22094
rect 69756 18284 69808 18290
rect 69756 18226 69808 18232
rect 69664 17672 69716 17678
rect 69664 17614 69716 17620
rect 69572 17536 69624 17542
rect 69572 17478 69624 17484
rect 69584 16969 69612 17478
rect 69676 17134 69704 17614
rect 69664 17128 69716 17134
rect 69664 17070 69716 17076
rect 69570 16960 69626 16969
rect 69570 16895 69626 16904
rect 69480 15972 69532 15978
rect 69480 15914 69532 15920
rect 68928 15496 68980 15502
rect 68980 15456 69060 15484
rect 68928 15438 68980 15444
rect 68928 14884 68980 14890
rect 68928 14826 68980 14832
rect 68940 14482 68968 14826
rect 68928 14476 68980 14482
rect 68928 14418 68980 14424
rect 68756 14062 68876 14090
rect 68926 14104 68982 14113
rect 68652 13932 68704 13938
rect 68652 13874 68704 13880
rect 68560 13184 68612 13190
rect 68560 13126 68612 13132
rect 68376 12980 68428 12986
rect 68376 12922 68428 12928
rect 68560 12436 68612 12442
rect 68560 12378 68612 12384
rect 68572 12170 68600 12378
rect 68664 12374 68692 13874
rect 68652 12368 68704 12374
rect 68652 12310 68704 12316
rect 68560 12164 68612 12170
rect 68560 12106 68612 12112
rect 68756 11529 68784 14062
rect 68926 14039 68982 14048
rect 68940 13938 68968 14039
rect 68928 13932 68980 13938
rect 68928 13874 68980 13880
rect 69032 13870 69060 15456
rect 69676 15314 69704 17070
rect 69768 16454 69796 18226
rect 69756 16448 69808 16454
rect 69756 16390 69808 16396
rect 69768 16182 69796 16390
rect 69756 16176 69808 16182
rect 69756 16118 69808 16124
rect 69676 15286 69796 15314
rect 69204 15156 69256 15162
rect 69204 15098 69256 15104
rect 69296 15156 69348 15162
rect 69296 15098 69348 15104
rect 69664 15156 69716 15162
rect 69664 15098 69716 15104
rect 69216 15026 69244 15098
rect 69204 15020 69256 15026
rect 69204 14962 69256 14968
rect 69216 14822 69244 14962
rect 69204 14816 69256 14822
rect 69204 14758 69256 14764
rect 69202 14376 69258 14385
rect 69202 14311 69204 14320
rect 69256 14311 69258 14320
rect 69204 14282 69256 14288
rect 69110 14240 69166 14249
rect 69110 14175 69166 14184
rect 69124 14006 69152 14175
rect 69112 14000 69164 14006
rect 69112 13942 69164 13948
rect 69020 13864 69072 13870
rect 69020 13806 69072 13812
rect 68928 13456 68980 13462
rect 68928 13398 68980 13404
rect 68836 13320 68888 13326
rect 68836 13262 68888 13268
rect 68848 12617 68876 13262
rect 68940 12918 68968 13398
rect 69308 13025 69336 15098
rect 69676 15042 69704 15098
rect 69492 15026 69704 15042
rect 69768 15026 69796 15286
rect 69860 15042 69888 22066
rect 70676 18896 70728 18902
rect 70676 18838 70728 18844
rect 70492 18284 70544 18290
rect 70492 18226 70544 18232
rect 70032 18216 70084 18222
rect 70032 18158 70084 18164
rect 69940 16108 69992 16114
rect 69940 16050 69992 16056
rect 69952 15638 69980 16050
rect 69940 15632 69992 15638
rect 69940 15574 69992 15580
rect 69480 15020 69704 15026
rect 69532 15014 69704 15020
rect 69756 15020 69808 15026
rect 69480 14962 69532 14968
rect 69860 15014 69980 15042
rect 69756 14962 69808 14968
rect 69952 14657 69980 15014
rect 69938 14648 69994 14657
rect 69938 14583 69994 14592
rect 70044 14482 70072 18158
rect 70216 18148 70268 18154
rect 70216 18090 70268 18096
rect 70228 17882 70256 18090
rect 70216 17876 70268 17882
rect 70216 17818 70268 17824
rect 70504 17542 70532 18226
rect 70688 18222 70716 18838
rect 70676 18216 70728 18222
rect 70676 18158 70728 18164
rect 70872 18154 70900 27406
rect 71516 27130 71544 27406
rect 71504 27124 71556 27130
rect 71504 27066 71556 27072
rect 71228 22772 71280 22778
rect 71228 22714 71280 22720
rect 70860 18148 70912 18154
rect 70860 18090 70912 18096
rect 70952 18080 71004 18086
rect 70952 18022 71004 18028
rect 70964 17678 70992 18022
rect 70952 17672 71004 17678
rect 70952 17614 71004 17620
rect 70492 17536 70544 17542
rect 70492 17478 70544 17484
rect 70768 17536 70820 17542
rect 70768 17478 70820 17484
rect 70504 17354 70532 17478
rect 70504 17326 70624 17354
rect 70596 17134 70624 17326
rect 70676 17264 70728 17270
rect 70676 17206 70728 17212
rect 70400 17128 70452 17134
rect 70400 17070 70452 17076
rect 70584 17128 70636 17134
rect 70584 17070 70636 17076
rect 70412 16946 70440 17070
rect 70688 16946 70716 17206
rect 70780 17202 70808 17478
rect 70768 17196 70820 17202
rect 70768 17138 70820 17144
rect 70412 16918 70716 16946
rect 70124 16448 70176 16454
rect 70124 16390 70176 16396
rect 70136 15502 70164 16390
rect 70124 15496 70176 15502
rect 70124 15438 70176 15444
rect 70308 15360 70360 15366
rect 70308 15302 70360 15308
rect 70400 15360 70452 15366
rect 70400 15302 70452 15308
rect 70032 14476 70084 14482
rect 70032 14418 70084 14424
rect 70320 14414 70348 15302
rect 70412 14550 70440 15302
rect 70688 14958 70716 16918
rect 71136 16652 71188 16658
rect 71136 16594 71188 16600
rect 70768 16584 70820 16590
rect 70768 16526 70820 16532
rect 70676 14952 70728 14958
rect 70676 14894 70728 14900
rect 70780 14550 70808 16526
rect 70858 15192 70914 15201
rect 70858 15127 70860 15136
rect 70912 15127 70914 15136
rect 70860 15098 70912 15104
rect 70400 14544 70452 14550
rect 70398 14512 70400 14521
rect 70768 14544 70820 14550
rect 70452 14512 70454 14521
rect 70768 14486 70820 14492
rect 70398 14447 70454 14456
rect 70308 14408 70360 14414
rect 70308 14350 70360 14356
rect 69480 14340 69532 14346
rect 69480 14282 69532 14288
rect 69492 14074 69520 14282
rect 69480 14068 69532 14074
rect 69480 14010 69532 14016
rect 70216 14068 70268 14074
rect 70216 14010 70268 14016
rect 70124 13932 70176 13938
rect 70124 13874 70176 13880
rect 69388 13864 69440 13870
rect 69440 13824 69704 13852
rect 69388 13806 69440 13812
rect 69386 13560 69442 13569
rect 69676 13546 69704 13824
rect 69676 13518 69888 13546
rect 69386 13495 69388 13504
rect 69440 13495 69442 13504
rect 69388 13466 69440 13472
rect 69664 13252 69716 13258
rect 69664 13194 69716 13200
rect 69388 13184 69440 13190
rect 69388 13126 69440 13132
rect 69478 13152 69534 13161
rect 69294 13016 69350 13025
rect 69294 12951 69350 12960
rect 68928 12912 68980 12918
rect 68928 12854 68980 12860
rect 69400 12850 69428 13126
rect 69478 13087 69534 13096
rect 69492 12850 69520 13087
rect 69112 12844 69164 12850
rect 69112 12786 69164 12792
rect 69388 12844 69440 12850
rect 69388 12786 69440 12792
rect 69480 12844 69532 12850
rect 69480 12786 69532 12792
rect 68834 12608 68890 12617
rect 68834 12543 68890 12552
rect 69124 12442 69152 12786
rect 69676 12782 69704 13194
rect 69860 13161 69888 13518
rect 69846 13152 69902 13161
rect 69846 13087 69902 13096
rect 69756 12844 69808 12850
rect 69756 12786 69808 12792
rect 69664 12776 69716 12782
rect 69664 12718 69716 12724
rect 69768 12714 69796 12786
rect 69860 12782 69888 13087
rect 70032 12980 70084 12986
rect 70032 12922 70084 12928
rect 69848 12776 69900 12782
rect 69848 12718 69900 12724
rect 69756 12708 69808 12714
rect 69756 12650 69808 12656
rect 69296 12640 69348 12646
rect 69296 12582 69348 12588
rect 69308 12442 69336 12582
rect 69112 12436 69164 12442
rect 69112 12378 69164 12384
rect 69296 12436 69348 12442
rect 69296 12378 69348 12384
rect 69480 12436 69532 12442
rect 69480 12378 69532 12384
rect 69388 12368 69440 12374
rect 69388 12310 69440 12316
rect 68928 12232 68980 12238
rect 68928 12174 68980 12180
rect 68940 12102 68968 12174
rect 69400 12170 69428 12310
rect 69492 12220 69520 12378
rect 69664 12232 69716 12238
rect 69492 12192 69664 12220
rect 69664 12174 69716 12180
rect 69754 12200 69810 12209
rect 69388 12164 69440 12170
rect 69754 12135 69810 12144
rect 69388 12106 69440 12112
rect 69768 12102 69796 12135
rect 68836 12096 68888 12102
rect 68836 12038 68888 12044
rect 68928 12096 68980 12102
rect 68928 12038 68980 12044
rect 69756 12096 69808 12102
rect 69756 12038 69808 12044
rect 68848 11830 68876 12038
rect 68836 11824 68888 11830
rect 68836 11766 68888 11772
rect 68940 11762 68968 12038
rect 69860 11898 69888 12718
rect 70044 12646 70072 12922
rect 70032 12640 70084 12646
rect 70032 12582 70084 12588
rect 70136 12170 70164 13874
rect 70228 13326 70256 14010
rect 70584 13796 70636 13802
rect 70584 13738 70636 13744
rect 70306 13560 70362 13569
rect 70306 13495 70362 13504
rect 70216 13320 70268 13326
rect 70216 13262 70268 13268
rect 70320 12918 70348 13495
rect 70308 12912 70360 12918
rect 70308 12854 70360 12860
rect 70216 12436 70268 12442
rect 70596 12434 70624 13738
rect 71044 13728 71096 13734
rect 71044 13670 71096 13676
rect 71056 13326 71084 13670
rect 70768 13320 70820 13326
rect 70768 13262 70820 13268
rect 71044 13320 71096 13326
rect 71044 13262 71096 13268
rect 70780 13161 70808 13262
rect 70766 13152 70822 13161
rect 70766 13087 70822 13096
rect 70216 12378 70268 12384
rect 70412 12406 70624 12434
rect 70228 12345 70256 12378
rect 70214 12336 70270 12345
rect 70214 12271 70270 12280
rect 70032 12164 70084 12170
rect 70032 12106 70084 12112
rect 70124 12164 70176 12170
rect 70124 12106 70176 12112
rect 70044 11898 70072 12106
rect 69112 11892 69164 11898
rect 69112 11834 69164 11840
rect 69204 11892 69256 11898
rect 69204 11834 69256 11840
rect 69848 11892 69900 11898
rect 69848 11834 69900 11840
rect 70032 11892 70084 11898
rect 70032 11834 70084 11840
rect 69124 11762 69152 11834
rect 69216 11762 69244 11834
rect 68928 11756 68980 11762
rect 68928 11698 68980 11704
rect 69112 11756 69164 11762
rect 69112 11698 69164 11704
rect 69204 11756 69256 11762
rect 69204 11698 69256 11704
rect 69018 11656 69074 11665
rect 69018 11591 69074 11600
rect 68742 11520 68798 11529
rect 68742 11455 68798 11464
rect 69032 11098 69060 11591
rect 69124 11286 69152 11698
rect 69216 11393 69244 11698
rect 69202 11384 69258 11393
rect 69202 11319 69258 11328
rect 69296 11348 69348 11354
rect 69296 11290 69348 11296
rect 69112 11280 69164 11286
rect 69112 11222 69164 11228
rect 69308 11121 69336 11290
rect 69388 11280 69440 11286
rect 69386 11248 69388 11257
rect 69440 11248 69442 11257
rect 69386 11183 69442 11192
rect 69294 11112 69350 11121
rect 69032 11082 69152 11098
rect 69032 11076 69164 11082
rect 69032 11070 69112 11076
rect 69294 11047 69350 11056
rect 69112 11018 69164 11024
rect 69020 9988 69072 9994
rect 69020 9930 69072 9936
rect 68284 9376 68336 9382
rect 68284 9318 68336 9324
rect 68192 9172 68244 9178
rect 68192 9114 68244 9120
rect 67548 9036 67600 9042
rect 67548 8978 67600 8984
rect 66794 8732 67102 8741
rect 66794 8730 66800 8732
rect 66856 8730 66880 8732
rect 66936 8730 66960 8732
rect 67016 8730 67040 8732
rect 67096 8730 67102 8732
rect 66856 8678 66858 8730
rect 67038 8678 67040 8730
rect 66794 8676 66800 8678
rect 66856 8676 66880 8678
rect 66936 8676 66960 8678
rect 67016 8676 67040 8678
rect 67096 8676 67102 8678
rect 66794 8667 67102 8676
rect 67560 8566 67588 8978
rect 68296 8974 68324 9318
rect 68284 8968 68336 8974
rect 68284 8910 68336 8916
rect 67548 8560 67600 8566
rect 67548 8502 67600 8508
rect 66794 7644 67102 7653
rect 66794 7642 66800 7644
rect 66856 7642 66880 7644
rect 66936 7642 66960 7644
rect 67016 7642 67040 7644
rect 67096 7642 67102 7644
rect 66856 7590 66858 7642
rect 67038 7590 67040 7642
rect 66794 7588 66800 7590
rect 66856 7588 66880 7590
rect 66936 7588 66960 7590
rect 67016 7588 67040 7590
rect 67096 7588 67102 7590
rect 66794 7579 67102 7588
rect 66794 6556 67102 6565
rect 66794 6554 66800 6556
rect 66856 6554 66880 6556
rect 66936 6554 66960 6556
rect 67016 6554 67040 6556
rect 67096 6554 67102 6556
rect 66856 6502 66858 6554
rect 67038 6502 67040 6554
rect 66794 6500 66800 6502
rect 66856 6500 66880 6502
rect 66936 6500 66960 6502
rect 67016 6500 67040 6502
rect 67096 6500 67102 6502
rect 66794 6491 67102 6500
rect 66794 5468 67102 5477
rect 66794 5466 66800 5468
rect 66856 5466 66880 5468
rect 66936 5466 66960 5468
rect 67016 5466 67040 5468
rect 67096 5466 67102 5468
rect 66856 5414 66858 5466
rect 67038 5414 67040 5466
rect 66794 5412 66800 5414
rect 66856 5412 66880 5414
rect 66936 5412 66960 5414
rect 67016 5412 67040 5414
rect 67096 5412 67102 5414
rect 66794 5403 67102 5412
rect 66794 4380 67102 4389
rect 66794 4378 66800 4380
rect 66856 4378 66880 4380
rect 66936 4378 66960 4380
rect 67016 4378 67040 4380
rect 67096 4378 67102 4380
rect 66856 4326 66858 4378
rect 67038 4326 67040 4378
rect 66794 4324 66800 4326
rect 66856 4324 66880 4326
rect 66936 4324 66960 4326
rect 67016 4324 67040 4326
rect 67096 4324 67102 4326
rect 66794 4315 67102 4324
rect 66794 3292 67102 3301
rect 66794 3290 66800 3292
rect 66856 3290 66880 3292
rect 66936 3290 66960 3292
rect 67016 3290 67040 3292
rect 67096 3290 67102 3292
rect 66856 3238 66858 3290
rect 67038 3238 67040 3290
rect 66794 3236 66800 3238
rect 66856 3236 66880 3238
rect 66936 3236 66960 3238
rect 67016 3236 67040 3238
rect 67096 3236 67102 3238
rect 66794 3227 67102 3236
rect 67456 2848 67508 2854
rect 67456 2790 67508 2796
rect 68376 2848 68428 2854
rect 68376 2790 68428 2796
rect 67468 2446 67496 2790
rect 68388 2446 68416 2790
rect 69032 2650 69060 9930
rect 70228 3534 70256 12271
rect 70308 12232 70360 12238
rect 70412 12220 70440 12406
rect 70780 12306 70808 13087
rect 70768 12300 70820 12306
rect 70768 12242 70820 12248
rect 70360 12192 70440 12220
rect 70308 12174 70360 12180
rect 70412 11558 70440 12192
rect 70860 11824 70912 11830
rect 70858 11792 70860 11801
rect 70912 11792 70914 11801
rect 70858 11727 70914 11736
rect 70400 11552 70452 11558
rect 70400 11494 70452 11500
rect 70768 8832 70820 8838
rect 70768 8774 70820 8780
rect 70676 5024 70728 5030
rect 70676 4966 70728 4972
rect 70688 4214 70716 4966
rect 70676 4208 70728 4214
rect 70676 4150 70728 4156
rect 70216 3528 70268 3534
rect 70216 3470 70268 3476
rect 70780 2650 70808 8774
rect 71148 4622 71176 16594
rect 71240 15570 71268 22714
rect 72068 22094 72096 27406
rect 72516 27328 72568 27334
rect 72516 27270 72568 27276
rect 71976 22066 72096 22094
rect 71976 18698 72004 22066
rect 71964 18692 72016 18698
rect 71964 18634 72016 18640
rect 71320 17128 71372 17134
rect 71320 17070 71372 17076
rect 71332 16590 71360 17070
rect 71320 16584 71372 16590
rect 71320 16526 71372 16532
rect 72424 16244 72476 16250
rect 72424 16186 72476 16192
rect 71872 16108 71924 16114
rect 71872 16050 71924 16056
rect 71504 16040 71556 16046
rect 71504 15982 71556 15988
rect 71516 15570 71544 15982
rect 71884 15706 71912 16050
rect 72056 15904 72108 15910
rect 72056 15846 72108 15852
rect 71872 15700 71924 15706
rect 71872 15642 71924 15648
rect 71228 15564 71280 15570
rect 71228 15506 71280 15512
rect 71504 15564 71556 15570
rect 71504 15506 71556 15512
rect 71228 14816 71280 14822
rect 71228 14758 71280 14764
rect 71240 13870 71268 14758
rect 71228 13864 71280 13870
rect 71228 13806 71280 13812
rect 71320 13796 71372 13802
rect 71320 13738 71372 13744
rect 71332 12434 71360 13738
rect 71240 12406 71360 12434
rect 71240 5030 71268 12406
rect 71320 12232 71372 12238
rect 71320 12174 71372 12180
rect 71332 11898 71360 12174
rect 71320 11892 71372 11898
rect 71320 11834 71372 11840
rect 71516 11762 71544 15506
rect 72068 15502 72096 15846
rect 72436 15502 72464 16186
rect 72056 15496 72108 15502
rect 72056 15438 72108 15444
rect 72424 15496 72476 15502
rect 72424 15438 72476 15444
rect 71964 15088 72016 15094
rect 71964 15030 72016 15036
rect 71780 14068 71832 14074
rect 71780 14010 71832 14016
rect 71686 13016 71742 13025
rect 71686 12951 71742 12960
rect 71700 12850 71728 12951
rect 71688 12844 71740 12850
rect 71688 12786 71740 12792
rect 71792 12646 71820 14010
rect 71976 13938 72004 15030
rect 72056 14816 72108 14822
rect 72056 14758 72108 14764
rect 72068 14346 72096 14758
rect 72056 14340 72108 14346
rect 72056 14282 72108 14288
rect 71872 13932 71924 13938
rect 71872 13874 71924 13880
rect 71964 13932 72016 13938
rect 71964 13874 72016 13880
rect 72240 13932 72292 13938
rect 72240 13874 72292 13880
rect 72332 13932 72384 13938
rect 72332 13874 72384 13880
rect 71884 13462 71912 13874
rect 71872 13456 71924 13462
rect 71872 13398 71924 13404
rect 72252 13258 72280 13874
rect 72344 13530 72372 13874
rect 72332 13524 72384 13530
rect 72332 13466 72384 13472
rect 72240 13252 72292 13258
rect 72240 13194 72292 13200
rect 72528 13190 72556 27270
rect 73080 27146 73108 29294
rect 73434 29294 73752 29322
rect 73434 29200 73490 29294
rect 73724 27470 73752 29294
rect 74078 29294 74304 29322
rect 74078 29200 74134 29294
rect 74276 27606 74304 29294
rect 74722 29294 74856 29322
rect 74722 29200 74778 29294
rect 74828 27606 74856 29294
rect 75366 29294 75500 29322
rect 75366 29200 75422 29294
rect 74264 27600 74316 27606
rect 74264 27542 74316 27548
rect 74816 27600 74868 27606
rect 74816 27542 74868 27548
rect 73712 27464 73764 27470
rect 73712 27406 73764 27412
rect 74448 27464 74500 27470
rect 74448 27406 74500 27412
rect 73804 27328 73856 27334
rect 73804 27270 73856 27276
rect 73080 27130 73200 27146
rect 73080 27124 73212 27130
rect 73080 27118 73160 27124
rect 73160 27066 73212 27072
rect 73528 26988 73580 26994
rect 73528 26930 73580 26936
rect 73436 22636 73488 22642
rect 73436 22578 73488 22584
rect 73068 16652 73120 16658
rect 73068 16594 73120 16600
rect 73080 16182 73108 16594
rect 73068 16176 73120 16182
rect 73068 16118 73120 16124
rect 73448 14550 73476 22578
rect 73540 18766 73568 26930
rect 73528 18760 73580 18766
rect 73528 18702 73580 18708
rect 73436 14544 73488 14550
rect 73436 14486 73488 14492
rect 73712 14272 73764 14278
rect 73712 14214 73764 14220
rect 73724 13938 73752 14214
rect 73712 13932 73764 13938
rect 73712 13874 73764 13880
rect 72516 13184 72568 13190
rect 72516 13126 72568 13132
rect 71872 12844 71924 12850
rect 71872 12786 71924 12792
rect 72332 12844 72384 12850
rect 72332 12786 72384 12792
rect 71780 12640 71832 12646
rect 71780 12582 71832 12588
rect 71504 11756 71556 11762
rect 71504 11698 71556 11704
rect 71412 11688 71464 11694
rect 71412 11630 71464 11636
rect 71228 5024 71280 5030
rect 71228 4966 71280 4972
rect 71136 4616 71188 4622
rect 71136 4558 71188 4564
rect 71148 4078 71176 4558
rect 71136 4072 71188 4078
rect 71136 4014 71188 4020
rect 71424 2650 71452 11630
rect 71884 8242 71912 12786
rect 72344 12374 72372 12786
rect 72424 12640 72476 12646
rect 72422 12608 72424 12617
rect 72476 12608 72478 12617
rect 72422 12543 72478 12552
rect 72332 12368 72384 12374
rect 72332 12310 72384 12316
rect 72344 11898 72372 12310
rect 72332 11892 72384 11898
rect 72332 11834 72384 11840
rect 73816 11354 73844 27270
rect 73896 26988 73948 26994
rect 73896 26930 73948 26936
rect 73908 14074 73936 26930
rect 74460 23526 74488 27406
rect 75092 27396 75144 27402
rect 75092 27338 75144 27344
rect 75104 27130 75132 27338
rect 75184 27328 75236 27334
rect 75184 27270 75236 27276
rect 75092 27124 75144 27130
rect 75092 27066 75144 27072
rect 73988 23520 74040 23526
rect 73988 23462 74040 23468
rect 74448 23520 74500 23526
rect 74448 23462 74500 23468
rect 73896 14068 73948 14074
rect 73896 14010 73948 14016
rect 73804 11348 73856 11354
rect 73804 11290 73856 11296
rect 74000 11286 74028 23462
rect 75196 17610 75224 27270
rect 75472 27130 75500 29294
rect 76010 29294 76328 29322
rect 76010 29200 76066 29294
rect 76300 27470 76328 29294
rect 76654 29294 76880 29322
rect 76654 29200 76710 29294
rect 76852 27606 76880 29294
rect 77298 29294 77432 29322
rect 77298 29200 77354 29294
rect 77404 27606 77432 29294
rect 77942 29294 78352 29322
rect 77942 29200 77998 29294
rect 77768 27772 78076 27781
rect 77768 27770 77774 27772
rect 77830 27770 77854 27772
rect 77910 27770 77934 27772
rect 77990 27770 78014 27772
rect 78070 27770 78076 27772
rect 77830 27718 77832 27770
rect 78012 27718 78014 27770
rect 77768 27716 77774 27718
rect 77830 27716 77854 27718
rect 77910 27716 77934 27718
rect 77990 27716 78014 27718
rect 78070 27716 78076 27718
rect 77768 27707 78076 27716
rect 76840 27600 76892 27606
rect 76840 27542 76892 27548
rect 77392 27600 77444 27606
rect 77392 27542 77444 27548
rect 78324 27470 78352 29294
rect 79230 29294 79456 29322
rect 79230 29200 79286 29294
rect 79428 27470 79456 29294
rect 79874 29200 79930 30000
rect 80518 29200 80574 30000
rect 81162 29322 81218 30000
rect 81806 29322 81862 30000
rect 82450 29322 82506 30000
rect 81162 29294 81388 29322
rect 81162 29200 81218 29294
rect 76288 27464 76340 27470
rect 76288 27406 76340 27412
rect 76380 27464 76432 27470
rect 76380 27406 76432 27412
rect 78312 27464 78364 27470
rect 78312 27406 78364 27412
rect 79416 27464 79468 27470
rect 79888 27452 79916 29200
rect 80060 27464 80112 27470
rect 79888 27424 80060 27452
rect 79416 27406 79468 27412
rect 81360 27452 81388 29294
rect 81806 29294 82032 29322
rect 81806 29200 81862 29294
rect 82004 27606 82032 29294
rect 82450 29294 82584 29322
rect 82450 29200 82506 29294
rect 81992 27600 82044 27606
rect 81992 27542 82044 27548
rect 82556 27470 82584 29294
rect 83094 29200 83150 30000
rect 83738 29322 83794 30000
rect 83738 29294 84148 29322
rect 83738 29200 83794 29294
rect 83108 27606 83136 29200
rect 83096 27600 83148 27606
rect 83096 27542 83148 27548
rect 83740 27600 83792 27606
rect 83740 27542 83792 27548
rect 84120 27554 84148 29294
rect 84382 29200 84438 30000
rect 85026 29322 85082 30000
rect 85026 29294 85160 29322
rect 85026 29200 85082 29294
rect 81440 27464 81492 27470
rect 81360 27424 81440 27452
rect 80060 27406 80112 27412
rect 81440 27406 81492 27412
rect 82176 27464 82228 27470
rect 82176 27406 82228 27412
rect 82544 27464 82596 27470
rect 82544 27406 82596 27412
rect 75460 27124 75512 27130
rect 75460 27066 75512 27072
rect 75644 26988 75696 26994
rect 75644 26930 75696 26936
rect 75656 26790 75684 26930
rect 75644 26784 75696 26790
rect 75644 26726 75696 26732
rect 76392 18426 76420 27406
rect 78128 27396 78180 27402
rect 78128 27338 78180 27344
rect 76748 26920 76800 26926
rect 76748 26862 76800 26868
rect 76380 18420 76432 18426
rect 76380 18362 76432 18368
rect 75184 17604 75236 17610
rect 75184 17546 75236 17552
rect 74816 14884 74868 14890
rect 74816 14826 74868 14832
rect 74828 14414 74856 14826
rect 74816 14408 74868 14414
rect 74816 14350 74868 14356
rect 73988 11280 74040 11286
rect 73988 11222 74040 11228
rect 71884 8214 72648 8242
rect 72620 4078 72648 8214
rect 72608 4072 72660 4078
rect 72608 4014 72660 4020
rect 71596 3936 71648 3942
rect 71596 3878 71648 3884
rect 71608 3058 71636 3878
rect 76760 3670 76788 26862
rect 77768 26684 78076 26693
rect 77768 26682 77774 26684
rect 77830 26682 77854 26684
rect 77910 26682 77934 26684
rect 77990 26682 78014 26684
rect 78070 26682 78076 26684
rect 77830 26630 77832 26682
rect 78012 26630 78014 26682
rect 77768 26628 77774 26630
rect 77830 26628 77854 26630
rect 77910 26628 77934 26630
rect 77990 26628 78014 26630
rect 78070 26628 78076 26630
rect 77768 26619 78076 26628
rect 77768 25596 78076 25605
rect 77768 25594 77774 25596
rect 77830 25594 77854 25596
rect 77910 25594 77934 25596
rect 77990 25594 78014 25596
rect 78070 25594 78076 25596
rect 77830 25542 77832 25594
rect 78012 25542 78014 25594
rect 77768 25540 77774 25542
rect 77830 25540 77854 25542
rect 77910 25540 77934 25542
rect 77990 25540 78014 25542
rect 78070 25540 78076 25542
rect 77768 25531 78076 25540
rect 77768 24508 78076 24517
rect 77768 24506 77774 24508
rect 77830 24506 77854 24508
rect 77910 24506 77934 24508
rect 77990 24506 78014 24508
rect 78070 24506 78076 24508
rect 77830 24454 77832 24506
rect 78012 24454 78014 24506
rect 77768 24452 77774 24454
rect 77830 24452 77854 24454
rect 77910 24452 77934 24454
rect 77990 24452 78014 24454
rect 78070 24452 78076 24454
rect 77768 24443 78076 24452
rect 77768 23420 78076 23429
rect 77768 23418 77774 23420
rect 77830 23418 77854 23420
rect 77910 23418 77934 23420
rect 77990 23418 78014 23420
rect 78070 23418 78076 23420
rect 77830 23366 77832 23418
rect 78012 23366 78014 23418
rect 77768 23364 77774 23366
rect 77830 23364 77854 23366
rect 77910 23364 77934 23366
rect 77990 23364 78014 23366
rect 78070 23364 78076 23366
rect 77768 23355 78076 23364
rect 77768 22332 78076 22341
rect 77768 22330 77774 22332
rect 77830 22330 77854 22332
rect 77910 22330 77934 22332
rect 77990 22330 78014 22332
rect 78070 22330 78076 22332
rect 77830 22278 77832 22330
rect 78012 22278 78014 22330
rect 77768 22276 77774 22278
rect 77830 22276 77854 22278
rect 77910 22276 77934 22278
rect 77990 22276 78014 22278
rect 78070 22276 78076 22278
rect 77768 22267 78076 22276
rect 77768 21244 78076 21253
rect 77768 21242 77774 21244
rect 77830 21242 77854 21244
rect 77910 21242 77934 21244
rect 77990 21242 78014 21244
rect 78070 21242 78076 21244
rect 77830 21190 77832 21242
rect 78012 21190 78014 21242
rect 77768 21188 77774 21190
rect 77830 21188 77854 21190
rect 77910 21188 77934 21190
rect 77990 21188 78014 21190
rect 78070 21188 78076 21190
rect 77768 21179 78076 21188
rect 77768 20156 78076 20165
rect 77768 20154 77774 20156
rect 77830 20154 77854 20156
rect 77910 20154 77934 20156
rect 77990 20154 78014 20156
rect 78070 20154 78076 20156
rect 77830 20102 77832 20154
rect 78012 20102 78014 20154
rect 77768 20100 77774 20102
rect 77830 20100 77854 20102
rect 77910 20100 77934 20102
rect 77990 20100 78014 20102
rect 78070 20100 78076 20102
rect 77768 20091 78076 20100
rect 77768 19068 78076 19077
rect 77768 19066 77774 19068
rect 77830 19066 77854 19068
rect 77910 19066 77934 19068
rect 77990 19066 78014 19068
rect 78070 19066 78076 19068
rect 77830 19014 77832 19066
rect 78012 19014 78014 19066
rect 77768 19012 77774 19014
rect 77830 19012 77854 19014
rect 77910 19012 77934 19014
rect 77990 19012 78014 19014
rect 78070 19012 78076 19014
rect 77768 19003 78076 19012
rect 78140 18358 78168 27338
rect 78956 27328 79008 27334
rect 78956 27270 79008 27276
rect 79600 27328 79652 27334
rect 79600 27270 79652 27276
rect 80244 27328 80296 27334
rect 80244 27270 80296 27276
rect 81532 27328 81584 27334
rect 81532 27270 81584 27276
rect 78968 18630 78996 27270
rect 78956 18624 79008 18630
rect 78956 18566 79008 18572
rect 78128 18352 78180 18358
rect 78128 18294 78180 18300
rect 77768 17980 78076 17989
rect 77768 17978 77774 17980
rect 77830 17978 77854 17980
rect 77910 17978 77934 17980
rect 77990 17978 78014 17980
rect 78070 17978 78076 17980
rect 77830 17926 77832 17978
rect 78012 17926 78014 17978
rect 77768 17924 77774 17926
rect 77830 17924 77854 17926
rect 77910 17924 77934 17926
rect 77990 17924 78014 17926
rect 78070 17924 78076 17926
rect 77768 17915 78076 17924
rect 77768 16892 78076 16901
rect 77768 16890 77774 16892
rect 77830 16890 77854 16892
rect 77910 16890 77934 16892
rect 77990 16890 78014 16892
rect 78070 16890 78076 16892
rect 77830 16838 77832 16890
rect 78012 16838 78014 16890
rect 77768 16836 77774 16838
rect 77830 16836 77854 16838
rect 77910 16836 77934 16838
rect 77990 16836 78014 16838
rect 78070 16836 78076 16838
rect 77768 16827 78076 16836
rect 77116 16720 77168 16726
rect 77116 16662 77168 16668
rect 76748 3664 76800 3670
rect 76748 3606 76800 3612
rect 73528 3596 73580 3602
rect 73528 3538 73580 3544
rect 71596 3052 71648 3058
rect 71596 2994 71648 3000
rect 71504 2848 71556 2854
rect 71504 2790 71556 2796
rect 69020 2644 69072 2650
rect 69020 2586 69072 2592
rect 70768 2644 70820 2650
rect 70768 2586 70820 2592
rect 71412 2644 71464 2650
rect 71412 2586 71464 2592
rect 68928 2576 68980 2582
rect 68848 2524 68928 2530
rect 68848 2518 68980 2524
rect 68848 2502 68968 2518
rect 68848 2446 68876 2502
rect 66260 2440 66312 2446
rect 66260 2382 66312 2388
rect 66444 2440 66496 2446
rect 66444 2382 66496 2388
rect 67456 2440 67508 2446
rect 67456 2382 67508 2388
rect 68376 2440 68428 2446
rect 68376 2382 68428 2388
rect 68836 2440 68888 2446
rect 68836 2382 68888 2388
rect 68928 2440 68980 2446
rect 68928 2382 68980 2388
rect 70216 2440 70268 2446
rect 70216 2382 70268 2388
rect 65064 2304 65116 2310
rect 65064 2246 65116 2252
rect 65708 2304 65760 2310
rect 65708 2246 65760 2252
rect 64696 2100 64748 2106
rect 64696 2042 64748 2048
rect 65076 800 65104 2246
rect 65720 800 65748 2246
rect 66456 1306 66484 2382
rect 66720 2304 66772 2310
rect 66720 2246 66772 2252
rect 67180 2304 67232 2310
rect 67180 2246 67232 2252
rect 67640 2304 67692 2310
rect 67640 2246 67692 2252
rect 66732 1970 66760 2246
rect 66794 2204 67102 2213
rect 66794 2202 66800 2204
rect 66856 2202 66880 2204
rect 66936 2202 66960 2204
rect 67016 2202 67040 2204
rect 67096 2202 67102 2204
rect 66856 2150 66858 2202
rect 67038 2150 67040 2202
rect 66794 2148 66800 2150
rect 66856 2148 66880 2150
rect 66936 2148 66960 2150
rect 67016 2148 67040 2150
rect 67096 2148 67102 2150
rect 66794 2139 67102 2148
rect 66720 1964 66772 1970
rect 66720 1906 66772 1912
rect 66364 1278 66484 1306
rect 66364 800 66392 1278
rect 67192 1170 67220 2246
rect 67008 1142 67220 1170
rect 67008 800 67036 1142
rect 67652 800 67680 2246
rect 68940 800 68968 2382
rect 69572 2304 69624 2310
rect 69572 2246 69624 2252
rect 69584 800 69612 2246
rect 70228 800 70256 2382
rect 70860 2372 70912 2378
rect 70860 2314 70912 2320
rect 70872 800 70900 2314
rect 71516 800 71544 2790
rect 71596 2644 71648 2650
rect 71596 2586 71648 2592
rect 71608 1494 71636 2586
rect 73540 2446 73568 3538
rect 75184 3528 75236 3534
rect 75184 3470 75236 3476
rect 75196 3194 75224 3470
rect 75184 3188 75236 3194
rect 75184 3130 75236 3136
rect 76760 3126 76788 3606
rect 77128 3126 77156 16662
rect 77768 15804 78076 15813
rect 77768 15802 77774 15804
rect 77830 15802 77854 15804
rect 77910 15802 77934 15804
rect 77990 15802 78014 15804
rect 78070 15802 78076 15804
rect 77830 15750 77832 15802
rect 78012 15750 78014 15802
rect 77768 15748 77774 15750
rect 77830 15748 77854 15750
rect 77910 15748 77934 15750
rect 77990 15748 78014 15750
rect 78070 15748 78076 15750
rect 77768 15739 78076 15748
rect 77768 14716 78076 14725
rect 77768 14714 77774 14716
rect 77830 14714 77854 14716
rect 77910 14714 77934 14716
rect 77990 14714 78014 14716
rect 78070 14714 78076 14716
rect 77830 14662 77832 14714
rect 78012 14662 78014 14714
rect 77768 14660 77774 14662
rect 77830 14660 77854 14662
rect 77910 14660 77934 14662
rect 77990 14660 78014 14662
rect 78070 14660 78076 14662
rect 77768 14651 78076 14660
rect 77768 13628 78076 13637
rect 77768 13626 77774 13628
rect 77830 13626 77854 13628
rect 77910 13626 77934 13628
rect 77990 13626 78014 13628
rect 78070 13626 78076 13628
rect 77830 13574 77832 13626
rect 78012 13574 78014 13626
rect 77768 13572 77774 13574
rect 77830 13572 77854 13574
rect 77910 13572 77934 13574
rect 77990 13572 78014 13574
rect 78070 13572 78076 13574
rect 77768 13563 78076 13572
rect 79612 13433 79640 27270
rect 80256 24177 80284 27270
rect 81544 27062 81572 27270
rect 81532 27056 81584 27062
rect 81532 26998 81584 27004
rect 80242 24168 80298 24177
rect 80242 24103 80298 24112
rect 79598 13424 79654 13433
rect 79598 13359 79654 13368
rect 77768 12540 78076 12549
rect 77768 12538 77774 12540
rect 77830 12538 77854 12540
rect 77910 12538 77934 12540
rect 77990 12538 78014 12540
rect 78070 12538 78076 12540
rect 77830 12486 77832 12538
rect 78012 12486 78014 12538
rect 77768 12484 77774 12486
rect 77830 12484 77854 12486
rect 77910 12484 77934 12486
rect 77990 12484 78014 12486
rect 78070 12484 78076 12486
rect 77768 12475 78076 12484
rect 82188 12442 82216 27406
rect 82728 27328 82780 27334
rect 82728 27270 82780 27276
rect 82740 26450 82768 27270
rect 82728 26444 82780 26450
rect 82728 26386 82780 26392
rect 83752 19990 83780 27542
rect 84120 27526 84240 27554
rect 84212 27470 84240 27526
rect 83832 27464 83884 27470
rect 83832 27406 83884 27412
rect 84200 27464 84252 27470
rect 84200 27406 84252 27412
rect 83844 27130 83872 27406
rect 83832 27124 83884 27130
rect 83832 27066 83884 27072
rect 84396 26994 84424 29200
rect 85132 27470 85160 29294
rect 85670 29200 85726 30000
rect 86314 29336 86370 29345
rect 86314 29271 86370 29280
rect 85684 27606 85712 29200
rect 85672 27600 85724 27606
rect 85672 27542 85724 27548
rect 86132 27532 86184 27538
rect 86132 27474 86184 27480
rect 85120 27464 85172 27470
rect 85120 27406 85172 27412
rect 84384 26988 84436 26994
rect 84384 26930 84436 26936
rect 85120 26988 85172 26994
rect 85120 26930 85172 26936
rect 85132 26382 85160 26930
rect 85396 26784 85448 26790
rect 85396 26726 85448 26732
rect 85408 26450 85436 26726
rect 85396 26444 85448 26450
rect 85396 26386 85448 26392
rect 85120 26376 85172 26382
rect 85120 26318 85172 26324
rect 84844 21004 84896 21010
rect 84844 20946 84896 20952
rect 83740 19984 83792 19990
rect 83740 19926 83792 19932
rect 82820 14476 82872 14482
rect 82820 14418 82872 14424
rect 82176 12436 82228 12442
rect 82176 12378 82228 12384
rect 77768 11452 78076 11461
rect 77768 11450 77774 11452
rect 77830 11450 77854 11452
rect 77910 11450 77934 11452
rect 77990 11450 78014 11452
rect 78070 11450 78076 11452
rect 77830 11398 77832 11450
rect 78012 11398 78014 11450
rect 77768 11396 77774 11398
rect 77830 11396 77854 11398
rect 77910 11396 77934 11398
rect 77990 11396 78014 11398
rect 78070 11396 78076 11398
rect 77768 11387 78076 11396
rect 77768 10364 78076 10373
rect 77768 10362 77774 10364
rect 77830 10362 77854 10364
rect 77910 10362 77934 10364
rect 77990 10362 78014 10364
rect 78070 10362 78076 10364
rect 77830 10310 77832 10362
rect 78012 10310 78014 10362
rect 77768 10308 77774 10310
rect 77830 10308 77854 10310
rect 77910 10308 77934 10310
rect 77990 10308 78014 10310
rect 78070 10308 78076 10310
rect 77768 10299 78076 10308
rect 77768 9276 78076 9285
rect 77768 9274 77774 9276
rect 77830 9274 77854 9276
rect 77910 9274 77934 9276
rect 77990 9274 78014 9276
rect 78070 9274 78076 9276
rect 77830 9222 77832 9274
rect 78012 9222 78014 9274
rect 77768 9220 77774 9222
rect 77830 9220 77854 9222
rect 77910 9220 77934 9222
rect 77990 9220 78014 9222
rect 78070 9220 78076 9222
rect 77768 9211 78076 9220
rect 82832 8362 82860 14418
rect 84856 14414 84884 20946
rect 84844 14408 84896 14414
rect 84844 14350 84896 14356
rect 82820 8356 82872 8362
rect 82820 8298 82872 8304
rect 77768 8188 78076 8197
rect 77768 8186 77774 8188
rect 77830 8186 77854 8188
rect 77910 8186 77934 8188
rect 77990 8186 78014 8188
rect 78070 8186 78076 8188
rect 77830 8134 77832 8186
rect 78012 8134 78014 8186
rect 77768 8132 77774 8134
rect 77830 8132 77854 8134
rect 77910 8132 77934 8134
rect 77990 8132 78014 8134
rect 78070 8132 78076 8134
rect 77768 8123 78076 8132
rect 77768 7100 78076 7109
rect 77768 7098 77774 7100
rect 77830 7098 77854 7100
rect 77910 7098 77934 7100
rect 77990 7098 78014 7100
rect 78070 7098 78076 7100
rect 77830 7046 77832 7098
rect 78012 7046 78014 7098
rect 77768 7044 77774 7046
rect 77830 7044 77854 7046
rect 77910 7044 77934 7046
rect 77990 7044 78014 7046
rect 78070 7044 78076 7046
rect 77768 7035 78076 7044
rect 77768 6012 78076 6021
rect 77768 6010 77774 6012
rect 77830 6010 77854 6012
rect 77910 6010 77934 6012
rect 77990 6010 78014 6012
rect 78070 6010 78076 6012
rect 77830 5958 77832 6010
rect 78012 5958 78014 6010
rect 77768 5956 77774 5958
rect 77830 5956 77854 5958
rect 77910 5956 77934 5958
rect 77990 5956 78014 5958
rect 78070 5956 78076 5958
rect 77768 5947 78076 5956
rect 77768 4924 78076 4933
rect 77768 4922 77774 4924
rect 77830 4922 77854 4924
rect 77910 4922 77934 4924
rect 77990 4922 78014 4924
rect 78070 4922 78076 4924
rect 77830 4870 77832 4922
rect 78012 4870 78014 4922
rect 77768 4868 77774 4870
rect 77830 4868 77854 4870
rect 77910 4868 77934 4870
rect 77990 4868 78014 4870
rect 78070 4868 78076 4870
rect 77768 4859 78076 4868
rect 83832 4820 83884 4826
rect 83832 4762 83884 4768
rect 81532 4004 81584 4010
rect 81532 3946 81584 3952
rect 77768 3836 78076 3845
rect 77768 3834 77774 3836
rect 77830 3834 77854 3836
rect 77910 3834 77934 3836
rect 77990 3834 78014 3836
rect 78070 3834 78076 3836
rect 77830 3782 77832 3834
rect 78012 3782 78014 3834
rect 77768 3780 77774 3782
rect 77830 3780 77854 3782
rect 77910 3780 77934 3782
rect 77990 3780 78014 3782
rect 78070 3780 78076 3782
rect 77768 3771 78076 3780
rect 76748 3120 76800 3126
rect 76748 3062 76800 3068
rect 77116 3120 77168 3126
rect 77116 3062 77168 3068
rect 79692 3120 79744 3126
rect 79692 3062 79744 3068
rect 76760 2990 76788 3062
rect 76748 2984 76800 2990
rect 76748 2926 76800 2932
rect 77768 2748 78076 2757
rect 77768 2746 77774 2748
rect 77830 2746 77854 2748
rect 77910 2746 77934 2748
rect 77990 2746 78014 2748
rect 78070 2746 78076 2748
rect 77830 2694 77832 2746
rect 78012 2694 78014 2746
rect 77768 2692 77774 2694
rect 77830 2692 77854 2694
rect 77910 2692 77934 2694
rect 77990 2692 78014 2694
rect 78070 2692 78076 2694
rect 77768 2683 78076 2692
rect 78588 2576 78640 2582
rect 78588 2518 78640 2524
rect 79232 2576 79284 2582
rect 79232 2518 79284 2524
rect 72148 2440 72200 2446
rect 72148 2382 72200 2388
rect 73528 2440 73580 2446
rect 73528 2382 73580 2388
rect 74080 2440 74132 2446
rect 74080 2382 74132 2388
rect 76748 2440 76800 2446
rect 76748 2382 76800 2388
rect 77024 2440 77076 2446
rect 77024 2382 77076 2388
rect 71596 1488 71648 1494
rect 71596 1430 71648 1436
rect 72160 800 72188 2382
rect 72424 2304 72476 2310
rect 72424 2246 72476 2252
rect 72792 2304 72844 2310
rect 72792 2246 72844 2252
rect 72436 1562 72464 2246
rect 72424 1556 72476 1562
rect 72424 1498 72476 1504
rect 72804 800 72832 2246
rect 74092 800 74120 2382
rect 74724 2372 74776 2378
rect 74724 2314 74776 2320
rect 74736 800 74764 2314
rect 75368 2304 75420 2310
rect 75368 2246 75420 2252
rect 76656 2304 76708 2310
rect 76656 2246 76708 2252
rect 75380 800 75408 2246
rect 76668 800 76696 2246
rect 76760 1902 76788 2382
rect 77036 2310 77064 2382
rect 77944 2372 77996 2378
rect 77944 2314 77996 2320
rect 77024 2304 77076 2310
rect 77024 2246 77076 2252
rect 77300 2304 77352 2310
rect 77300 2246 77352 2252
rect 76748 1896 76800 1902
rect 76748 1838 76800 1844
rect 77036 1494 77064 2246
rect 77024 1488 77076 1494
rect 77024 1430 77076 1436
rect 77312 800 77340 2246
rect 77956 800 77984 2314
rect 78600 800 78628 2518
rect 79244 800 79272 2518
rect 79508 2440 79560 2446
rect 79508 2382 79560 2388
rect 79520 1698 79548 2382
rect 79704 2378 79732 3062
rect 81544 3058 81572 3946
rect 81532 3052 81584 3058
rect 81532 2994 81584 3000
rect 79968 2848 80020 2854
rect 79968 2790 80020 2796
rect 81808 2848 81860 2854
rect 81808 2790 81860 2796
rect 79980 2446 80008 2790
rect 80796 2576 80848 2582
rect 80794 2544 80796 2553
rect 81164 2576 81216 2582
rect 80848 2544 80850 2553
rect 81164 2518 81216 2524
rect 80794 2479 80850 2488
rect 79968 2440 80020 2446
rect 79968 2382 80020 2388
rect 80520 2440 80572 2446
rect 80520 2382 80572 2388
rect 79692 2372 79744 2378
rect 79692 2314 79744 2320
rect 80060 2304 80112 2310
rect 79888 2264 80060 2292
rect 79508 1692 79560 1698
rect 79508 1634 79560 1640
rect 79888 800 79916 2264
rect 80060 2246 80112 2252
rect 80532 800 80560 2382
rect 81176 800 81204 2518
rect 81440 2304 81492 2310
rect 81440 2246 81492 2252
rect 81452 2038 81480 2246
rect 81440 2032 81492 2038
rect 81440 1974 81492 1980
rect 81820 800 81848 2790
rect 83844 2446 83872 4762
rect 85132 2990 85160 26318
rect 85408 26234 85436 26386
rect 85224 26206 85436 26234
rect 85028 2984 85080 2990
rect 85028 2926 85080 2932
rect 85120 2984 85172 2990
rect 85120 2926 85172 2932
rect 85040 2802 85068 2926
rect 85224 2802 85252 26206
rect 86144 26042 86172 27474
rect 86328 27130 86356 29271
rect 86958 29200 87014 30000
rect 87602 29200 87658 30000
rect 88246 29200 88302 30000
rect 88890 29200 88946 30000
rect 89534 29200 89590 30000
rect 86408 27464 86460 27470
rect 86408 27406 86460 27412
rect 86316 27124 86368 27130
rect 86316 27066 86368 27072
rect 86132 26036 86184 26042
rect 86132 25978 86184 25984
rect 86420 8906 86448 27406
rect 86972 27130 87000 29200
rect 87510 27976 87566 27985
rect 87510 27911 87566 27920
rect 86960 27124 87012 27130
rect 86960 27066 87012 27072
rect 87236 26988 87288 26994
rect 87236 26930 87288 26936
rect 86592 26852 86644 26858
rect 86592 26794 86644 26800
rect 86500 23656 86552 23662
rect 86500 23598 86552 23604
rect 86512 22438 86540 23598
rect 86500 22432 86552 22438
rect 86500 22374 86552 22380
rect 86604 16046 86632 26794
rect 87052 26376 87104 26382
rect 87052 26318 87104 26324
rect 86776 26036 86828 26042
rect 86776 25978 86828 25984
rect 86788 25906 86816 25978
rect 86776 25900 86828 25906
rect 86776 25842 86828 25848
rect 86776 24200 86828 24206
rect 86776 24142 86828 24148
rect 86788 23866 86816 24142
rect 86776 23860 86828 23866
rect 86776 23802 86828 23808
rect 87064 17066 87092 26318
rect 87144 25696 87196 25702
rect 87144 25638 87196 25644
rect 87052 17060 87104 17066
rect 87052 17002 87104 17008
rect 86592 16040 86644 16046
rect 86592 15982 86644 15988
rect 86776 13320 86828 13326
rect 86776 13262 86828 13268
rect 86788 12986 86816 13262
rect 86776 12980 86828 12986
rect 86776 12922 86828 12928
rect 86960 12844 87012 12850
rect 86960 12786 87012 12792
rect 87052 12844 87104 12850
rect 87052 12786 87104 12792
rect 86972 12753 87000 12786
rect 86958 12744 87014 12753
rect 86958 12679 87014 12688
rect 86592 10260 86644 10266
rect 86592 10202 86644 10208
rect 86408 8900 86460 8906
rect 86408 8842 86460 8848
rect 86604 3534 86632 10202
rect 86972 6914 87000 12679
rect 87064 10742 87092 12786
rect 87156 12374 87184 25638
rect 87248 14550 87276 26930
rect 87420 26920 87472 26926
rect 87420 26862 87472 26868
rect 87432 26625 87460 26862
rect 87418 26616 87474 26625
rect 87418 26551 87474 26560
rect 87524 26042 87552 27911
rect 87616 27538 87644 29200
rect 87694 28656 87750 28665
rect 87694 28591 87750 28600
rect 87604 27532 87656 27538
rect 87604 27474 87656 27480
rect 87708 26042 87736 28591
rect 87788 27464 87840 27470
rect 87788 27406 87840 27412
rect 87512 26036 87564 26042
rect 87512 25978 87564 25984
rect 87696 26036 87748 26042
rect 87696 25978 87748 25984
rect 87800 25514 87828 27406
rect 87880 27328 87932 27334
rect 87880 27270 87932 27276
rect 87970 27296 88026 27305
rect 87340 25486 87828 25514
rect 87340 16794 87368 25486
rect 87892 25378 87920 27270
rect 87970 27231 88026 27240
rect 87984 26382 88012 27231
rect 88260 26586 88288 29200
rect 88248 26580 88300 26586
rect 88248 26522 88300 26528
rect 87972 26376 88024 26382
rect 87972 26318 88024 26324
rect 88904 26314 88932 29200
rect 89548 27606 89576 29200
rect 89536 27600 89588 27606
rect 89536 27542 89588 27548
rect 88892 26308 88944 26314
rect 88892 26250 88944 26256
rect 88156 26240 88208 26246
rect 88156 26182 88208 26188
rect 88168 25974 88196 26182
rect 88156 25968 88208 25974
rect 88156 25910 88208 25916
rect 87800 25350 87920 25378
rect 87604 21888 87656 21894
rect 87604 21830 87656 21836
rect 87512 21344 87564 21350
rect 87512 21286 87564 21292
rect 87420 20936 87472 20942
rect 87420 20878 87472 20884
rect 87432 20505 87460 20878
rect 87418 20496 87474 20505
rect 87418 20431 87474 20440
rect 87328 16788 87380 16794
rect 87328 16730 87380 16736
rect 87236 14544 87288 14550
rect 87236 14486 87288 14492
rect 87144 12368 87196 12374
rect 87144 12310 87196 12316
rect 87524 11218 87552 21286
rect 87616 17270 87644 21830
rect 87696 19712 87748 19718
rect 87696 19654 87748 19660
rect 87708 19514 87736 19654
rect 87696 19508 87748 19514
rect 87696 19450 87748 19456
rect 87604 17264 87656 17270
rect 87604 17206 87656 17212
rect 87800 12889 87828 25350
rect 87878 25256 87934 25265
rect 87878 25191 87880 25200
rect 87932 25191 87934 25200
rect 87880 25162 87932 25168
rect 87972 25152 88024 25158
rect 87972 25094 88024 25100
rect 87880 16584 87932 16590
rect 87880 16526 87932 16532
rect 87786 12880 87842 12889
rect 87786 12815 87842 12824
rect 87512 11212 87564 11218
rect 87512 11154 87564 11160
rect 87420 11144 87472 11150
rect 87420 11086 87472 11092
rect 87432 10985 87460 11086
rect 87696 11008 87748 11014
rect 87418 10976 87474 10985
rect 87696 10950 87748 10956
rect 87418 10911 87474 10920
rect 87708 10810 87736 10950
rect 87696 10804 87748 10810
rect 87696 10746 87748 10752
rect 87052 10736 87104 10742
rect 87052 10678 87104 10684
rect 87420 8968 87472 8974
rect 87418 8936 87420 8945
rect 87472 8936 87474 8945
rect 87418 8871 87474 8880
rect 86972 6886 87092 6914
rect 86868 4140 86920 4146
rect 86868 4082 86920 4088
rect 86880 3942 86908 4082
rect 86868 3936 86920 3942
rect 86868 3878 86920 3884
rect 86684 3664 86736 3670
rect 86684 3606 86736 3612
rect 86592 3528 86644 3534
rect 86592 3470 86644 3476
rect 85488 2916 85540 2922
rect 85488 2858 85540 2864
rect 85040 2774 85252 2802
rect 85500 2514 85528 2858
rect 86316 2576 86368 2582
rect 86316 2518 86368 2524
rect 85488 2508 85540 2514
rect 85488 2450 85540 2456
rect 83832 2440 83884 2446
rect 83832 2382 83884 2388
rect 85028 2440 85080 2446
rect 85028 2382 85080 2388
rect 82452 2372 82504 2378
rect 82452 2314 82504 2320
rect 82464 800 82492 2314
rect 82728 2304 82780 2310
rect 82728 2246 82780 2252
rect 83096 2304 83148 2310
rect 83096 2246 83148 2252
rect 84200 2304 84252 2310
rect 84200 2246 84252 2252
rect 84384 2304 84436 2310
rect 84384 2246 84436 2252
rect 82740 2106 82768 2246
rect 82728 2100 82780 2106
rect 82728 2042 82780 2048
rect 83108 800 83136 2246
rect 84212 1834 84240 2246
rect 84200 1828 84252 1834
rect 84200 1770 84252 1776
rect 84396 800 84424 2246
rect 85040 800 85068 2382
rect 85304 2304 85356 2310
rect 85304 2246 85356 2252
rect 85672 2304 85724 2310
rect 85672 2246 85724 2252
rect 85316 1630 85344 2246
rect 85304 1624 85356 1630
rect 85304 1566 85356 1572
rect 85684 800 85712 2246
rect 86328 800 86356 2518
rect 47780 734 47992 762
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 84382 0 84438 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86696 105 86724 3606
rect 86868 2984 86920 2990
rect 86868 2926 86920 2932
rect 86880 921 86908 2926
rect 86960 2848 87012 2854
rect 86960 2790 87012 2796
rect 86866 912 86922 921
rect 86866 847 86922 856
rect 86972 800 87000 2790
rect 87064 2310 87092 6886
rect 87420 6248 87472 6254
rect 87418 6216 87420 6225
rect 87696 6248 87748 6254
rect 87472 6216 87474 6225
rect 87696 6190 87748 6196
rect 87418 6151 87474 6160
rect 87708 5642 87736 6190
rect 87696 5636 87748 5642
rect 87696 5578 87748 5584
rect 87892 4146 87920 16526
rect 87984 13977 88012 25094
rect 88248 24812 88300 24818
rect 88248 24754 88300 24760
rect 88064 24608 88116 24614
rect 88062 24576 88064 24585
rect 88116 24576 88118 24585
rect 88062 24511 88118 24520
rect 88064 24064 88116 24070
rect 88064 24006 88116 24012
rect 88076 23905 88104 24006
rect 88062 23896 88118 23905
rect 88062 23831 88118 23840
rect 88064 23520 88116 23526
rect 88064 23462 88116 23468
rect 88076 23225 88104 23462
rect 88062 23216 88118 23225
rect 88062 23151 88118 23160
rect 88064 22636 88116 22642
rect 88064 22578 88116 22584
rect 88076 22545 88104 22578
rect 88062 22536 88118 22545
rect 88062 22471 88118 22480
rect 88156 22432 88208 22438
rect 88156 22374 88208 22380
rect 88064 21888 88116 21894
rect 88062 21856 88064 21865
rect 88116 21856 88118 21865
rect 88062 21791 88118 21800
rect 88064 21344 88116 21350
rect 88064 21286 88116 21292
rect 88076 21185 88104 21286
rect 88062 21176 88118 21185
rect 88062 21111 88118 21120
rect 88168 20058 88196 22374
rect 88260 20262 88288 24754
rect 88248 20256 88300 20262
rect 88248 20198 88300 20204
rect 88156 20052 88208 20058
rect 88156 19994 88208 20000
rect 88062 19816 88118 19825
rect 88062 19751 88118 19760
rect 88076 19718 88104 19751
rect 88064 19712 88116 19718
rect 88064 19654 88116 19660
rect 88064 19168 88116 19174
rect 88062 19136 88064 19145
rect 88116 19136 88118 19145
rect 88062 19071 88118 19080
rect 88248 18760 88300 18766
rect 88248 18702 88300 18708
rect 88064 18624 88116 18630
rect 88064 18566 88116 18572
rect 88076 18222 88104 18566
rect 88260 18465 88288 18702
rect 88246 18456 88302 18465
rect 88246 18391 88302 18400
rect 88064 18216 88116 18222
rect 88064 18158 88116 18164
rect 88062 17096 88118 17105
rect 88062 17031 88064 17040
rect 88116 17031 88118 17040
rect 88064 17002 88116 17008
rect 88064 16448 88116 16454
rect 88062 16416 88064 16425
rect 88116 16416 88118 16425
rect 88062 16351 88118 16360
rect 88064 15904 88116 15910
rect 88064 15846 88116 15852
rect 88076 15745 88104 15846
rect 88062 15736 88118 15745
rect 88062 15671 88118 15680
rect 88064 15428 88116 15434
rect 88064 15370 88116 15376
rect 88076 15065 88104 15370
rect 88156 15360 88208 15366
rect 88156 15302 88208 15308
rect 88062 15056 88118 15065
rect 88168 15026 88196 15302
rect 88248 15088 88300 15094
rect 88248 15030 88300 15036
rect 88062 14991 88118 15000
rect 88156 15020 88208 15026
rect 88156 14962 88208 14968
rect 88062 14376 88118 14385
rect 88062 14311 88064 14320
rect 88116 14311 88118 14320
rect 88064 14282 88116 14288
rect 88156 14272 88208 14278
rect 88156 14214 88208 14220
rect 87970 13968 88026 13977
rect 87970 13903 88026 13912
rect 88064 13728 88116 13734
rect 88062 13696 88064 13705
rect 88116 13696 88118 13705
rect 88062 13631 88118 13640
rect 88064 13184 88116 13190
rect 88064 13126 88116 13132
rect 88076 13025 88104 13126
rect 88062 13016 88118 13025
rect 88062 12951 88118 12960
rect 88168 12918 88196 14214
rect 88156 12912 88208 12918
rect 88156 12854 88208 12860
rect 88064 12640 88116 12646
rect 88064 12582 88116 12588
rect 88076 12345 88104 12582
rect 88062 12336 88118 12345
rect 88062 12271 88118 12280
rect 88260 11762 88288 15030
rect 88248 11756 88300 11762
rect 88248 11698 88300 11704
rect 88062 11656 88118 11665
rect 88062 11591 88064 11600
rect 88116 11591 88118 11600
rect 88064 11562 88116 11568
rect 88064 10464 88116 10470
rect 88064 10406 88116 10412
rect 88076 10305 88104 10406
rect 88062 10296 88118 10305
rect 88062 10231 88118 10240
rect 88248 8492 88300 8498
rect 88248 8434 88300 8440
rect 88260 8265 88288 8434
rect 88246 8256 88302 8265
rect 88246 8191 88302 8200
rect 88064 7744 88116 7750
rect 88064 7686 88116 7692
rect 88076 7585 88104 7686
rect 88062 7576 88118 7585
rect 88062 7511 88118 7520
rect 88064 7404 88116 7410
rect 88064 7346 88116 7352
rect 88076 6905 88104 7346
rect 88062 6896 88118 6905
rect 88062 6831 88118 6840
rect 87972 5704 88024 5710
rect 87972 5646 88024 5652
rect 87984 5545 88012 5646
rect 87970 5536 88026 5545
rect 87970 5471 88026 5480
rect 88064 5024 88116 5030
rect 88064 4966 88116 4972
rect 88076 4865 88104 4966
rect 88062 4856 88118 4865
rect 88062 4791 88118 4800
rect 88064 4480 88116 4486
rect 88064 4422 88116 4428
rect 88076 4185 88104 4422
rect 88062 4176 88118 4185
rect 87696 4140 87748 4146
rect 87696 4082 87748 4088
rect 87880 4140 87932 4146
rect 88062 4111 88118 4120
rect 87880 4082 87932 4088
rect 87604 3664 87656 3670
rect 87604 3606 87656 3612
rect 87052 2304 87104 2310
rect 87052 2246 87104 2252
rect 87616 800 87644 3606
rect 87708 3194 87736 4082
rect 88248 4004 88300 4010
rect 88248 3946 88300 3952
rect 87880 3936 87932 3942
rect 87880 3878 87932 3884
rect 88064 3936 88116 3942
rect 88064 3878 88116 3884
rect 87892 3738 87920 3878
rect 87788 3732 87840 3738
rect 87788 3674 87840 3680
rect 87880 3732 87932 3738
rect 87880 3674 87932 3680
rect 87800 3194 87828 3674
rect 87696 3188 87748 3194
rect 87696 3130 87748 3136
rect 87788 3188 87840 3194
rect 87788 3130 87840 3136
rect 88076 2825 88104 3878
rect 88156 3528 88208 3534
rect 88156 3470 88208 3476
rect 88062 2816 88118 2825
rect 88062 2751 88118 2760
rect 87972 2304 88024 2310
rect 87972 2246 88024 2252
rect 87984 1766 88012 2246
rect 88168 2145 88196 3470
rect 88154 2136 88210 2145
rect 88154 2071 88210 2080
rect 87972 1760 88024 1766
rect 87972 1702 88024 1708
rect 88260 800 88288 3946
rect 89536 3732 89588 3738
rect 89536 3674 89588 3680
rect 88338 3496 88394 3505
rect 88338 3431 88394 3440
rect 88352 3194 88380 3431
rect 88340 3188 88392 3194
rect 88340 3130 88392 3136
rect 88892 2372 88944 2378
rect 88892 2314 88944 2320
rect 88904 800 88932 2314
rect 89548 800 89576 3674
rect 86682 96 86738 105
rect 86682 31 86738 40
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 89534 0 89590 800
<< via2 >>
rect 1766 28600 1822 28656
rect 1490 27920 1546 27976
rect 2778 29144 2834 29200
rect 1674 26560 1730 26616
rect 1398 25880 1454 25936
rect 1398 25236 1400 25256
rect 1400 25236 1452 25256
rect 1452 25236 1454 25256
rect 1398 25200 1454 25236
rect 1398 24520 1454 24576
rect 1766 23160 1822 23216
rect 1582 22516 1584 22536
rect 1584 22516 1636 22536
rect 1636 22516 1638 22536
rect 1582 22480 1638 22516
rect 1398 21836 1400 21856
rect 1400 21836 1452 21856
rect 1452 21836 1454 21856
rect 1398 21800 1454 21836
rect 1398 21120 1454 21176
rect 1398 20440 1454 20496
rect 1398 19796 1400 19816
rect 1400 19796 1452 19816
rect 1452 19796 1454 19816
rect 1398 19760 1454 19796
rect 1398 18400 1454 18456
rect 1398 17720 1454 17776
rect 1398 16396 1400 16416
rect 1400 16396 1452 16416
rect 1452 16396 1454 16416
rect 1398 16360 1454 16396
rect 1398 15000 1454 15056
rect 1582 15000 1638 15056
rect 1582 14356 1584 14376
rect 1584 14356 1636 14376
rect 1636 14356 1638 14376
rect 1582 14320 1638 14356
rect 1398 13676 1400 13696
rect 1400 13676 1452 13696
rect 1452 13676 1454 13696
rect 1398 13640 1454 13676
rect 1582 12960 1638 13016
rect 1398 12280 1454 12336
rect 1766 19080 1822 19136
rect 3054 27240 3110 27296
rect 1766 17040 1822 17096
rect 1398 11620 1454 11656
rect 1398 11600 1400 11620
rect 1400 11600 1452 11620
rect 1452 11600 1454 11620
rect 1398 10956 1400 10976
rect 1400 10956 1452 10976
rect 1452 10956 1454 10976
rect 1398 10920 1454 10956
rect 1582 10668 1638 10704
rect 1582 10648 1584 10668
rect 1584 10648 1636 10668
rect 1636 10648 1638 10668
rect 1398 10240 1454 10296
rect 1398 9560 1454 9616
rect 1582 8916 1584 8936
rect 1584 8916 1636 8936
rect 1636 8916 1638 8936
rect 1582 8880 1638 8916
rect 1398 8200 1454 8256
rect 1398 6840 1454 6896
rect 1398 5516 1400 5536
rect 1400 5516 1452 5536
rect 1452 5516 1454 5536
rect 1398 5480 1454 5516
rect 1582 4120 1638 4176
rect 1398 3440 1454 3496
rect 1766 6160 1822 6216
rect 1490 2760 1546 2816
rect 2686 2372 2742 2408
rect 2686 2352 2688 2372
rect 2688 2352 2740 2372
rect 2740 2352 2742 2372
rect 11930 27770 11986 27772
rect 12010 27770 12066 27772
rect 12090 27770 12146 27772
rect 12170 27770 12226 27772
rect 11930 27718 11976 27770
rect 11976 27718 11986 27770
rect 12010 27718 12040 27770
rect 12040 27718 12052 27770
rect 12052 27718 12066 27770
rect 12090 27718 12104 27770
rect 12104 27718 12116 27770
rect 12116 27718 12146 27770
rect 12170 27718 12180 27770
rect 12180 27718 12226 27770
rect 11930 27716 11986 27718
rect 12010 27716 12066 27718
rect 12090 27716 12146 27718
rect 12170 27716 12226 27718
rect 11930 26682 11986 26684
rect 12010 26682 12066 26684
rect 12090 26682 12146 26684
rect 12170 26682 12226 26684
rect 11930 26630 11976 26682
rect 11976 26630 11986 26682
rect 12010 26630 12040 26682
rect 12040 26630 12052 26682
rect 12052 26630 12066 26682
rect 12090 26630 12104 26682
rect 12104 26630 12116 26682
rect 12116 26630 12146 26682
rect 12170 26630 12180 26682
rect 12180 26630 12226 26682
rect 11930 26628 11986 26630
rect 12010 26628 12066 26630
rect 12090 26628 12146 26630
rect 12170 26628 12226 26630
rect 11930 25594 11986 25596
rect 12010 25594 12066 25596
rect 12090 25594 12146 25596
rect 12170 25594 12226 25596
rect 11930 25542 11976 25594
rect 11976 25542 11986 25594
rect 12010 25542 12040 25594
rect 12040 25542 12052 25594
rect 12052 25542 12066 25594
rect 12090 25542 12104 25594
rect 12104 25542 12116 25594
rect 12116 25542 12146 25594
rect 12170 25542 12180 25594
rect 12180 25542 12226 25594
rect 11930 25540 11986 25542
rect 12010 25540 12066 25542
rect 12090 25540 12146 25542
rect 12170 25540 12226 25542
rect 11930 24506 11986 24508
rect 12010 24506 12066 24508
rect 12090 24506 12146 24508
rect 12170 24506 12226 24508
rect 11930 24454 11976 24506
rect 11976 24454 11986 24506
rect 12010 24454 12040 24506
rect 12040 24454 12052 24506
rect 12052 24454 12066 24506
rect 12090 24454 12104 24506
rect 12104 24454 12116 24506
rect 12116 24454 12146 24506
rect 12170 24454 12180 24506
rect 12180 24454 12226 24506
rect 11930 24452 11986 24454
rect 12010 24452 12066 24454
rect 12090 24452 12146 24454
rect 12170 24452 12226 24454
rect 11930 23418 11986 23420
rect 12010 23418 12066 23420
rect 12090 23418 12146 23420
rect 12170 23418 12226 23420
rect 11930 23366 11976 23418
rect 11976 23366 11986 23418
rect 12010 23366 12040 23418
rect 12040 23366 12052 23418
rect 12052 23366 12066 23418
rect 12090 23366 12104 23418
rect 12104 23366 12116 23418
rect 12116 23366 12146 23418
rect 12170 23366 12180 23418
rect 12180 23366 12226 23418
rect 11930 23364 11986 23366
rect 12010 23364 12066 23366
rect 12090 23364 12146 23366
rect 12170 23364 12226 23366
rect 11930 22330 11986 22332
rect 12010 22330 12066 22332
rect 12090 22330 12146 22332
rect 12170 22330 12226 22332
rect 11930 22278 11976 22330
rect 11976 22278 11986 22330
rect 12010 22278 12040 22330
rect 12040 22278 12052 22330
rect 12052 22278 12066 22330
rect 12090 22278 12104 22330
rect 12104 22278 12116 22330
rect 12116 22278 12146 22330
rect 12170 22278 12180 22330
rect 12180 22278 12226 22330
rect 11930 22276 11986 22278
rect 12010 22276 12066 22278
rect 12090 22276 12146 22278
rect 12170 22276 12226 22278
rect 11930 21242 11986 21244
rect 12010 21242 12066 21244
rect 12090 21242 12146 21244
rect 12170 21242 12226 21244
rect 11930 21190 11976 21242
rect 11976 21190 11986 21242
rect 12010 21190 12040 21242
rect 12040 21190 12052 21242
rect 12052 21190 12066 21242
rect 12090 21190 12104 21242
rect 12104 21190 12116 21242
rect 12116 21190 12146 21242
rect 12170 21190 12180 21242
rect 12180 21190 12226 21242
rect 11930 21188 11986 21190
rect 12010 21188 12066 21190
rect 12090 21188 12146 21190
rect 12170 21188 12226 21190
rect 11930 20154 11986 20156
rect 12010 20154 12066 20156
rect 12090 20154 12146 20156
rect 12170 20154 12226 20156
rect 11930 20102 11976 20154
rect 11976 20102 11986 20154
rect 12010 20102 12040 20154
rect 12040 20102 12052 20154
rect 12052 20102 12066 20154
rect 12090 20102 12104 20154
rect 12104 20102 12116 20154
rect 12116 20102 12146 20154
rect 12170 20102 12180 20154
rect 12180 20102 12226 20154
rect 11930 20100 11986 20102
rect 12010 20100 12066 20102
rect 12090 20100 12146 20102
rect 12170 20100 12226 20102
rect 11930 19066 11986 19068
rect 12010 19066 12066 19068
rect 12090 19066 12146 19068
rect 12170 19066 12226 19068
rect 11930 19014 11976 19066
rect 11976 19014 11986 19066
rect 12010 19014 12040 19066
rect 12040 19014 12052 19066
rect 12052 19014 12066 19066
rect 12090 19014 12104 19066
rect 12104 19014 12116 19066
rect 12116 19014 12146 19066
rect 12170 19014 12180 19066
rect 12180 19014 12226 19066
rect 11930 19012 11986 19014
rect 12010 19012 12066 19014
rect 12090 19012 12146 19014
rect 12170 19012 12226 19014
rect 12254 18264 12310 18320
rect 11930 17978 11986 17980
rect 12010 17978 12066 17980
rect 12090 17978 12146 17980
rect 12170 17978 12226 17980
rect 11930 17926 11976 17978
rect 11976 17926 11986 17978
rect 12010 17926 12040 17978
rect 12040 17926 12052 17978
rect 12052 17926 12066 17978
rect 12090 17926 12104 17978
rect 12104 17926 12116 17978
rect 12116 17926 12146 17978
rect 12170 17926 12180 17978
rect 12180 17926 12226 17978
rect 11930 17924 11986 17926
rect 12010 17924 12066 17926
rect 12090 17924 12146 17926
rect 12170 17924 12226 17926
rect 11930 16890 11986 16892
rect 12010 16890 12066 16892
rect 12090 16890 12146 16892
rect 12170 16890 12226 16892
rect 11930 16838 11976 16890
rect 11976 16838 11986 16890
rect 12010 16838 12040 16890
rect 12040 16838 12052 16890
rect 12052 16838 12066 16890
rect 12090 16838 12104 16890
rect 12104 16838 12116 16890
rect 12116 16838 12146 16890
rect 12170 16838 12180 16890
rect 12180 16838 12226 16890
rect 11930 16836 11986 16838
rect 12010 16836 12066 16838
rect 12090 16836 12146 16838
rect 12170 16836 12226 16838
rect 11930 15802 11986 15804
rect 12010 15802 12066 15804
rect 12090 15802 12146 15804
rect 12170 15802 12226 15804
rect 11930 15750 11976 15802
rect 11976 15750 11986 15802
rect 12010 15750 12040 15802
rect 12040 15750 12052 15802
rect 12052 15750 12066 15802
rect 12090 15750 12104 15802
rect 12104 15750 12116 15802
rect 12116 15750 12146 15802
rect 12170 15750 12180 15802
rect 12180 15750 12226 15802
rect 11930 15748 11986 15750
rect 12010 15748 12066 15750
rect 12090 15748 12146 15750
rect 12170 15748 12226 15750
rect 11930 14714 11986 14716
rect 12010 14714 12066 14716
rect 12090 14714 12146 14716
rect 12170 14714 12226 14716
rect 11930 14662 11976 14714
rect 11976 14662 11986 14714
rect 12010 14662 12040 14714
rect 12040 14662 12052 14714
rect 12052 14662 12066 14714
rect 12090 14662 12104 14714
rect 12104 14662 12116 14714
rect 12116 14662 12146 14714
rect 12170 14662 12180 14714
rect 12180 14662 12226 14714
rect 11930 14660 11986 14662
rect 12010 14660 12066 14662
rect 12090 14660 12146 14662
rect 12170 14660 12226 14662
rect 11930 13626 11986 13628
rect 12010 13626 12066 13628
rect 12090 13626 12146 13628
rect 12170 13626 12226 13628
rect 11930 13574 11976 13626
rect 11976 13574 11986 13626
rect 12010 13574 12040 13626
rect 12040 13574 12052 13626
rect 12052 13574 12066 13626
rect 12090 13574 12104 13626
rect 12104 13574 12116 13626
rect 12116 13574 12146 13626
rect 12170 13574 12180 13626
rect 12180 13574 12226 13626
rect 11930 13572 11986 13574
rect 12010 13572 12066 13574
rect 12090 13572 12146 13574
rect 12170 13572 12226 13574
rect 11930 12538 11986 12540
rect 12010 12538 12066 12540
rect 12090 12538 12146 12540
rect 12170 12538 12226 12540
rect 11930 12486 11976 12538
rect 11976 12486 11986 12538
rect 12010 12486 12040 12538
rect 12040 12486 12052 12538
rect 12052 12486 12066 12538
rect 12090 12486 12104 12538
rect 12104 12486 12116 12538
rect 12116 12486 12146 12538
rect 12170 12486 12180 12538
rect 12180 12486 12226 12538
rect 11930 12484 11986 12486
rect 12010 12484 12066 12486
rect 12090 12484 12146 12486
rect 12170 12484 12226 12486
rect 11930 11450 11986 11452
rect 12010 11450 12066 11452
rect 12090 11450 12146 11452
rect 12170 11450 12226 11452
rect 11930 11398 11976 11450
rect 11976 11398 11986 11450
rect 12010 11398 12040 11450
rect 12040 11398 12052 11450
rect 12052 11398 12066 11450
rect 12090 11398 12104 11450
rect 12104 11398 12116 11450
rect 12116 11398 12146 11450
rect 12170 11398 12180 11450
rect 12180 11398 12226 11450
rect 11930 11396 11986 11398
rect 12010 11396 12066 11398
rect 12090 11396 12146 11398
rect 12170 11396 12226 11398
rect 14462 11348 14518 11384
rect 15106 15408 15162 15464
rect 14462 11328 14464 11348
rect 14464 11328 14516 11348
rect 14516 11328 14518 11348
rect 11930 10362 11986 10364
rect 12010 10362 12066 10364
rect 12090 10362 12146 10364
rect 12170 10362 12226 10364
rect 11930 10310 11976 10362
rect 11976 10310 11986 10362
rect 12010 10310 12040 10362
rect 12040 10310 12052 10362
rect 12052 10310 12066 10362
rect 12090 10310 12104 10362
rect 12104 10310 12116 10362
rect 12116 10310 12146 10362
rect 12170 10310 12180 10362
rect 12180 10310 12226 10362
rect 11930 10308 11986 10310
rect 12010 10308 12066 10310
rect 12090 10308 12146 10310
rect 12170 10308 12226 10310
rect 11930 9274 11986 9276
rect 12010 9274 12066 9276
rect 12090 9274 12146 9276
rect 12170 9274 12226 9276
rect 11930 9222 11976 9274
rect 11976 9222 11986 9274
rect 12010 9222 12040 9274
rect 12040 9222 12052 9274
rect 12052 9222 12066 9274
rect 12090 9222 12104 9274
rect 12104 9222 12116 9274
rect 12116 9222 12146 9274
rect 12170 9222 12180 9274
rect 12180 9222 12226 9274
rect 11930 9220 11986 9222
rect 12010 9220 12066 9222
rect 12090 9220 12146 9222
rect 12170 9220 12226 9222
rect 11930 8186 11986 8188
rect 12010 8186 12066 8188
rect 12090 8186 12146 8188
rect 12170 8186 12226 8188
rect 11930 8134 11976 8186
rect 11976 8134 11986 8186
rect 12010 8134 12040 8186
rect 12040 8134 12052 8186
rect 12052 8134 12066 8186
rect 12090 8134 12104 8186
rect 12104 8134 12116 8186
rect 12116 8134 12146 8186
rect 12170 8134 12180 8186
rect 12180 8134 12226 8186
rect 11930 8132 11986 8134
rect 12010 8132 12066 8134
rect 12090 8132 12146 8134
rect 12170 8132 12226 8134
rect 11930 7098 11986 7100
rect 12010 7098 12066 7100
rect 12090 7098 12146 7100
rect 12170 7098 12226 7100
rect 11930 7046 11976 7098
rect 11976 7046 11986 7098
rect 12010 7046 12040 7098
rect 12040 7046 12052 7098
rect 12052 7046 12066 7098
rect 12090 7046 12104 7098
rect 12104 7046 12116 7098
rect 12116 7046 12146 7098
rect 12170 7046 12180 7098
rect 12180 7046 12226 7098
rect 11930 7044 11986 7046
rect 12010 7044 12066 7046
rect 12090 7044 12146 7046
rect 12170 7044 12226 7046
rect 11930 6010 11986 6012
rect 12010 6010 12066 6012
rect 12090 6010 12146 6012
rect 12170 6010 12226 6012
rect 11930 5958 11976 6010
rect 11976 5958 11986 6010
rect 12010 5958 12040 6010
rect 12040 5958 12052 6010
rect 12052 5958 12066 6010
rect 12090 5958 12104 6010
rect 12104 5958 12116 6010
rect 12116 5958 12146 6010
rect 12170 5958 12180 6010
rect 12180 5958 12226 6010
rect 11930 5956 11986 5958
rect 12010 5956 12066 5958
rect 12090 5956 12146 5958
rect 12170 5956 12226 5958
rect 11930 4922 11986 4924
rect 12010 4922 12066 4924
rect 12090 4922 12146 4924
rect 12170 4922 12226 4924
rect 11930 4870 11976 4922
rect 11976 4870 11986 4922
rect 12010 4870 12040 4922
rect 12040 4870 12052 4922
rect 12052 4870 12066 4922
rect 12090 4870 12104 4922
rect 12104 4870 12116 4922
rect 12116 4870 12146 4922
rect 12170 4870 12180 4922
rect 12180 4870 12226 4922
rect 11930 4868 11986 4870
rect 12010 4868 12066 4870
rect 12090 4868 12146 4870
rect 12170 4868 12226 4870
rect 11930 3834 11986 3836
rect 12010 3834 12066 3836
rect 12090 3834 12146 3836
rect 12170 3834 12226 3836
rect 11930 3782 11976 3834
rect 11976 3782 11986 3834
rect 12010 3782 12040 3834
rect 12040 3782 12052 3834
rect 12052 3782 12066 3834
rect 12090 3782 12104 3834
rect 12104 3782 12116 3834
rect 12116 3782 12146 3834
rect 12170 3782 12180 3834
rect 12180 3782 12226 3834
rect 11930 3780 11986 3782
rect 12010 3780 12066 3782
rect 12090 3780 12146 3782
rect 12170 3780 12226 3782
rect 2962 2080 3018 2136
rect 2778 1400 2834 1456
rect 4066 856 4122 912
rect 11930 2746 11986 2748
rect 12010 2746 12066 2748
rect 12090 2746 12146 2748
rect 12170 2746 12226 2748
rect 11930 2694 11976 2746
rect 11976 2694 11986 2746
rect 12010 2694 12040 2746
rect 12040 2694 12052 2746
rect 12052 2694 12066 2746
rect 12090 2694 12104 2746
rect 12104 2694 12116 2746
rect 12116 2694 12146 2746
rect 12170 2694 12180 2746
rect 12180 2694 12226 2746
rect 11930 2692 11986 2694
rect 12010 2692 12066 2694
rect 12090 2692 12146 2694
rect 12170 2692 12226 2694
rect 18878 11328 18934 11384
rect 19890 13640 19946 13696
rect 20074 13504 20130 13560
rect 19982 12552 20038 12608
rect 21822 16904 21878 16960
rect 21178 13232 21234 13288
rect 21086 11600 21142 11656
rect 22006 14864 22062 14920
rect 21914 14320 21970 14376
rect 22098 13912 22154 13968
rect 22374 17584 22430 17640
rect 22904 27226 22960 27228
rect 22984 27226 23040 27228
rect 23064 27226 23120 27228
rect 23144 27226 23200 27228
rect 22904 27174 22950 27226
rect 22950 27174 22960 27226
rect 22984 27174 23014 27226
rect 23014 27174 23026 27226
rect 23026 27174 23040 27226
rect 23064 27174 23078 27226
rect 23078 27174 23090 27226
rect 23090 27174 23120 27226
rect 23144 27174 23154 27226
rect 23154 27174 23200 27226
rect 22904 27172 22960 27174
rect 22984 27172 23040 27174
rect 23064 27172 23120 27174
rect 23144 27172 23200 27174
rect 23386 26696 23442 26752
rect 22904 26138 22960 26140
rect 22984 26138 23040 26140
rect 23064 26138 23120 26140
rect 23144 26138 23200 26140
rect 22904 26086 22950 26138
rect 22950 26086 22960 26138
rect 22984 26086 23014 26138
rect 23014 26086 23026 26138
rect 23026 26086 23040 26138
rect 23064 26086 23078 26138
rect 23078 26086 23090 26138
rect 23090 26086 23120 26138
rect 23144 26086 23154 26138
rect 23154 26086 23200 26138
rect 22904 26084 22960 26086
rect 22984 26084 23040 26086
rect 23064 26084 23120 26086
rect 23144 26084 23200 26086
rect 22904 25050 22960 25052
rect 22984 25050 23040 25052
rect 23064 25050 23120 25052
rect 23144 25050 23200 25052
rect 22904 24998 22950 25050
rect 22950 24998 22960 25050
rect 22984 24998 23014 25050
rect 23014 24998 23026 25050
rect 23026 24998 23040 25050
rect 23064 24998 23078 25050
rect 23078 24998 23090 25050
rect 23090 24998 23120 25050
rect 23144 24998 23154 25050
rect 23154 24998 23200 25050
rect 22904 24996 22960 24998
rect 22984 24996 23040 24998
rect 23064 24996 23120 24998
rect 23144 24996 23200 24998
rect 22904 23962 22960 23964
rect 22984 23962 23040 23964
rect 23064 23962 23120 23964
rect 23144 23962 23200 23964
rect 22904 23910 22950 23962
rect 22950 23910 22960 23962
rect 22984 23910 23014 23962
rect 23014 23910 23026 23962
rect 23026 23910 23040 23962
rect 23064 23910 23078 23962
rect 23078 23910 23090 23962
rect 23090 23910 23120 23962
rect 23144 23910 23154 23962
rect 23154 23910 23200 23962
rect 22904 23908 22960 23910
rect 22984 23908 23040 23910
rect 23064 23908 23120 23910
rect 23144 23908 23200 23910
rect 22904 22874 22960 22876
rect 22984 22874 23040 22876
rect 23064 22874 23120 22876
rect 23144 22874 23200 22876
rect 22904 22822 22950 22874
rect 22950 22822 22960 22874
rect 22984 22822 23014 22874
rect 23014 22822 23026 22874
rect 23026 22822 23040 22874
rect 23064 22822 23078 22874
rect 23078 22822 23090 22874
rect 23090 22822 23120 22874
rect 23144 22822 23154 22874
rect 23154 22822 23200 22874
rect 22904 22820 22960 22822
rect 22984 22820 23040 22822
rect 23064 22820 23120 22822
rect 23144 22820 23200 22822
rect 22904 21786 22960 21788
rect 22984 21786 23040 21788
rect 23064 21786 23120 21788
rect 23144 21786 23200 21788
rect 22904 21734 22950 21786
rect 22950 21734 22960 21786
rect 22984 21734 23014 21786
rect 23014 21734 23026 21786
rect 23026 21734 23040 21786
rect 23064 21734 23078 21786
rect 23078 21734 23090 21786
rect 23090 21734 23120 21786
rect 23144 21734 23154 21786
rect 23154 21734 23200 21786
rect 22904 21732 22960 21734
rect 22984 21732 23040 21734
rect 23064 21732 23120 21734
rect 23144 21732 23200 21734
rect 22904 20698 22960 20700
rect 22984 20698 23040 20700
rect 23064 20698 23120 20700
rect 23144 20698 23200 20700
rect 22904 20646 22950 20698
rect 22950 20646 22960 20698
rect 22984 20646 23014 20698
rect 23014 20646 23026 20698
rect 23026 20646 23040 20698
rect 23064 20646 23078 20698
rect 23078 20646 23090 20698
rect 23090 20646 23120 20698
rect 23144 20646 23154 20698
rect 23154 20646 23200 20698
rect 22904 20644 22960 20646
rect 22984 20644 23040 20646
rect 23064 20644 23120 20646
rect 23144 20644 23200 20646
rect 22904 19610 22960 19612
rect 22984 19610 23040 19612
rect 23064 19610 23120 19612
rect 23144 19610 23200 19612
rect 22904 19558 22950 19610
rect 22950 19558 22960 19610
rect 22984 19558 23014 19610
rect 23014 19558 23026 19610
rect 23026 19558 23040 19610
rect 23064 19558 23078 19610
rect 23078 19558 23090 19610
rect 23090 19558 23120 19610
rect 23144 19558 23154 19610
rect 23154 19558 23200 19610
rect 22904 19556 22960 19558
rect 22984 19556 23040 19558
rect 23064 19556 23120 19558
rect 23144 19556 23200 19558
rect 22904 18522 22960 18524
rect 22984 18522 23040 18524
rect 23064 18522 23120 18524
rect 23144 18522 23200 18524
rect 22904 18470 22950 18522
rect 22950 18470 22960 18522
rect 22984 18470 23014 18522
rect 23014 18470 23026 18522
rect 23026 18470 23040 18522
rect 23064 18470 23078 18522
rect 23078 18470 23090 18522
rect 23090 18470 23120 18522
rect 23144 18470 23154 18522
rect 23154 18470 23200 18522
rect 22904 18468 22960 18470
rect 22984 18468 23040 18470
rect 23064 18468 23120 18470
rect 23144 18468 23200 18470
rect 22904 17434 22960 17436
rect 22984 17434 23040 17436
rect 23064 17434 23120 17436
rect 23144 17434 23200 17436
rect 22904 17382 22950 17434
rect 22950 17382 22960 17434
rect 22984 17382 23014 17434
rect 23014 17382 23026 17434
rect 23026 17382 23040 17434
rect 23064 17382 23078 17434
rect 23078 17382 23090 17434
rect 23090 17382 23120 17434
rect 23144 17382 23154 17434
rect 23154 17382 23200 17434
rect 22904 17380 22960 17382
rect 22984 17380 23040 17382
rect 23064 17380 23120 17382
rect 23144 17380 23200 17382
rect 22904 16346 22960 16348
rect 22984 16346 23040 16348
rect 23064 16346 23120 16348
rect 23144 16346 23200 16348
rect 22904 16294 22950 16346
rect 22950 16294 22960 16346
rect 22984 16294 23014 16346
rect 23014 16294 23026 16346
rect 23026 16294 23040 16346
rect 23064 16294 23078 16346
rect 23078 16294 23090 16346
rect 23090 16294 23120 16346
rect 23144 16294 23154 16346
rect 23154 16294 23200 16346
rect 22904 16292 22960 16294
rect 22984 16292 23040 16294
rect 23064 16292 23120 16294
rect 23144 16292 23200 16294
rect 22098 13796 22154 13832
rect 22098 13776 22100 13796
rect 22100 13776 22152 13796
rect 22152 13776 22154 13796
rect 21546 11328 21602 11384
rect 22904 15258 22960 15260
rect 22984 15258 23040 15260
rect 23064 15258 23120 15260
rect 23144 15258 23200 15260
rect 22904 15206 22950 15258
rect 22950 15206 22960 15258
rect 22984 15206 23014 15258
rect 23014 15206 23026 15258
rect 23026 15206 23040 15258
rect 23064 15206 23078 15258
rect 23078 15206 23090 15258
rect 23090 15206 23120 15258
rect 23144 15206 23154 15258
rect 23154 15206 23200 15258
rect 22904 15204 22960 15206
rect 22984 15204 23040 15206
rect 23064 15204 23120 15206
rect 23144 15204 23200 15206
rect 25410 27396 25466 27432
rect 25410 27376 25412 27396
rect 25412 27376 25464 27396
rect 25464 27376 25466 27396
rect 23386 15272 23442 15328
rect 23110 14764 23112 14784
rect 23112 14764 23164 14784
rect 23164 14764 23166 14784
rect 23110 14728 23166 14764
rect 22834 14456 22890 14512
rect 23294 14320 23350 14376
rect 22904 14170 22960 14172
rect 22984 14170 23040 14172
rect 23064 14170 23120 14172
rect 23144 14170 23200 14172
rect 22904 14118 22950 14170
rect 22950 14118 22960 14170
rect 22984 14118 23014 14170
rect 23014 14118 23026 14170
rect 23026 14118 23040 14170
rect 23064 14118 23078 14170
rect 23078 14118 23090 14170
rect 23090 14118 23120 14170
rect 23144 14118 23154 14170
rect 23154 14118 23200 14170
rect 22904 14116 22960 14118
rect 22984 14116 23040 14118
rect 23064 14116 23120 14118
rect 23144 14116 23200 14118
rect 22834 13932 22890 13968
rect 22834 13912 22836 13932
rect 22836 13912 22888 13932
rect 22888 13912 22890 13932
rect 22904 13082 22960 13084
rect 22984 13082 23040 13084
rect 23064 13082 23120 13084
rect 23144 13082 23200 13084
rect 22904 13030 22950 13082
rect 22950 13030 22960 13082
rect 22984 13030 23014 13082
rect 23014 13030 23026 13082
rect 23026 13030 23040 13082
rect 23064 13030 23078 13082
rect 23078 13030 23090 13082
rect 23090 13030 23120 13082
rect 23144 13030 23154 13082
rect 23154 13030 23200 13082
rect 22904 13028 22960 13030
rect 22984 13028 23040 13030
rect 23064 13028 23120 13030
rect 23144 13028 23200 13030
rect 23938 14184 23994 14240
rect 24214 15680 24270 15736
rect 24122 14592 24178 14648
rect 22904 11994 22960 11996
rect 22984 11994 23040 11996
rect 23064 11994 23120 11996
rect 23144 11994 23200 11996
rect 22904 11942 22950 11994
rect 22950 11942 22960 11994
rect 22984 11942 23014 11994
rect 23014 11942 23026 11994
rect 23026 11942 23040 11994
rect 23064 11942 23078 11994
rect 23078 11942 23090 11994
rect 23090 11942 23120 11994
rect 23144 11942 23154 11994
rect 23154 11942 23200 11994
rect 22904 11940 22960 11942
rect 22984 11940 23040 11942
rect 23064 11940 23120 11942
rect 23144 11940 23200 11942
rect 22904 10906 22960 10908
rect 22984 10906 23040 10908
rect 23064 10906 23120 10908
rect 23144 10906 23200 10908
rect 22904 10854 22950 10906
rect 22950 10854 22960 10906
rect 22984 10854 23014 10906
rect 23014 10854 23026 10906
rect 23026 10854 23040 10906
rect 23064 10854 23078 10906
rect 23078 10854 23090 10906
rect 23090 10854 23120 10906
rect 23144 10854 23154 10906
rect 23154 10854 23200 10906
rect 22904 10852 22960 10854
rect 22984 10852 23040 10854
rect 23064 10852 23120 10854
rect 23144 10852 23200 10854
rect 22904 9818 22960 9820
rect 22984 9818 23040 9820
rect 23064 9818 23120 9820
rect 23144 9818 23200 9820
rect 22904 9766 22950 9818
rect 22950 9766 22960 9818
rect 22984 9766 23014 9818
rect 23014 9766 23026 9818
rect 23026 9766 23040 9818
rect 23064 9766 23078 9818
rect 23078 9766 23090 9818
rect 23090 9766 23120 9818
rect 23144 9766 23154 9818
rect 23154 9766 23200 9818
rect 22904 9764 22960 9766
rect 22984 9764 23040 9766
rect 23064 9764 23120 9766
rect 23144 9764 23200 9766
rect 22904 8730 22960 8732
rect 22984 8730 23040 8732
rect 23064 8730 23120 8732
rect 23144 8730 23200 8732
rect 22904 8678 22950 8730
rect 22950 8678 22960 8730
rect 22984 8678 23014 8730
rect 23014 8678 23026 8730
rect 23026 8678 23040 8730
rect 23064 8678 23078 8730
rect 23078 8678 23090 8730
rect 23090 8678 23120 8730
rect 23144 8678 23154 8730
rect 23154 8678 23200 8730
rect 22904 8676 22960 8678
rect 22984 8676 23040 8678
rect 23064 8676 23120 8678
rect 23144 8676 23200 8678
rect 22904 7642 22960 7644
rect 22984 7642 23040 7644
rect 23064 7642 23120 7644
rect 23144 7642 23200 7644
rect 22904 7590 22950 7642
rect 22950 7590 22960 7642
rect 22984 7590 23014 7642
rect 23014 7590 23026 7642
rect 23026 7590 23040 7642
rect 23064 7590 23078 7642
rect 23078 7590 23090 7642
rect 23090 7590 23120 7642
rect 23144 7590 23154 7642
rect 23154 7590 23200 7642
rect 22904 7588 22960 7590
rect 22984 7588 23040 7590
rect 23064 7588 23120 7590
rect 23144 7588 23200 7590
rect 22904 6554 22960 6556
rect 22984 6554 23040 6556
rect 23064 6554 23120 6556
rect 23144 6554 23200 6556
rect 22904 6502 22950 6554
rect 22950 6502 22960 6554
rect 22984 6502 23014 6554
rect 23014 6502 23026 6554
rect 23026 6502 23040 6554
rect 23064 6502 23078 6554
rect 23078 6502 23090 6554
rect 23090 6502 23120 6554
rect 23144 6502 23154 6554
rect 23154 6502 23200 6554
rect 22904 6500 22960 6502
rect 22984 6500 23040 6502
rect 23064 6500 23120 6502
rect 23144 6500 23200 6502
rect 22904 5466 22960 5468
rect 22984 5466 23040 5468
rect 23064 5466 23120 5468
rect 23144 5466 23200 5468
rect 22904 5414 22950 5466
rect 22950 5414 22960 5466
rect 22984 5414 23014 5466
rect 23014 5414 23026 5466
rect 23026 5414 23040 5466
rect 23064 5414 23078 5466
rect 23078 5414 23090 5466
rect 23090 5414 23120 5466
rect 23144 5414 23154 5466
rect 23154 5414 23200 5466
rect 22904 5412 22960 5414
rect 22984 5412 23040 5414
rect 23064 5412 23120 5414
rect 23144 5412 23200 5414
rect 22904 4378 22960 4380
rect 22984 4378 23040 4380
rect 23064 4378 23120 4380
rect 23144 4378 23200 4380
rect 22904 4326 22950 4378
rect 22950 4326 22960 4378
rect 22984 4326 23014 4378
rect 23014 4326 23026 4378
rect 23026 4326 23040 4378
rect 23064 4326 23078 4378
rect 23078 4326 23090 4378
rect 23090 4326 23120 4378
rect 23144 4326 23154 4378
rect 23154 4326 23200 4378
rect 22904 4324 22960 4326
rect 22984 4324 23040 4326
rect 23064 4324 23120 4326
rect 23144 4324 23200 4326
rect 22904 3290 22960 3292
rect 22984 3290 23040 3292
rect 23064 3290 23120 3292
rect 23144 3290 23200 3292
rect 22904 3238 22950 3290
rect 22950 3238 22960 3290
rect 22984 3238 23014 3290
rect 23014 3238 23026 3290
rect 23026 3238 23040 3290
rect 23064 3238 23078 3290
rect 23078 3238 23090 3290
rect 23090 3238 23120 3290
rect 23144 3238 23154 3290
rect 23154 3238 23200 3290
rect 22904 3236 22960 3238
rect 22984 3236 23040 3238
rect 23064 3236 23120 3238
rect 23144 3236 23200 3238
rect 22904 2202 22960 2204
rect 22984 2202 23040 2204
rect 23064 2202 23120 2204
rect 23144 2202 23200 2204
rect 22904 2150 22950 2202
rect 22950 2150 22960 2202
rect 22984 2150 23014 2202
rect 23014 2150 23026 2202
rect 23026 2150 23040 2202
rect 23064 2150 23078 2202
rect 23078 2150 23090 2202
rect 23090 2150 23120 2202
rect 23144 2150 23154 2202
rect 23154 2150 23200 2202
rect 22904 2148 22960 2150
rect 22984 2148 23040 2150
rect 23064 2148 23120 2150
rect 23144 2148 23200 2150
rect 23938 13096 23994 13152
rect 24582 17484 24584 17504
rect 24584 17484 24636 17504
rect 24636 17484 24638 17504
rect 24582 17448 24638 17484
rect 24674 17076 24676 17096
rect 24676 17076 24728 17096
rect 24728 17076 24730 17096
rect 24674 17040 24730 17076
rect 25042 16224 25098 16280
rect 24030 12824 24086 12880
rect 24214 12960 24270 13016
rect 25410 15816 25466 15872
rect 25870 16768 25926 16824
rect 25778 16224 25834 16280
rect 26422 26560 26478 26616
rect 26330 17484 26332 17504
rect 26332 17484 26384 17504
rect 26384 17484 26386 17504
rect 26330 17448 26386 17484
rect 26146 16224 26202 16280
rect 26054 16088 26110 16144
rect 25594 14456 25650 14512
rect 25870 14320 25926 14376
rect 25042 13368 25098 13424
rect 27342 26560 27398 26616
rect 26146 14320 26202 14376
rect 27526 26424 27582 26480
rect 27802 26696 27858 26752
rect 26974 16224 27030 16280
rect 24674 12416 24730 12472
rect 24306 11192 24362 11248
rect 24306 11076 24362 11112
rect 24306 11056 24308 11076
rect 24308 11056 24360 11076
rect 24360 11056 24362 11076
rect 25134 12280 25190 12336
rect 25226 12180 25228 12200
rect 25228 12180 25280 12200
rect 25280 12180 25282 12200
rect 25226 12144 25282 12180
rect 25318 12008 25374 12064
rect 25042 11872 25098 11928
rect 25686 11736 25742 11792
rect 26054 13232 26110 13288
rect 26146 12960 26202 13016
rect 26330 13096 26386 13152
rect 26698 14356 26700 14376
rect 26700 14356 26752 14376
rect 26752 14356 26754 14376
rect 26698 14320 26754 14356
rect 26514 12844 26570 12880
rect 26514 12824 26516 12844
rect 26516 12824 26568 12844
rect 26568 12824 26570 12844
rect 26790 13640 26846 13696
rect 26054 12688 26110 12744
rect 26330 12552 26386 12608
rect 26882 13504 26938 13560
rect 25594 11500 25596 11520
rect 25596 11500 25648 11520
rect 25648 11500 25650 11520
rect 25594 11464 25650 11500
rect 25870 11328 25926 11384
rect 26054 11600 26110 11656
rect 24214 2216 24270 2272
rect 26422 12008 26478 12064
rect 26514 11872 26570 11928
rect 26330 11464 26386 11520
rect 26238 11192 26294 11248
rect 25962 3052 26018 3088
rect 25962 3032 25964 3052
rect 25964 3032 26016 3052
rect 26016 3032 26018 3052
rect 27158 17720 27214 17776
rect 27342 15952 27398 16008
rect 27434 15680 27490 15736
rect 27342 15156 27398 15192
rect 27710 15952 27766 16008
rect 27342 15136 27344 15156
rect 27344 15136 27396 15156
rect 27396 15136 27398 15156
rect 27066 14456 27122 14512
rect 26974 12552 27030 12608
rect 27802 15816 27858 15872
rect 27894 15564 27950 15600
rect 27894 15544 27896 15564
rect 27896 15544 27948 15564
rect 27948 15544 27950 15564
rect 28078 16768 28134 16824
rect 28446 17584 28502 17640
rect 28354 17076 28356 17096
rect 28356 17076 28408 17096
rect 28408 17076 28410 17096
rect 28354 17040 28410 17076
rect 28262 16904 28318 16960
rect 28538 16940 28540 16960
rect 28540 16940 28592 16960
rect 28592 16940 28594 16960
rect 28538 16904 28594 16940
rect 27802 13912 27858 13968
rect 27894 13404 27896 13424
rect 27896 13404 27948 13424
rect 27948 13404 27950 13424
rect 27894 13368 27950 13404
rect 28262 16224 28318 16280
rect 28170 14592 28226 14648
rect 28078 13948 28080 13968
rect 28080 13948 28132 13968
rect 28132 13948 28134 13968
rect 28078 13912 28134 13948
rect 26330 2488 26386 2544
rect 26330 1828 26386 1864
rect 26330 1808 26332 1828
rect 26332 1808 26384 1828
rect 26384 1808 26386 1828
rect 27986 12280 28042 12336
rect 28538 14864 28594 14920
rect 28538 14764 28540 14784
rect 28540 14764 28592 14784
rect 28592 14764 28594 14784
rect 28538 14728 28594 14764
rect 29366 26832 29422 26888
rect 29642 26560 29698 26616
rect 28998 17720 29054 17776
rect 29182 15988 29184 16008
rect 29184 15988 29236 16008
rect 29236 15988 29238 16008
rect 29182 15952 29238 15988
rect 28906 15272 28962 15328
rect 28814 14184 28870 14240
rect 28354 12416 28410 12472
rect 28262 12316 28264 12336
rect 28264 12316 28316 12336
rect 28316 12316 28318 12336
rect 28262 12280 28318 12316
rect 28354 12008 28410 12064
rect 28538 3032 28594 3088
rect 27250 1536 27306 1592
rect 28262 2252 28264 2272
rect 28264 2252 28316 2272
rect 28316 2252 28318 2272
rect 28262 2216 28318 2252
rect 28814 12280 28870 12336
rect 28906 12044 28908 12064
rect 28908 12044 28960 12064
rect 28960 12044 28962 12064
rect 28906 12008 28962 12044
rect 28814 11736 28870 11792
rect 28906 11056 28962 11112
rect 29642 13252 29698 13288
rect 29642 13232 29644 13252
rect 29644 13232 29696 13252
rect 29696 13232 29698 13252
rect 29550 12008 29606 12064
rect 30286 14864 30342 14920
rect 30562 15816 30618 15872
rect 30838 14184 30894 14240
rect 30930 13776 30986 13832
rect 30010 12144 30066 12200
rect 29826 11872 29882 11928
rect 29734 10920 29790 10976
rect 30746 11092 30748 11112
rect 30748 11092 30800 11112
rect 30800 11092 30802 11112
rect 30746 11056 30802 11092
rect 31206 27376 31262 27432
rect 31114 22616 31170 22672
rect 31114 17448 31170 17504
rect 33878 27770 33934 27772
rect 33958 27770 34014 27772
rect 34038 27770 34094 27772
rect 34118 27770 34174 27772
rect 33878 27718 33924 27770
rect 33924 27718 33934 27770
rect 33958 27718 33988 27770
rect 33988 27718 34000 27770
rect 34000 27718 34014 27770
rect 34038 27718 34052 27770
rect 34052 27718 34064 27770
rect 34064 27718 34094 27770
rect 34118 27718 34128 27770
rect 34128 27718 34174 27770
rect 33878 27716 33934 27718
rect 33958 27716 34014 27718
rect 34038 27716 34094 27718
rect 34118 27716 34174 27718
rect 33046 26424 33102 26480
rect 31758 17312 31814 17368
rect 31482 15136 31538 15192
rect 31942 15544 31998 15600
rect 31114 13796 31170 13832
rect 31114 13776 31116 13796
rect 31116 13776 31168 13796
rect 31168 13776 31170 13796
rect 31850 14456 31906 14512
rect 32770 17448 32826 17504
rect 32494 15544 32550 15600
rect 32402 14728 32458 14784
rect 32862 13640 32918 13696
rect 31758 11736 31814 11792
rect 31482 10804 31538 10840
rect 31482 10784 31484 10804
rect 31484 10784 31536 10804
rect 31536 10784 31538 10804
rect 30286 1944 30342 2000
rect 33138 15816 33194 15872
rect 33322 14864 33378 14920
rect 33322 14184 33378 14240
rect 33878 26682 33934 26684
rect 33958 26682 34014 26684
rect 34038 26682 34094 26684
rect 34118 26682 34174 26684
rect 33878 26630 33924 26682
rect 33924 26630 33934 26682
rect 33958 26630 33988 26682
rect 33988 26630 34000 26682
rect 34000 26630 34014 26682
rect 34038 26630 34052 26682
rect 34052 26630 34064 26682
rect 34064 26630 34094 26682
rect 34118 26630 34128 26682
rect 34128 26630 34174 26682
rect 33878 26628 33934 26630
rect 33958 26628 34014 26630
rect 34038 26628 34094 26630
rect 34118 26628 34174 26630
rect 33878 25594 33934 25596
rect 33958 25594 34014 25596
rect 34038 25594 34094 25596
rect 34118 25594 34174 25596
rect 33878 25542 33924 25594
rect 33924 25542 33934 25594
rect 33958 25542 33988 25594
rect 33988 25542 34000 25594
rect 34000 25542 34014 25594
rect 34038 25542 34052 25594
rect 34052 25542 34064 25594
rect 34064 25542 34094 25594
rect 34118 25542 34128 25594
rect 34128 25542 34174 25594
rect 33878 25540 33934 25542
rect 33958 25540 34014 25542
rect 34038 25540 34094 25542
rect 34118 25540 34174 25542
rect 33878 24506 33934 24508
rect 33958 24506 34014 24508
rect 34038 24506 34094 24508
rect 34118 24506 34174 24508
rect 33878 24454 33924 24506
rect 33924 24454 33934 24506
rect 33958 24454 33988 24506
rect 33988 24454 34000 24506
rect 34000 24454 34014 24506
rect 34038 24454 34052 24506
rect 34052 24454 34064 24506
rect 34064 24454 34094 24506
rect 34118 24454 34128 24506
rect 34128 24454 34174 24506
rect 33878 24452 33934 24454
rect 33958 24452 34014 24454
rect 34038 24452 34094 24454
rect 34118 24452 34174 24454
rect 33878 23418 33934 23420
rect 33958 23418 34014 23420
rect 34038 23418 34094 23420
rect 34118 23418 34174 23420
rect 33878 23366 33924 23418
rect 33924 23366 33934 23418
rect 33958 23366 33988 23418
rect 33988 23366 34000 23418
rect 34000 23366 34014 23418
rect 34038 23366 34052 23418
rect 34052 23366 34064 23418
rect 34064 23366 34094 23418
rect 34118 23366 34128 23418
rect 34128 23366 34174 23418
rect 33878 23364 33934 23366
rect 33958 23364 34014 23366
rect 34038 23364 34094 23366
rect 34118 23364 34174 23366
rect 33878 22330 33934 22332
rect 33958 22330 34014 22332
rect 34038 22330 34094 22332
rect 34118 22330 34174 22332
rect 33878 22278 33924 22330
rect 33924 22278 33934 22330
rect 33958 22278 33988 22330
rect 33988 22278 34000 22330
rect 34000 22278 34014 22330
rect 34038 22278 34052 22330
rect 34052 22278 34064 22330
rect 34064 22278 34094 22330
rect 34118 22278 34128 22330
rect 34128 22278 34174 22330
rect 33878 22276 33934 22278
rect 33958 22276 34014 22278
rect 34038 22276 34094 22278
rect 34118 22276 34174 22278
rect 33878 21242 33934 21244
rect 33958 21242 34014 21244
rect 34038 21242 34094 21244
rect 34118 21242 34174 21244
rect 33878 21190 33924 21242
rect 33924 21190 33934 21242
rect 33958 21190 33988 21242
rect 33988 21190 34000 21242
rect 34000 21190 34014 21242
rect 34038 21190 34052 21242
rect 34052 21190 34064 21242
rect 34064 21190 34094 21242
rect 34118 21190 34128 21242
rect 34128 21190 34174 21242
rect 33878 21188 33934 21190
rect 33958 21188 34014 21190
rect 34038 21188 34094 21190
rect 34118 21188 34174 21190
rect 33878 20154 33934 20156
rect 33958 20154 34014 20156
rect 34038 20154 34094 20156
rect 34118 20154 34174 20156
rect 33878 20102 33924 20154
rect 33924 20102 33934 20154
rect 33958 20102 33988 20154
rect 33988 20102 34000 20154
rect 34000 20102 34014 20154
rect 34038 20102 34052 20154
rect 34052 20102 34064 20154
rect 34064 20102 34094 20154
rect 34118 20102 34128 20154
rect 34128 20102 34174 20154
rect 33878 20100 33934 20102
rect 33958 20100 34014 20102
rect 34038 20100 34094 20102
rect 34118 20100 34174 20102
rect 33878 19066 33934 19068
rect 33958 19066 34014 19068
rect 34038 19066 34094 19068
rect 34118 19066 34174 19068
rect 33878 19014 33924 19066
rect 33924 19014 33934 19066
rect 33958 19014 33988 19066
rect 33988 19014 34000 19066
rect 34000 19014 34014 19066
rect 34038 19014 34052 19066
rect 34052 19014 34064 19066
rect 34064 19014 34094 19066
rect 34118 19014 34128 19066
rect 34128 19014 34174 19066
rect 33878 19012 33934 19014
rect 33958 19012 34014 19014
rect 34038 19012 34094 19014
rect 34118 19012 34174 19014
rect 33598 17196 33654 17232
rect 33598 17176 33600 17196
rect 33600 17176 33652 17196
rect 33652 17176 33654 17196
rect 33598 15680 33654 15736
rect 33506 14728 33562 14784
rect 33878 17978 33934 17980
rect 33958 17978 34014 17980
rect 34038 17978 34094 17980
rect 34118 17978 34174 17980
rect 33878 17926 33924 17978
rect 33924 17926 33934 17978
rect 33958 17926 33988 17978
rect 33988 17926 34000 17978
rect 34000 17926 34014 17978
rect 34038 17926 34052 17978
rect 34052 17926 34064 17978
rect 34064 17926 34094 17978
rect 34118 17926 34128 17978
rect 34128 17926 34174 17978
rect 33878 17924 33934 17926
rect 33958 17924 34014 17926
rect 34038 17924 34094 17926
rect 34118 17924 34174 17926
rect 33878 16890 33934 16892
rect 33958 16890 34014 16892
rect 34038 16890 34094 16892
rect 34118 16890 34174 16892
rect 33878 16838 33924 16890
rect 33924 16838 33934 16890
rect 33958 16838 33988 16890
rect 33988 16838 34000 16890
rect 34000 16838 34014 16890
rect 34038 16838 34052 16890
rect 34052 16838 34064 16890
rect 34064 16838 34094 16890
rect 34118 16838 34128 16890
rect 34128 16838 34174 16890
rect 33878 16836 33934 16838
rect 33958 16836 34014 16838
rect 34038 16836 34094 16838
rect 34118 16836 34174 16838
rect 34334 16496 34390 16552
rect 33878 15802 33934 15804
rect 33958 15802 34014 15804
rect 34038 15802 34094 15804
rect 34118 15802 34174 15804
rect 33878 15750 33924 15802
rect 33924 15750 33934 15802
rect 33958 15750 33988 15802
rect 33988 15750 34000 15802
rect 34000 15750 34014 15802
rect 34038 15750 34052 15802
rect 34052 15750 34064 15802
rect 34064 15750 34094 15802
rect 34118 15750 34128 15802
rect 34128 15750 34174 15802
rect 33878 15748 33934 15750
rect 33958 15748 34014 15750
rect 34038 15748 34094 15750
rect 34118 15748 34174 15750
rect 35070 17176 35126 17232
rect 33966 14864 34022 14920
rect 33878 14714 33934 14716
rect 33958 14714 34014 14716
rect 34038 14714 34094 14716
rect 34118 14714 34174 14716
rect 33878 14662 33924 14714
rect 33924 14662 33934 14714
rect 33958 14662 33988 14714
rect 33988 14662 34000 14714
rect 34000 14662 34014 14714
rect 34038 14662 34052 14714
rect 34052 14662 34064 14714
rect 34064 14662 34094 14714
rect 34118 14662 34128 14714
rect 34128 14662 34174 14714
rect 33878 14660 33934 14662
rect 33958 14660 34014 14662
rect 34038 14660 34094 14662
rect 34118 14660 34174 14662
rect 34242 14456 34298 14512
rect 33414 13796 33470 13832
rect 33414 13776 33416 13796
rect 33416 13776 33468 13796
rect 33468 13776 33470 13796
rect 33874 14048 33930 14104
rect 33230 12280 33286 12336
rect 32862 11600 32918 11656
rect 33322 12008 33378 12064
rect 33878 13626 33934 13628
rect 33958 13626 34014 13628
rect 34038 13626 34094 13628
rect 34118 13626 34174 13628
rect 33878 13574 33924 13626
rect 33924 13574 33934 13626
rect 33958 13574 33988 13626
rect 33988 13574 34000 13626
rect 34000 13574 34014 13626
rect 34038 13574 34052 13626
rect 34052 13574 34064 13626
rect 34064 13574 34094 13626
rect 34118 13574 34128 13626
rect 34128 13574 34174 13626
rect 33878 13572 33934 13574
rect 33958 13572 34014 13574
rect 34038 13572 34094 13574
rect 34118 13572 34174 13574
rect 34150 13096 34206 13152
rect 33878 12538 33934 12540
rect 33958 12538 34014 12540
rect 34038 12538 34094 12540
rect 34118 12538 34174 12540
rect 33878 12486 33924 12538
rect 33924 12486 33934 12538
rect 33958 12486 33988 12538
rect 33988 12486 34000 12538
rect 34000 12486 34014 12538
rect 34038 12486 34052 12538
rect 34052 12486 34064 12538
rect 34064 12486 34094 12538
rect 34118 12486 34128 12538
rect 34128 12486 34174 12538
rect 33878 12484 33934 12486
rect 33958 12484 34014 12486
rect 34038 12484 34094 12486
rect 34118 12484 34174 12486
rect 33874 11872 33930 11928
rect 33878 11450 33934 11452
rect 33958 11450 34014 11452
rect 34038 11450 34094 11452
rect 34118 11450 34174 11452
rect 33878 11398 33924 11450
rect 33924 11398 33934 11450
rect 33958 11398 33988 11450
rect 33988 11398 34000 11450
rect 34000 11398 34014 11450
rect 34038 11398 34052 11450
rect 34052 11398 34064 11450
rect 34064 11398 34094 11450
rect 34118 11398 34128 11450
rect 34128 11398 34174 11450
rect 33878 11396 33934 11398
rect 33958 11396 34014 11398
rect 34038 11396 34094 11398
rect 34118 11396 34174 11398
rect 34978 14356 34980 14376
rect 34980 14356 35032 14376
rect 35032 14356 35034 14376
rect 34978 14320 35034 14356
rect 34610 13524 34666 13560
rect 34610 13504 34612 13524
rect 34612 13504 34664 13524
rect 34664 13504 34666 13524
rect 34886 13640 34942 13696
rect 34334 11736 34390 11792
rect 33878 10362 33934 10364
rect 33958 10362 34014 10364
rect 34038 10362 34094 10364
rect 34118 10362 34174 10364
rect 33878 10310 33924 10362
rect 33924 10310 33934 10362
rect 33958 10310 33988 10362
rect 33988 10310 34000 10362
rect 34000 10310 34014 10362
rect 34038 10310 34052 10362
rect 34052 10310 34064 10362
rect 34064 10310 34094 10362
rect 34118 10310 34128 10362
rect 34128 10310 34174 10362
rect 33878 10308 33934 10310
rect 33958 10308 34014 10310
rect 34038 10308 34094 10310
rect 34118 10308 34174 10310
rect 33878 9274 33934 9276
rect 33958 9274 34014 9276
rect 34038 9274 34094 9276
rect 34118 9274 34174 9276
rect 33878 9222 33924 9274
rect 33924 9222 33934 9274
rect 33958 9222 33988 9274
rect 33988 9222 34000 9274
rect 34000 9222 34014 9274
rect 34038 9222 34052 9274
rect 34052 9222 34064 9274
rect 34064 9222 34094 9274
rect 34118 9222 34128 9274
rect 34128 9222 34174 9274
rect 33878 9220 33934 9222
rect 33958 9220 34014 9222
rect 34038 9220 34094 9222
rect 34118 9220 34174 9222
rect 33878 8186 33934 8188
rect 33958 8186 34014 8188
rect 34038 8186 34094 8188
rect 34118 8186 34174 8188
rect 33878 8134 33924 8186
rect 33924 8134 33934 8186
rect 33958 8134 33988 8186
rect 33988 8134 34000 8186
rect 34000 8134 34014 8186
rect 34038 8134 34052 8186
rect 34052 8134 34064 8186
rect 34064 8134 34094 8186
rect 34118 8134 34128 8186
rect 34128 8134 34174 8186
rect 33878 8132 33934 8134
rect 33958 8132 34014 8134
rect 34038 8132 34094 8134
rect 34118 8132 34174 8134
rect 33878 7098 33934 7100
rect 33958 7098 34014 7100
rect 34038 7098 34094 7100
rect 34118 7098 34174 7100
rect 33878 7046 33924 7098
rect 33924 7046 33934 7098
rect 33958 7046 33988 7098
rect 33988 7046 34000 7098
rect 34000 7046 34014 7098
rect 34038 7046 34052 7098
rect 34052 7046 34064 7098
rect 34064 7046 34094 7098
rect 34118 7046 34128 7098
rect 34128 7046 34174 7098
rect 33878 7044 33934 7046
rect 33958 7044 34014 7046
rect 34038 7044 34094 7046
rect 34118 7044 34174 7046
rect 35254 14048 35310 14104
rect 35070 12008 35126 12064
rect 35254 12008 35310 12064
rect 33878 6010 33934 6012
rect 33958 6010 34014 6012
rect 34038 6010 34094 6012
rect 34118 6010 34174 6012
rect 33878 5958 33924 6010
rect 33924 5958 33934 6010
rect 33958 5958 33988 6010
rect 33988 5958 34000 6010
rect 34000 5958 34014 6010
rect 34038 5958 34052 6010
rect 34052 5958 34064 6010
rect 34064 5958 34094 6010
rect 34118 5958 34128 6010
rect 34128 5958 34174 6010
rect 33878 5956 33934 5958
rect 33958 5956 34014 5958
rect 34038 5956 34094 5958
rect 34118 5956 34174 5958
rect 33878 4922 33934 4924
rect 33958 4922 34014 4924
rect 34038 4922 34094 4924
rect 34118 4922 34174 4924
rect 33878 4870 33924 4922
rect 33924 4870 33934 4922
rect 33958 4870 33988 4922
rect 33988 4870 34000 4922
rect 34000 4870 34014 4922
rect 34038 4870 34052 4922
rect 34052 4870 34064 4922
rect 34064 4870 34094 4922
rect 34118 4870 34128 4922
rect 34128 4870 34174 4922
rect 33878 4868 33934 4870
rect 33958 4868 34014 4870
rect 34038 4868 34094 4870
rect 34118 4868 34174 4870
rect 33878 3834 33934 3836
rect 33958 3834 34014 3836
rect 34038 3834 34094 3836
rect 34118 3834 34174 3836
rect 33878 3782 33924 3834
rect 33924 3782 33934 3834
rect 33958 3782 33988 3834
rect 33988 3782 34000 3834
rect 34000 3782 34014 3834
rect 34038 3782 34052 3834
rect 34052 3782 34064 3834
rect 34064 3782 34094 3834
rect 34118 3782 34128 3834
rect 34128 3782 34174 3834
rect 33878 3780 33934 3782
rect 33958 3780 34014 3782
rect 34038 3780 34094 3782
rect 34118 3780 34174 3782
rect 31850 1944 31906 2000
rect 31666 1844 31668 1864
rect 31668 1844 31720 1864
rect 31720 1844 31722 1864
rect 31666 1808 31722 1844
rect 31758 1672 31814 1728
rect 31850 1556 31906 1592
rect 31850 1536 31852 1556
rect 31852 1536 31904 1556
rect 31904 1536 31906 1556
rect 33878 2746 33934 2748
rect 33958 2746 34014 2748
rect 34038 2746 34094 2748
rect 34118 2746 34174 2748
rect 33878 2694 33924 2746
rect 33924 2694 33934 2746
rect 33958 2694 33988 2746
rect 33988 2694 34000 2746
rect 34000 2694 34014 2746
rect 34038 2694 34052 2746
rect 34052 2694 34064 2746
rect 34064 2694 34094 2746
rect 34118 2694 34128 2746
rect 34128 2694 34174 2746
rect 33878 2692 33934 2694
rect 33958 2692 34014 2694
rect 34038 2692 34094 2694
rect 34118 2692 34174 2694
rect 36450 18300 36452 18320
rect 36452 18300 36504 18320
rect 36504 18300 36506 18320
rect 36450 18264 36506 18300
rect 37646 17196 37702 17232
rect 37646 17176 37648 17196
rect 37648 17176 37700 17196
rect 37700 17176 37702 17196
rect 35806 14048 35862 14104
rect 35714 13504 35770 13560
rect 35530 12824 35586 12880
rect 35438 12144 35494 12200
rect 35438 11736 35494 11792
rect 36174 15136 36230 15192
rect 36266 14900 36268 14920
rect 36268 14900 36320 14920
rect 36320 14900 36322 14920
rect 36266 14864 36322 14900
rect 35806 11872 35862 11928
rect 35806 11600 35862 11656
rect 36266 12044 36268 12064
rect 36268 12044 36320 12064
rect 36320 12044 36322 12064
rect 36266 12008 36322 12044
rect 36266 11636 36268 11656
rect 36268 11636 36320 11656
rect 36320 11636 36322 11656
rect 36266 11600 36322 11636
rect 34058 2080 34114 2136
rect 36634 14320 36690 14376
rect 36450 13640 36506 13696
rect 37002 14220 37004 14240
rect 37004 14220 37056 14240
rect 37056 14220 37058 14240
rect 37002 14184 37058 14220
rect 37002 13776 37058 13832
rect 36910 13132 36912 13152
rect 36912 13132 36964 13152
rect 36964 13132 36966 13152
rect 36910 13096 36966 13132
rect 37370 14864 37426 14920
rect 37370 14184 37426 14240
rect 37278 14048 37334 14104
rect 37278 13096 37334 13152
rect 37186 12144 37242 12200
rect 36726 11756 36782 11792
rect 36726 11736 36728 11756
rect 36728 11736 36780 11756
rect 36780 11736 36782 11756
rect 37094 11192 37150 11248
rect 37094 10784 37150 10840
rect 37554 13796 37610 13832
rect 37554 13776 37556 13796
rect 37556 13776 37608 13796
rect 37608 13776 37610 13796
rect 38198 26832 38254 26888
rect 38750 16652 38806 16688
rect 38750 16632 38752 16652
rect 38752 16632 38804 16652
rect 38804 16632 38806 16652
rect 37922 14864 37978 14920
rect 39302 15136 39358 15192
rect 38290 14356 38292 14376
rect 38292 14356 38344 14376
rect 38344 14356 38346 14376
rect 38290 14320 38346 14356
rect 37738 11872 37794 11928
rect 37738 10956 37740 10976
rect 37740 10956 37792 10976
rect 37792 10956 37794 10976
rect 37738 10920 37794 10956
rect 39578 16768 39634 16824
rect 38750 13504 38806 13560
rect 39394 13640 39450 13696
rect 38566 12280 38622 12336
rect 38290 11328 38346 11384
rect 38106 11092 38108 11112
rect 38108 11092 38160 11112
rect 38160 11092 38162 11112
rect 38106 11056 38162 11092
rect 38566 10512 38622 10568
rect 39394 13504 39450 13560
rect 38842 12280 38898 12336
rect 39026 12008 39082 12064
rect 38934 11192 38990 11248
rect 38842 10784 38898 10840
rect 38658 9988 38714 10024
rect 38658 9968 38660 9988
rect 38660 9968 38712 9988
rect 38712 9968 38714 9988
rect 40682 26968 40738 27024
rect 40682 26324 40684 26344
rect 40684 26324 40736 26344
rect 40736 26324 40738 26344
rect 40682 26288 40738 26324
rect 40682 17856 40738 17912
rect 40498 17176 40554 17232
rect 39946 14456 40002 14512
rect 40130 13776 40186 13832
rect 40314 13796 40370 13832
rect 40314 13776 40316 13796
rect 40316 13776 40368 13796
rect 40368 13776 40370 13796
rect 39394 11736 39450 11792
rect 39486 10784 39542 10840
rect 40038 12180 40040 12200
rect 40040 12180 40092 12200
rect 40092 12180 40094 12200
rect 40038 12144 40094 12180
rect 40590 13096 40646 13152
rect 39118 9968 39174 10024
rect 35714 1672 35770 1728
rect 38658 1808 38714 1864
rect 39946 2896 40002 2952
rect 40774 15136 40830 15192
rect 41510 17720 41566 17776
rect 41326 17448 41382 17504
rect 42614 27396 42670 27432
rect 42614 27376 42616 27396
rect 42616 27376 42668 27396
rect 42668 27376 42670 27396
rect 41786 26968 41842 27024
rect 42706 26968 42762 27024
rect 41694 26288 41750 26344
rect 41694 17484 41696 17504
rect 41696 17484 41748 17504
rect 41748 17484 41750 17504
rect 41694 17448 41750 17484
rect 41602 14592 41658 14648
rect 41418 14184 41474 14240
rect 41510 14068 41566 14104
rect 41510 14048 41512 14068
rect 41512 14048 41564 14068
rect 41564 14048 41566 14068
rect 41786 14456 41842 14512
rect 41694 13776 41750 13832
rect 40958 13640 41014 13696
rect 40958 13096 41014 13152
rect 41326 13640 41382 13696
rect 41786 12824 41842 12880
rect 41510 12688 41566 12744
rect 41694 12144 41750 12200
rect 42154 22616 42210 22672
rect 42246 17720 42302 17776
rect 42338 17040 42394 17096
rect 42338 16768 42394 16824
rect 42982 16668 42984 16688
rect 42984 16668 43036 16688
rect 43036 16668 43038 16688
rect 42982 16632 43038 16668
rect 42614 15680 42670 15736
rect 42890 15816 42946 15872
rect 42798 14864 42854 14920
rect 42890 14764 42892 14784
rect 42892 14764 42944 14784
rect 42944 14764 42946 14784
rect 42890 14728 42946 14764
rect 41142 11212 41198 11248
rect 41142 11192 41144 11212
rect 41144 11192 41196 11212
rect 41196 11192 41198 11212
rect 41142 10956 41144 10976
rect 41144 10956 41196 10976
rect 41196 10956 41198 10976
rect 41142 10920 41198 10956
rect 41418 10512 41474 10568
rect 40958 2760 41014 2816
rect 40314 2080 40370 2136
rect 42154 10240 42210 10296
rect 42890 13504 42946 13560
rect 42798 12824 42854 12880
rect 42614 3732 42670 3768
rect 42614 3712 42616 3732
rect 42616 3712 42668 3732
rect 42668 3712 42670 3732
rect 44852 27226 44908 27228
rect 44932 27226 44988 27228
rect 45012 27226 45068 27228
rect 45092 27226 45148 27228
rect 44852 27174 44898 27226
rect 44898 27174 44908 27226
rect 44932 27174 44962 27226
rect 44962 27174 44974 27226
rect 44974 27174 44988 27226
rect 45012 27174 45026 27226
rect 45026 27174 45038 27226
rect 45038 27174 45068 27226
rect 45092 27174 45102 27226
rect 45102 27174 45148 27226
rect 44852 27172 44908 27174
rect 44932 27172 44988 27174
rect 45012 27172 45068 27174
rect 45092 27172 45148 27174
rect 44822 26988 44878 27024
rect 44822 26968 44824 26988
rect 44824 26968 44876 26988
rect 44876 26968 44878 26988
rect 43442 17740 43498 17776
rect 43442 17720 43444 17740
rect 43444 17720 43496 17740
rect 43496 17720 43498 17740
rect 43902 15816 43958 15872
rect 43902 14592 43958 14648
rect 43442 12960 43498 13016
rect 43350 11872 43406 11928
rect 43810 13640 43866 13696
rect 44852 26138 44908 26140
rect 44932 26138 44988 26140
rect 45012 26138 45068 26140
rect 45092 26138 45148 26140
rect 44852 26086 44898 26138
rect 44898 26086 44908 26138
rect 44932 26086 44962 26138
rect 44962 26086 44974 26138
rect 44974 26086 44988 26138
rect 45012 26086 45026 26138
rect 45026 26086 45038 26138
rect 45038 26086 45068 26138
rect 45092 26086 45102 26138
rect 45102 26086 45148 26138
rect 44852 26084 44908 26086
rect 44932 26084 44988 26086
rect 45012 26084 45068 26086
rect 45092 26084 45148 26086
rect 44270 15544 44326 15600
rect 44852 25050 44908 25052
rect 44932 25050 44988 25052
rect 45012 25050 45068 25052
rect 45092 25050 45148 25052
rect 44852 24998 44898 25050
rect 44898 24998 44908 25050
rect 44932 24998 44962 25050
rect 44962 24998 44974 25050
rect 44974 24998 44988 25050
rect 45012 24998 45026 25050
rect 45026 24998 45038 25050
rect 45038 24998 45068 25050
rect 45092 24998 45102 25050
rect 45102 24998 45148 25050
rect 44852 24996 44908 24998
rect 44932 24996 44988 24998
rect 45012 24996 45068 24998
rect 45092 24996 45148 24998
rect 44852 23962 44908 23964
rect 44932 23962 44988 23964
rect 45012 23962 45068 23964
rect 45092 23962 45148 23964
rect 44852 23910 44898 23962
rect 44898 23910 44908 23962
rect 44932 23910 44962 23962
rect 44962 23910 44974 23962
rect 44974 23910 44988 23962
rect 45012 23910 45026 23962
rect 45026 23910 45038 23962
rect 45038 23910 45068 23962
rect 45092 23910 45102 23962
rect 45102 23910 45148 23962
rect 44852 23908 44908 23910
rect 44932 23908 44988 23910
rect 45012 23908 45068 23910
rect 45092 23908 45148 23910
rect 44852 22874 44908 22876
rect 44932 22874 44988 22876
rect 45012 22874 45068 22876
rect 45092 22874 45148 22876
rect 44852 22822 44898 22874
rect 44898 22822 44908 22874
rect 44932 22822 44962 22874
rect 44962 22822 44974 22874
rect 44974 22822 44988 22874
rect 45012 22822 45026 22874
rect 45026 22822 45038 22874
rect 45038 22822 45068 22874
rect 45092 22822 45102 22874
rect 45102 22822 45148 22874
rect 44852 22820 44908 22822
rect 44932 22820 44988 22822
rect 45012 22820 45068 22822
rect 45092 22820 45148 22822
rect 44852 21786 44908 21788
rect 44932 21786 44988 21788
rect 45012 21786 45068 21788
rect 45092 21786 45148 21788
rect 44852 21734 44898 21786
rect 44898 21734 44908 21786
rect 44932 21734 44962 21786
rect 44962 21734 44974 21786
rect 44974 21734 44988 21786
rect 45012 21734 45026 21786
rect 45026 21734 45038 21786
rect 45038 21734 45068 21786
rect 45092 21734 45102 21786
rect 45102 21734 45148 21786
rect 44852 21732 44908 21734
rect 44932 21732 44988 21734
rect 45012 21732 45068 21734
rect 45092 21732 45148 21734
rect 44852 20698 44908 20700
rect 44932 20698 44988 20700
rect 45012 20698 45068 20700
rect 45092 20698 45148 20700
rect 44852 20646 44898 20698
rect 44898 20646 44908 20698
rect 44932 20646 44962 20698
rect 44962 20646 44974 20698
rect 44974 20646 44988 20698
rect 45012 20646 45026 20698
rect 45026 20646 45038 20698
rect 45038 20646 45068 20698
rect 45092 20646 45102 20698
rect 45102 20646 45148 20698
rect 44852 20644 44908 20646
rect 44932 20644 44988 20646
rect 45012 20644 45068 20646
rect 45092 20644 45148 20646
rect 44852 19610 44908 19612
rect 44932 19610 44988 19612
rect 45012 19610 45068 19612
rect 45092 19610 45148 19612
rect 44852 19558 44898 19610
rect 44898 19558 44908 19610
rect 44932 19558 44962 19610
rect 44962 19558 44974 19610
rect 44974 19558 44988 19610
rect 45012 19558 45026 19610
rect 45026 19558 45038 19610
rect 45038 19558 45068 19610
rect 45092 19558 45102 19610
rect 45102 19558 45148 19610
rect 44852 19556 44908 19558
rect 44932 19556 44988 19558
rect 45012 19556 45068 19558
rect 45092 19556 45148 19558
rect 44852 18522 44908 18524
rect 44932 18522 44988 18524
rect 45012 18522 45068 18524
rect 45092 18522 45148 18524
rect 44852 18470 44898 18522
rect 44898 18470 44908 18522
rect 44932 18470 44962 18522
rect 44962 18470 44974 18522
rect 44974 18470 44988 18522
rect 45012 18470 45026 18522
rect 45026 18470 45038 18522
rect 45038 18470 45068 18522
rect 45092 18470 45102 18522
rect 45102 18470 45148 18522
rect 44852 18468 44908 18470
rect 44932 18468 44988 18470
rect 45012 18468 45068 18470
rect 45092 18468 45148 18470
rect 44852 17434 44908 17436
rect 44932 17434 44988 17436
rect 45012 17434 45068 17436
rect 45092 17434 45148 17436
rect 44852 17382 44898 17434
rect 44898 17382 44908 17434
rect 44932 17382 44962 17434
rect 44962 17382 44974 17434
rect 44974 17382 44988 17434
rect 45012 17382 45026 17434
rect 45026 17382 45038 17434
rect 45038 17382 45068 17434
rect 45092 17382 45102 17434
rect 45102 17382 45148 17434
rect 44852 17380 44908 17382
rect 44932 17380 44988 17382
rect 45012 17380 45068 17382
rect 45092 17380 45148 17382
rect 46754 27396 46810 27432
rect 46754 27376 46756 27396
rect 46756 27376 46808 27396
rect 46808 27376 46810 27396
rect 45650 17856 45706 17912
rect 46294 17720 46350 17776
rect 45650 17312 45706 17368
rect 44730 16632 44786 16688
rect 44852 16346 44908 16348
rect 44932 16346 44988 16348
rect 45012 16346 45068 16348
rect 45092 16346 45148 16348
rect 44852 16294 44898 16346
rect 44898 16294 44908 16346
rect 44932 16294 44962 16346
rect 44962 16294 44974 16346
rect 44974 16294 44988 16346
rect 45012 16294 45026 16346
rect 45026 16294 45038 16346
rect 45038 16294 45068 16346
rect 45092 16294 45102 16346
rect 45102 16294 45148 16346
rect 44852 16292 44908 16294
rect 44932 16292 44988 16294
rect 45012 16292 45068 16294
rect 45092 16292 45148 16294
rect 46294 17584 46350 17640
rect 46754 17584 46810 17640
rect 45926 16904 45982 16960
rect 46202 16360 46258 16416
rect 44852 15258 44908 15260
rect 44932 15258 44988 15260
rect 45012 15258 45068 15260
rect 45092 15258 45148 15260
rect 44852 15206 44898 15258
rect 44898 15206 44908 15258
rect 44932 15206 44962 15258
rect 44962 15206 44974 15258
rect 44974 15206 44988 15258
rect 45012 15206 45026 15258
rect 45026 15206 45038 15258
rect 45038 15206 45068 15258
rect 45092 15206 45102 15258
rect 45102 15206 45148 15258
rect 44852 15204 44908 15206
rect 44932 15204 44988 15206
rect 45012 15204 45068 15206
rect 45092 15204 45148 15206
rect 44638 15136 44694 15192
rect 44086 13504 44142 13560
rect 44546 14184 44602 14240
rect 43902 13096 43958 13152
rect 43626 12280 43682 12336
rect 43718 11464 43774 11520
rect 43718 11192 43774 11248
rect 43350 10104 43406 10160
rect 43442 4004 43498 4040
rect 43442 3984 43444 4004
rect 43444 3984 43496 4004
rect 43496 3984 43498 4004
rect 43442 3476 43444 3496
rect 43444 3476 43496 3496
rect 43496 3476 43498 3496
rect 43442 3440 43498 3476
rect 43994 12008 44050 12064
rect 44362 11192 44418 11248
rect 44852 14170 44908 14172
rect 44932 14170 44988 14172
rect 45012 14170 45068 14172
rect 45092 14170 45148 14172
rect 44852 14118 44898 14170
rect 44898 14118 44908 14170
rect 44932 14118 44962 14170
rect 44962 14118 44974 14170
rect 44974 14118 44988 14170
rect 45012 14118 45026 14170
rect 45026 14118 45038 14170
rect 45038 14118 45068 14170
rect 45092 14118 45102 14170
rect 45102 14118 45148 14170
rect 44852 14116 44908 14118
rect 44932 14116 44988 14118
rect 45012 14116 45068 14118
rect 45092 14116 45148 14118
rect 45282 14048 45338 14104
rect 44730 13504 44786 13560
rect 44852 13082 44908 13084
rect 44932 13082 44988 13084
rect 45012 13082 45068 13084
rect 45092 13082 45148 13084
rect 44852 13030 44898 13082
rect 44898 13030 44908 13082
rect 44932 13030 44962 13082
rect 44962 13030 44974 13082
rect 44974 13030 44988 13082
rect 45012 13030 45026 13082
rect 45026 13030 45038 13082
rect 45038 13030 45068 13082
rect 45092 13030 45102 13082
rect 45102 13030 45148 13082
rect 44852 13028 44908 13030
rect 44932 13028 44988 13030
rect 45012 13028 45068 13030
rect 45092 13028 45148 13030
rect 45282 12824 45338 12880
rect 45558 13504 45614 13560
rect 45466 12960 45522 13016
rect 44852 11994 44908 11996
rect 44932 11994 44988 11996
rect 45012 11994 45068 11996
rect 45092 11994 45148 11996
rect 44852 11942 44898 11994
rect 44898 11942 44908 11994
rect 44932 11942 44962 11994
rect 44962 11942 44974 11994
rect 44974 11942 44988 11994
rect 45012 11942 45026 11994
rect 45026 11942 45038 11994
rect 45038 11942 45068 11994
rect 45092 11942 45102 11994
rect 45102 11942 45148 11994
rect 44852 11940 44908 11942
rect 44932 11940 44988 11942
rect 45012 11940 45068 11942
rect 45092 11940 45148 11942
rect 44822 11056 44878 11112
rect 44852 10906 44908 10908
rect 44932 10906 44988 10908
rect 45012 10906 45068 10908
rect 45092 10906 45148 10908
rect 44852 10854 44898 10906
rect 44898 10854 44908 10906
rect 44932 10854 44962 10906
rect 44962 10854 44974 10906
rect 44974 10854 44988 10906
rect 45012 10854 45026 10906
rect 45026 10854 45038 10906
rect 45038 10854 45068 10906
rect 45092 10854 45102 10906
rect 45102 10854 45148 10906
rect 44852 10852 44908 10854
rect 44932 10852 44988 10854
rect 45012 10852 45068 10854
rect 45092 10852 45148 10854
rect 46662 16224 46718 16280
rect 46386 16108 46442 16144
rect 46386 16088 46388 16108
rect 46388 16088 46440 16108
rect 46440 16088 46442 16108
rect 48134 17620 48136 17640
rect 48136 17620 48188 17640
rect 48188 17620 48190 17640
rect 48134 17584 48190 17620
rect 47858 17176 47914 17232
rect 48134 16768 48190 16824
rect 48870 17448 48926 17504
rect 48686 17312 48742 17368
rect 48410 16632 48466 16688
rect 47582 16532 47584 16552
rect 47584 16532 47636 16552
rect 47636 16532 47638 16552
rect 47582 16496 47638 16532
rect 48134 16496 48190 16552
rect 46846 15816 46902 15872
rect 46846 15136 46902 15192
rect 46938 14884 46994 14920
rect 46938 14864 46940 14884
rect 46940 14864 46992 14884
rect 46992 14864 46994 14884
rect 46662 14728 46718 14784
rect 46478 14320 46534 14376
rect 46018 13640 46074 13696
rect 45834 13096 45890 13152
rect 45926 12688 45982 12744
rect 46110 12688 46166 12744
rect 46846 12960 46902 13016
rect 46570 12552 46626 12608
rect 46386 12144 46442 12200
rect 45282 10512 45338 10568
rect 45834 11056 45890 11112
rect 45190 10376 45246 10432
rect 44852 9818 44908 9820
rect 44932 9818 44988 9820
rect 45012 9818 45068 9820
rect 45092 9818 45148 9820
rect 44852 9766 44898 9818
rect 44898 9766 44908 9818
rect 44932 9766 44962 9818
rect 44962 9766 44974 9818
rect 44974 9766 44988 9818
rect 45012 9766 45026 9818
rect 45026 9766 45038 9818
rect 45038 9766 45068 9818
rect 45092 9766 45102 9818
rect 45102 9766 45148 9818
rect 44852 9764 44908 9766
rect 44932 9764 44988 9766
rect 45012 9764 45068 9766
rect 45092 9764 45148 9766
rect 44852 8730 44908 8732
rect 44932 8730 44988 8732
rect 45012 8730 45068 8732
rect 45092 8730 45148 8732
rect 44852 8678 44898 8730
rect 44898 8678 44908 8730
rect 44932 8678 44962 8730
rect 44962 8678 44974 8730
rect 44974 8678 44988 8730
rect 45012 8678 45026 8730
rect 45026 8678 45038 8730
rect 45038 8678 45068 8730
rect 45092 8678 45102 8730
rect 45102 8678 45148 8730
rect 44852 8676 44908 8678
rect 44932 8676 44988 8678
rect 45012 8676 45068 8678
rect 45092 8676 45148 8678
rect 44852 7642 44908 7644
rect 44932 7642 44988 7644
rect 45012 7642 45068 7644
rect 45092 7642 45148 7644
rect 44852 7590 44898 7642
rect 44898 7590 44908 7642
rect 44932 7590 44962 7642
rect 44962 7590 44974 7642
rect 44974 7590 44988 7642
rect 45012 7590 45026 7642
rect 45026 7590 45038 7642
rect 45038 7590 45068 7642
rect 45092 7590 45102 7642
rect 45102 7590 45148 7642
rect 44852 7588 44908 7590
rect 44932 7588 44988 7590
rect 45012 7588 45068 7590
rect 45092 7588 45148 7590
rect 44852 6554 44908 6556
rect 44932 6554 44988 6556
rect 45012 6554 45068 6556
rect 45092 6554 45148 6556
rect 44852 6502 44898 6554
rect 44898 6502 44908 6554
rect 44932 6502 44962 6554
rect 44962 6502 44974 6554
rect 44974 6502 44988 6554
rect 45012 6502 45026 6554
rect 45026 6502 45038 6554
rect 45038 6502 45068 6554
rect 45092 6502 45102 6554
rect 45102 6502 45148 6554
rect 44852 6500 44908 6502
rect 44932 6500 44988 6502
rect 45012 6500 45068 6502
rect 45092 6500 45148 6502
rect 44852 5466 44908 5468
rect 44932 5466 44988 5468
rect 45012 5466 45068 5468
rect 45092 5466 45148 5468
rect 44852 5414 44898 5466
rect 44898 5414 44908 5466
rect 44932 5414 44962 5466
rect 44962 5414 44974 5466
rect 44974 5414 44988 5466
rect 45012 5414 45026 5466
rect 45026 5414 45038 5466
rect 45038 5414 45068 5466
rect 45092 5414 45102 5466
rect 45102 5414 45148 5466
rect 44852 5412 44908 5414
rect 44932 5412 44988 5414
rect 45012 5412 45068 5414
rect 45092 5412 45148 5414
rect 44852 4378 44908 4380
rect 44932 4378 44988 4380
rect 45012 4378 45068 4380
rect 45092 4378 45148 4380
rect 44852 4326 44898 4378
rect 44898 4326 44908 4378
rect 44932 4326 44962 4378
rect 44962 4326 44974 4378
rect 44974 4326 44988 4378
rect 45012 4326 45026 4378
rect 45026 4326 45038 4378
rect 45038 4326 45068 4378
rect 45092 4326 45102 4378
rect 45102 4326 45148 4378
rect 44852 4324 44908 4326
rect 44932 4324 44988 4326
rect 45012 4324 45068 4326
rect 45092 4324 45148 4326
rect 44852 3290 44908 3292
rect 44932 3290 44988 3292
rect 45012 3290 45068 3292
rect 45092 3290 45148 3292
rect 44852 3238 44898 3290
rect 44898 3238 44908 3290
rect 44932 3238 44962 3290
rect 44962 3238 44974 3290
rect 44974 3238 44988 3290
rect 45012 3238 45026 3290
rect 45026 3238 45038 3290
rect 45038 3238 45068 3290
rect 45092 3238 45102 3290
rect 45102 3238 45148 3290
rect 44852 3236 44908 3238
rect 44932 3236 44988 3238
rect 45012 3236 45068 3238
rect 45092 3236 45148 3238
rect 45282 2896 45338 2952
rect 45466 2896 45522 2952
rect 45558 2760 45614 2816
rect 44852 2202 44908 2204
rect 44932 2202 44988 2204
rect 45012 2202 45068 2204
rect 45092 2202 45148 2204
rect 44852 2150 44898 2202
rect 44898 2150 44908 2202
rect 44932 2150 44962 2202
rect 44962 2150 44974 2202
rect 44974 2150 44988 2202
rect 45012 2150 45026 2202
rect 45026 2150 45038 2202
rect 45038 2150 45068 2202
rect 45092 2150 45102 2202
rect 45102 2150 45148 2202
rect 44852 2148 44908 2150
rect 44932 2148 44988 2150
rect 45012 2148 45068 2150
rect 45092 2148 45148 2150
rect 45558 1980 45560 2000
rect 45560 1980 45612 2000
rect 45612 1980 45614 2000
rect 45558 1944 45614 1980
rect 45558 1692 45614 1728
rect 45558 1672 45560 1692
rect 45560 1672 45612 1692
rect 45612 1672 45614 1692
rect 46478 4004 46534 4040
rect 46478 3984 46480 4004
rect 46480 3984 46532 4004
rect 46532 3984 46534 4004
rect 47122 12552 47178 12608
rect 46754 12008 46810 12064
rect 46754 11872 46810 11928
rect 47122 11328 47178 11384
rect 47306 11328 47362 11384
rect 46754 10512 46810 10568
rect 47214 10412 47216 10432
rect 47216 10412 47268 10432
rect 47268 10412 47270 10432
rect 47214 10376 47270 10412
rect 48042 16360 48098 16416
rect 48226 16224 48282 16280
rect 48226 15700 48282 15736
rect 48226 15680 48228 15700
rect 48228 15680 48280 15700
rect 48280 15680 48282 15700
rect 48502 15680 48558 15736
rect 48042 15544 48098 15600
rect 48318 15272 48374 15328
rect 48778 15272 48834 15328
rect 48410 14728 48466 14784
rect 47674 14456 47730 14512
rect 47490 14220 47492 14240
rect 47492 14220 47544 14240
rect 47544 14220 47546 14240
rect 47490 14184 47546 14220
rect 47858 13776 47914 13832
rect 48318 13776 48374 13832
rect 48226 13504 48282 13560
rect 48134 12416 48190 12472
rect 48410 12824 48466 12880
rect 48042 12008 48098 12064
rect 48410 12416 48466 12472
rect 48410 12008 48466 12064
rect 48870 14900 48872 14920
rect 48872 14900 48924 14920
rect 48924 14900 48926 14920
rect 48870 14864 48926 14900
rect 48686 12416 48742 12472
rect 48502 11464 48558 11520
rect 47858 10104 47914 10160
rect 46570 2760 46626 2816
rect 48226 3712 48282 3768
rect 48134 3440 48190 3496
rect 48870 13504 48926 13560
rect 49422 17176 49478 17232
rect 49698 17312 49754 17368
rect 50066 17312 50122 17368
rect 49606 16224 49662 16280
rect 49422 15816 49478 15872
rect 49238 13640 49294 13696
rect 49238 13504 49294 13560
rect 48870 12008 48926 12064
rect 49238 11464 49294 11520
rect 48870 3476 48872 3496
rect 48872 3476 48924 3496
rect 48924 3476 48926 3496
rect 48870 3440 48926 3476
rect 45834 1808 45890 1864
rect 48870 1980 48872 2000
rect 48872 1980 48924 2000
rect 48924 1980 48926 2000
rect 48870 1944 48926 1980
rect 48502 1672 48558 1728
rect 49238 3168 49294 3224
rect 49974 17060 50030 17096
rect 49974 17040 49976 17060
rect 49976 17040 50028 17060
rect 50028 17040 50030 17060
rect 50250 16768 50306 16824
rect 49422 13096 49478 13152
rect 49606 13096 49662 13152
rect 49514 12960 49570 13016
rect 50158 15816 50214 15872
rect 49974 15544 50030 15600
rect 50526 18128 50582 18184
rect 50618 16632 50674 16688
rect 50434 14340 50490 14376
rect 50434 14320 50436 14340
rect 50436 14320 50488 14340
rect 50488 14320 50490 14340
rect 50342 14048 50398 14104
rect 50986 16940 50988 16960
rect 50988 16940 51040 16960
rect 51040 16940 51042 16960
rect 50986 16904 51042 16940
rect 51354 16360 51410 16416
rect 51170 15952 51226 16008
rect 51078 15272 51134 15328
rect 50986 15136 51042 15192
rect 50618 14592 50674 14648
rect 50894 14612 50950 14648
rect 50894 14592 50896 14612
rect 50896 14592 50948 14612
rect 50948 14592 50950 14612
rect 50618 14220 50620 14240
rect 50620 14220 50672 14240
rect 50672 14220 50674 14240
rect 50618 14184 50674 14220
rect 50802 14184 50858 14240
rect 50158 13504 50214 13560
rect 49606 11056 49662 11112
rect 49514 10784 49570 10840
rect 50158 12724 50160 12744
rect 50160 12724 50212 12744
rect 50212 12724 50214 12744
rect 50158 12688 50214 12724
rect 49974 12280 50030 12336
rect 50434 12300 50490 12336
rect 50434 12280 50436 12300
rect 50436 12280 50488 12300
rect 50488 12280 50490 12300
rect 49514 3460 49570 3496
rect 49514 3440 49516 3460
rect 49516 3440 49568 3460
rect 49568 3440 49570 3460
rect 49790 2896 49846 2952
rect 50250 3304 50306 3360
rect 50986 13504 51042 13560
rect 50894 12960 50950 13016
rect 51170 13504 51226 13560
rect 51446 15272 51502 15328
rect 51354 14592 51410 14648
rect 51538 14592 51594 14648
rect 51630 14456 51686 14512
rect 51906 16768 51962 16824
rect 51998 15544 52054 15600
rect 51170 13232 51226 13288
rect 51538 13232 51594 13288
rect 51354 12008 51410 12064
rect 51354 11500 51356 11520
rect 51356 11500 51408 11520
rect 51408 11500 51410 11520
rect 51354 11464 51410 11500
rect 50894 10920 50950 10976
rect 50802 10104 50858 10160
rect 51354 10920 51410 10976
rect 53010 17584 53066 17640
rect 52274 15544 52330 15600
rect 52274 14864 52330 14920
rect 52182 14320 52238 14376
rect 52826 16496 52882 16552
rect 53194 16244 53250 16280
rect 53194 16224 53196 16244
rect 53196 16224 53248 16244
rect 53248 16224 53250 16244
rect 52826 15952 52882 16008
rect 52550 15272 52606 15328
rect 53470 16904 53526 16960
rect 53470 15680 53526 15736
rect 53194 15136 53250 15192
rect 52826 14456 52882 14512
rect 52458 14320 52514 14376
rect 52274 14048 52330 14104
rect 52090 10240 52146 10296
rect 52366 13776 52422 13832
rect 53746 16224 53802 16280
rect 53930 15952 53986 16008
rect 53102 14864 53158 14920
rect 52918 13796 52974 13832
rect 52918 13776 52920 13796
rect 52920 13776 52972 13796
rect 52972 13776 52974 13796
rect 52826 12980 52882 13016
rect 52826 12960 52828 12980
rect 52828 12960 52880 12980
rect 52880 12960 52882 12980
rect 53010 12960 53066 13016
rect 53010 12416 53066 12472
rect 52918 12144 52974 12200
rect 52274 11056 52330 11112
rect 52642 10512 52698 10568
rect 52550 10376 52606 10432
rect 50526 3476 50528 3496
rect 50528 3476 50580 3496
rect 50580 3476 50582 3496
rect 50526 3440 50582 3476
rect 50618 2760 50674 2816
rect 51446 4020 51448 4040
rect 51448 4020 51500 4040
rect 51500 4020 51502 4040
rect 51446 3984 51502 4020
rect 51814 3440 51870 3496
rect 52550 3984 52606 4040
rect 52918 3440 52974 3496
rect 52182 3304 52238 3360
rect 51998 3188 52054 3224
rect 51998 3168 52000 3188
rect 52000 3168 52052 3188
rect 52052 3168 52054 3188
rect 53286 12724 53288 12744
rect 53288 12724 53340 12744
rect 53340 12724 53342 12744
rect 53286 12688 53342 12724
rect 53378 12416 53434 12472
rect 53378 10784 53434 10840
rect 53746 12280 53802 12336
rect 53838 11464 53894 11520
rect 53838 11328 53894 11384
rect 53746 10920 53802 10976
rect 53654 10784 53710 10840
rect 53470 10512 53526 10568
rect 55826 27770 55882 27772
rect 55906 27770 55962 27772
rect 55986 27770 56042 27772
rect 56066 27770 56122 27772
rect 55826 27718 55872 27770
rect 55872 27718 55882 27770
rect 55906 27718 55936 27770
rect 55936 27718 55948 27770
rect 55948 27718 55962 27770
rect 55986 27718 56000 27770
rect 56000 27718 56012 27770
rect 56012 27718 56042 27770
rect 56066 27718 56076 27770
rect 56076 27718 56122 27770
rect 55826 27716 55882 27718
rect 55906 27716 55962 27718
rect 55986 27716 56042 27718
rect 56066 27716 56122 27718
rect 55310 17756 55312 17776
rect 55312 17756 55364 17776
rect 55364 17756 55366 17776
rect 55310 17720 55366 17756
rect 54482 17312 54538 17368
rect 54666 16904 54722 16960
rect 54298 14864 54354 14920
rect 54206 14728 54262 14784
rect 54114 12960 54170 13016
rect 54482 16360 54538 16416
rect 54390 14456 54446 14512
rect 55402 16768 55458 16824
rect 54942 15816 54998 15872
rect 54758 15680 54814 15736
rect 54390 11872 54446 11928
rect 55826 26682 55882 26684
rect 55906 26682 55962 26684
rect 55986 26682 56042 26684
rect 56066 26682 56122 26684
rect 55826 26630 55872 26682
rect 55872 26630 55882 26682
rect 55906 26630 55936 26682
rect 55936 26630 55948 26682
rect 55948 26630 55962 26682
rect 55986 26630 56000 26682
rect 56000 26630 56012 26682
rect 56012 26630 56042 26682
rect 56066 26630 56076 26682
rect 56076 26630 56122 26682
rect 55826 26628 55882 26630
rect 55906 26628 55962 26630
rect 55986 26628 56042 26630
rect 56066 26628 56122 26630
rect 55826 25594 55882 25596
rect 55906 25594 55962 25596
rect 55986 25594 56042 25596
rect 56066 25594 56122 25596
rect 55826 25542 55872 25594
rect 55872 25542 55882 25594
rect 55906 25542 55936 25594
rect 55936 25542 55948 25594
rect 55948 25542 55962 25594
rect 55986 25542 56000 25594
rect 56000 25542 56012 25594
rect 56012 25542 56042 25594
rect 56066 25542 56076 25594
rect 56076 25542 56122 25594
rect 55826 25540 55882 25542
rect 55906 25540 55962 25542
rect 55986 25540 56042 25542
rect 56066 25540 56122 25542
rect 55826 24506 55882 24508
rect 55906 24506 55962 24508
rect 55986 24506 56042 24508
rect 56066 24506 56122 24508
rect 55826 24454 55872 24506
rect 55872 24454 55882 24506
rect 55906 24454 55936 24506
rect 55936 24454 55948 24506
rect 55948 24454 55962 24506
rect 55986 24454 56000 24506
rect 56000 24454 56012 24506
rect 56012 24454 56042 24506
rect 56066 24454 56076 24506
rect 56076 24454 56122 24506
rect 55826 24452 55882 24454
rect 55906 24452 55962 24454
rect 55986 24452 56042 24454
rect 56066 24452 56122 24454
rect 55826 23418 55882 23420
rect 55906 23418 55962 23420
rect 55986 23418 56042 23420
rect 56066 23418 56122 23420
rect 55826 23366 55872 23418
rect 55872 23366 55882 23418
rect 55906 23366 55936 23418
rect 55936 23366 55948 23418
rect 55948 23366 55962 23418
rect 55986 23366 56000 23418
rect 56000 23366 56012 23418
rect 56012 23366 56042 23418
rect 56066 23366 56076 23418
rect 56076 23366 56122 23418
rect 55826 23364 55882 23366
rect 55906 23364 55962 23366
rect 55986 23364 56042 23366
rect 56066 23364 56122 23366
rect 55826 22330 55882 22332
rect 55906 22330 55962 22332
rect 55986 22330 56042 22332
rect 56066 22330 56122 22332
rect 55826 22278 55872 22330
rect 55872 22278 55882 22330
rect 55906 22278 55936 22330
rect 55936 22278 55948 22330
rect 55948 22278 55962 22330
rect 55986 22278 56000 22330
rect 56000 22278 56012 22330
rect 56012 22278 56042 22330
rect 56066 22278 56076 22330
rect 56076 22278 56122 22330
rect 55826 22276 55882 22278
rect 55906 22276 55962 22278
rect 55986 22276 56042 22278
rect 56066 22276 56122 22278
rect 55826 21242 55882 21244
rect 55906 21242 55962 21244
rect 55986 21242 56042 21244
rect 56066 21242 56122 21244
rect 55826 21190 55872 21242
rect 55872 21190 55882 21242
rect 55906 21190 55936 21242
rect 55936 21190 55948 21242
rect 55948 21190 55962 21242
rect 55986 21190 56000 21242
rect 56000 21190 56012 21242
rect 56012 21190 56042 21242
rect 56066 21190 56076 21242
rect 56076 21190 56122 21242
rect 55826 21188 55882 21190
rect 55906 21188 55962 21190
rect 55986 21188 56042 21190
rect 56066 21188 56122 21190
rect 55826 20154 55882 20156
rect 55906 20154 55962 20156
rect 55986 20154 56042 20156
rect 56066 20154 56122 20156
rect 55826 20102 55872 20154
rect 55872 20102 55882 20154
rect 55906 20102 55936 20154
rect 55936 20102 55948 20154
rect 55948 20102 55962 20154
rect 55986 20102 56000 20154
rect 56000 20102 56012 20154
rect 56012 20102 56042 20154
rect 56066 20102 56076 20154
rect 56076 20102 56122 20154
rect 55826 20100 55882 20102
rect 55906 20100 55962 20102
rect 55986 20100 56042 20102
rect 56066 20100 56122 20102
rect 55826 19066 55882 19068
rect 55906 19066 55962 19068
rect 55986 19066 56042 19068
rect 56066 19066 56122 19068
rect 55826 19014 55872 19066
rect 55872 19014 55882 19066
rect 55906 19014 55936 19066
rect 55936 19014 55948 19066
rect 55948 19014 55962 19066
rect 55986 19014 56000 19066
rect 56000 19014 56012 19066
rect 56012 19014 56042 19066
rect 56066 19014 56076 19066
rect 56076 19014 56122 19066
rect 55826 19012 55882 19014
rect 55906 19012 55962 19014
rect 55986 19012 56042 19014
rect 56066 19012 56122 19014
rect 55826 17978 55882 17980
rect 55906 17978 55962 17980
rect 55986 17978 56042 17980
rect 56066 17978 56122 17980
rect 55826 17926 55872 17978
rect 55872 17926 55882 17978
rect 55906 17926 55936 17978
rect 55936 17926 55948 17978
rect 55948 17926 55962 17978
rect 55986 17926 56000 17978
rect 56000 17926 56012 17978
rect 56012 17926 56042 17978
rect 56066 17926 56076 17978
rect 56076 17926 56122 17978
rect 55826 17924 55882 17926
rect 55906 17924 55962 17926
rect 55986 17924 56042 17926
rect 56066 17924 56122 17926
rect 55826 16890 55882 16892
rect 55906 16890 55962 16892
rect 55986 16890 56042 16892
rect 56066 16890 56122 16892
rect 55826 16838 55872 16890
rect 55872 16838 55882 16890
rect 55906 16838 55936 16890
rect 55936 16838 55948 16890
rect 55948 16838 55962 16890
rect 55986 16838 56000 16890
rect 56000 16838 56012 16890
rect 56012 16838 56042 16890
rect 56066 16838 56076 16890
rect 56076 16838 56122 16890
rect 55826 16836 55882 16838
rect 55906 16836 55962 16838
rect 55986 16836 56042 16838
rect 56066 16836 56122 16838
rect 55494 16088 55550 16144
rect 55678 15952 55734 16008
rect 55826 15802 55882 15804
rect 55906 15802 55962 15804
rect 55986 15802 56042 15804
rect 56066 15802 56122 15804
rect 55826 15750 55872 15802
rect 55872 15750 55882 15802
rect 55906 15750 55936 15802
rect 55936 15750 55948 15802
rect 55948 15750 55962 15802
rect 55986 15750 56000 15802
rect 56000 15750 56012 15802
rect 56012 15750 56042 15802
rect 56066 15750 56076 15802
rect 56076 15750 56122 15802
rect 55826 15748 55882 15750
rect 55906 15748 55962 15750
rect 55986 15748 56042 15750
rect 56066 15748 56122 15750
rect 56322 18284 56378 18320
rect 56322 18264 56324 18284
rect 56324 18264 56376 18284
rect 56376 18264 56378 18284
rect 56414 18128 56470 18184
rect 56874 17584 56930 17640
rect 56782 17196 56838 17232
rect 56782 17176 56784 17196
rect 56784 17176 56836 17196
rect 56836 17176 56838 17196
rect 56598 15952 56654 16008
rect 56322 15544 56378 15600
rect 54942 14184 54998 14240
rect 55126 14184 55182 14240
rect 54758 12960 54814 13016
rect 55826 14714 55882 14716
rect 55906 14714 55962 14716
rect 55986 14714 56042 14716
rect 56066 14714 56122 14716
rect 55826 14662 55872 14714
rect 55872 14662 55882 14714
rect 55906 14662 55936 14714
rect 55936 14662 55948 14714
rect 55948 14662 55962 14714
rect 55986 14662 56000 14714
rect 56000 14662 56012 14714
rect 56012 14662 56042 14714
rect 56066 14662 56076 14714
rect 56076 14662 56122 14714
rect 55826 14660 55882 14662
rect 55906 14660 55962 14662
rect 55986 14660 56042 14662
rect 56066 14660 56122 14662
rect 54666 11892 54722 11928
rect 54666 11872 54668 11892
rect 54668 11872 54720 11892
rect 54720 11872 54722 11892
rect 55678 13640 55734 13696
rect 55826 13626 55882 13628
rect 55906 13626 55962 13628
rect 55986 13626 56042 13628
rect 56066 13626 56122 13628
rect 55826 13574 55872 13626
rect 55872 13574 55882 13626
rect 55906 13574 55936 13626
rect 55936 13574 55948 13626
rect 55948 13574 55962 13626
rect 55986 13574 56000 13626
rect 56000 13574 56012 13626
rect 56012 13574 56042 13626
rect 56066 13574 56076 13626
rect 56076 13574 56122 13626
rect 55826 13572 55882 13574
rect 55906 13572 55962 13574
rect 55986 13572 56042 13574
rect 56066 13572 56122 13574
rect 55678 13096 55734 13152
rect 56046 12960 56102 13016
rect 55826 12538 55882 12540
rect 55906 12538 55962 12540
rect 55986 12538 56042 12540
rect 56066 12538 56122 12540
rect 55826 12486 55872 12538
rect 55872 12486 55882 12538
rect 55906 12486 55936 12538
rect 55936 12486 55948 12538
rect 55948 12486 55962 12538
rect 55986 12486 56000 12538
rect 56000 12486 56012 12538
rect 56012 12486 56042 12538
rect 56066 12486 56076 12538
rect 56076 12486 56122 12538
rect 55826 12484 55882 12486
rect 55906 12484 55962 12486
rect 55986 12484 56042 12486
rect 56066 12484 56122 12486
rect 55218 11464 55274 11520
rect 55826 11450 55882 11452
rect 55906 11450 55962 11452
rect 55986 11450 56042 11452
rect 56066 11450 56122 11452
rect 55826 11398 55872 11450
rect 55872 11398 55882 11450
rect 55906 11398 55936 11450
rect 55936 11398 55948 11450
rect 55948 11398 55962 11450
rect 55986 11398 56000 11450
rect 56000 11398 56012 11450
rect 56012 11398 56042 11450
rect 56066 11398 56076 11450
rect 56076 11398 56122 11450
rect 55826 11396 55882 11398
rect 55906 11396 55962 11398
rect 55986 11396 56042 11398
rect 56066 11396 56122 11398
rect 55218 11092 55220 11112
rect 55220 11092 55272 11112
rect 55272 11092 55274 11112
rect 55218 11056 55274 11092
rect 55402 10376 55458 10432
rect 55826 10362 55882 10364
rect 55906 10362 55962 10364
rect 55986 10362 56042 10364
rect 56066 10362 56122 10364
rect 55826 10310 55872 10362
rect 55872 10310 55882 10362
rect 55906 10310 55936 10362
rect 55936 10310 55948 10362
rect 55948 10310 55962 10362
rect 55986 10310 56000 10362
rect 56000 10310 56012 10362
rect 56012 10310 56042 10362
rect 56066 10310 56076 10362
rect 56076 10310 56122 10362
rect 55826 10308 55882 10310
rect 55906 10308 55962 10310
rect 55986 10308 56042 10310
rect 56066 10308 56122 10310
rect 56874 15136 56930 15192
rect 56966 14900 56968 14920
rect 56968 14900 57020 14920
rect 57020 14900 57022 14920
rect 56966 14864 57022 14900
rect 56874 14728 56930 14784
rect 57886 17448 57942 17504
rect 57426 16632 57482 16688
rect 57058 14048 57114 14104
rect 56874 13776 56930 13832
rect 57058 13504 57114 13560
rect 57518 16496 57574 16552
rect 57610 14456 57666 14512
rect 57242 14048 57298 14104
rect 56598 12552 56654 12608
rect 56414 11464 56470 11520
rect 55826 9274 55882 9276
rect 55906 9274 55962 9276
rect 55986 9274 56042 9276
rect 56066 9274 56122 9276
rect 55826 9222 55872 9274
rect 55872 9222 55882 9274
rect 55906 9222 55936 9274
rect 55936 9222 55948 9274
rect 55948 9222 55962 9274
rect 55986 9222 56000 9274
rect 56000 9222 56012 9274
rect 56012 9222 56042 9274
rect 56066 9222 56076 9274
rect 56076 9222 56122 9274
rect 55826 9220 55882 9222
rect 55906 9220 55962 9222
rect 55986 9220 56042 9222
rect 56066 9220 56122 9222
rect 55826 8186 55882 8188
rect 55906 8186 55962 8188
rect 55986 8186 56042 8188
rect 56066 8186 56122 8188
rect 55826 8134 55872 8186
rect 55872 8134 55882 8186
rect 55906 8134 55936 8186
rect 55936 8134 55948 8186
rect 55948 8134 55962 8186
rect 55986 8134 56000 8186
rect 56000 8134 56012 8186
rect 56012 8134 56042 8186
rect 56066 8134 56076 8186
rect 56076 8134 56122 8186
rect 55826 8132 55882 8134
rect 55906 8132 55962 8134
rect 55986 8132 56042 8134
rect 56066 8132 56122 8134
rect 55826 7098 55882 7100
rect 55906 7098 55962 7100
rect 55986 7098 56042 7100
rect 56066 7098 56122 7100
rect 55826 7046 55872 7098
rect 55872 7046 55882 7098
rect 55906 7046 55936 7098
rect 55936 7046 55948 7098
rect 55948 7046 55962 7098
rect 55986 7046 56000 7098
rect 56000 7046 56012 7098
rect 56012 7046 56042 7098
rect 56066 7046 56076 7098
rect 56076 7046 56122 7098
rect 55826 7044 55882 7046
rect 55906 7044 55962 7046
rect 55986 7044 56042 7046
rect 56066 7044 56122 7046
rect 55826 6010 55882 6012
rect 55906 6010 55962 6012
rect 55986 6010 56042 6012
rect 56066 6010 56122 6012
rect 55826 5958 55872 6010
rect 55872 5958 55882 6010
rect 55906 5958 55936 6010
rect 55936 5958 55948 6010
rect 55948 5958 55962 6010
rect 55986 5958 56000 6010
rect 56000 5958 56012 6010
rect 56012 5958 56042 6010
rect 56066 5958 56076 6010
rect 56076 5958 56122 6010
rect 55826 5956 55882 5958
rect 55906 5956 55962 5958
rect 55986 5956 56042 5958
rect 56066 5956 56122 5958
rect 55826 4922 55882 4924
rect 55906 4922 55962 4924
rect 55986 4922 56042 4924
rect 56066 4922 56122 4924
rect 55826 4870 55872 4922
rect 55872 4870 55882 4922
rect 55906 4870 55936 4922
rect 55936 4870 55948 4922
rect 55948 4870 55962 4922
rect 55986 4870 56000 4922
rect 56000 4870 56012 4922
rect 56012 4870 56042 4922
rect 56066 4870 56076 4922
rect 56076 4870 56122 4922
rect 55826 4868 55882 4870
rect 55906 4868 55962 4870
rect 55986 4868 56042 4870
rect 56066 4868 56122 4870
rect 55826 3834 55882 3836
rect 55906 3834 55962 3836
rect 55986 3834 56042 3836
rect 56066 3834 56122 3836
rect 55826 3782 55872 3834
rect 55872 3782 55882 3834
rect 55906 3782 55936 3834
rect 55936 3782 55948 3834
rect 55948 3782 55962 3834
rect 55986 3782 56000 3834
rect 56000 3782 56012 3834
rect 56012 3782 56042 3834
rect 56066 3782 56076 3834
rect 56076 3782 56122 3834
rect 55826 3780 55882 3782
rect 55906 3780 55962 3782
rect 55986 3780 56042 3782
rect 56066 3780 56122 3782
rect 56598 11500 56600 11520
rect 56600 11500 56652 11520
rect 56652 11500 56654 11520
rect 56598 11464 56654 11500
rect 57426 13640 57482 13696
rect 56966 10648 57022 10704
rect 57518 11464 57574 11520
rect 55826 2746 55882 2748
rect 55906 2746 55962 2748
rect 55986 2746 56042 2748
rect 56066 2746 56122 2748
rect 55826 2694 55872 2746
rect 55872 2694 55882 2746
rect 55906 2694 55936 2746
rect 55936 2694 55948 2746
rect 55948 2694 55962 2746
rect 55986 2694 56000 2746
rect 56000 2694 56012 2746
rect 56012 2694 56042 2746
rect 56066 2694 56076 2746
rect 56076 2694 56122 2746
rect 55826 2692 55882 2694
rect 55906 2692 55962 2694
rect 55986 2692 56042 2694
rect 56066 2692 56122 2694
rect 57610 10104 57666 10160
rect 59266 21392 59322 21448
rect 58622 17720 58678 17776
rect 58622 17176 58678 17232
rect 57978 16088 58034 16144
rect 58806 17040 58862 17096
rect 58254 16108 58310 16144
rect 58622 16224 58678 16280
rect 58254 16088 58256 16108
rect 58256 16088 58308 16108
rect 58308 16088 58310 16108
rect 57794 14340 57850 14376
rect 57794 14320 57796 14340
rect 57796 14320 57848 14340
rect 57848 14320 57850 14340
rect 57978 15988 57980 16008
rect 57980 15988 58032 16008
rect 58032 15988 58034 16008
rect 57978 15952 58034 15988
rect 57978 14592 58034 14648
rect 58070 13232 58126 13288
rect 58162 12960 58218 13016
rect 58070 11192 58126 11248
rect 58622 15564 58678 15600
rect 58622 15544 58624 15564
rect 58624 15544 58676 15564
rect 58676 15544 58678 15564
rect 58530 14456 58586 14512
rect 58346 13268 58348 13288
rect 58348 13268 58400 13288
rect 58400 13268 58402 13288
rect 58346 13232 58402 13268
rect 58346 12960 58402 13016
rect 58714 12416 58770 12472
rect 58346 11464 58402 11520
rect 58898 16768 58954 16824
rect 58898 16496 58954 16552
rect 59082 17484 59084 17504
rect 59084 17484 59136 17504
rect 59136 17484 59138 17504
rect 59082 17448 59138 17484
rect 58806 11192 58862 11248
rect 56506 2352 56562 2408
rect 60462 17756 60464 17776
rect 60464 17756 60516 17776
rect 60516 17756 60518 17776
rect 60462 17720 60518 17756
rect 60830 17740 60886 17776
rect 60830 17720 60832 17740
rect 60832 17720 60884 17740
rect 60884 17720 60886 17740
rect 60278 17312 60334 17368
rect 59266 15952 59322 16008
rect 59542 16632 59598 16688
rect 59450 13232 59506 13288
rect 59266 11872 59322 11928
rect 59358 10920 59414 10976
rect 59910 15136 59966 15192
rect 60002 14728 60058 14784
rect 60002 13776 60058 13832
rect 60646 17040 60702 17096
rect 59910 12280 59966 12336
rect 60738 16360 60794 16416
rect 60554 15308 60556 15328
rect 60556 15308 60608 15328
rect 60608 15308 60610 15328
rect 60554 15272 60610 15308
rect 60830 14900 60832 14920
rect 60832 14900 60884 14920
rect 60884 14900 60886 14920
rect 60830 14864 60886 14900
rect 61842 15428 61898 15464
rect 61842 15408 61844 15428
rect 61844 15408 61896 15428
rect 61896 15408 61898 15428
rect 62210 15544 62266 15600
rect 62118 14476 62174 14512
rect 62118 14456 62120 14476
rect 62120 14456 62172 14476
rect 62172 14456 62174 14476
rect 60278 14184 60334 14240
rect 60278 13504 60334 13560
rect 60554 14184 60610 14240
rect 60646 13812 60648 13832
rect 60648 13812 60700 13832
rect 60700 13812 60702 13832
rect 60646 13776 60702 13812
rect 60830 13776 60886 13832
rect 61014 13812 61016 13832
rect 61016 13812 61068 13832
rect 61068 13812 61070 13832
rect 61014 13776 61070 13812
rect 60554 13504 60610 13560
rect 60554 13268 60556 13288
rect 60556 13268 60608 13288
rect 60608 13268 60610 13288
rect 60554 13232 60610 13268
rect 60738 13232 60794 13288
rect 60370 12416 60426 12472
rect 60278 12280 60334 12336
rect 60830 13096 60886 13152
rect 60462 12008 60518 12064
rect 60646 12044 60648 12064
rect 60648 12044 60700 12064
rect 60700 12044 60702 12064
rect 60646 12008 60702 12044
rect 60278 11464 60334 11520
rect 60554 11464 60610 11520
rect 60646 10920 60702 10976
rect 61106 12280 61162 12336
rect 61106 11736 61162 11792
rect 59634 10512 59690 10568
rect 61566 14068 61622 14104
rect 61566 14048 61568 14068
rect 61568 14048 61620 14068
rect 61620 14048 61622 14068
rect 61382 13640 61438 13696
rect 61842 14048 61898 14104
rect 61842 10376 61898 10432
rect 62118 13676 62120 13696
rect 62120 13676 62172 13696
rect 62172 13676 62174 13696
rect 62118 13640 62174 13676
rect 62302 15136 62358 15192
rect 62394 15020 62450 15056
rect 62394 15000 62396 15020
rect 62396 15000 62448 15020
rect 62448 15000 62450 15020
rect 62578 17484 62580 17504
rect 62580 17484 62632 17504
rect 62632 17484 62634 17504
rect 62578 17448 62634 17484
rect 63038 16668 63040 16688
rect 63040 16668 63092 16688
rect 63092 16668 63094 16688
rect 63038 16632 63094 16668
rect 62670 15564 62726 15600
rect 62670 15544 62672 15564
rect 62672 15544 62724 15564
rect 62724 15544 62726 15564
rect 62578 15000 62634 15056
rect 62302 13504 62358 13560
rect 62486 12280 62542 12336
rect 62302 12008 62358 12064
rect 62762 12552 62818 12608
rect 62670 12416 62726 12472
rect 62670 11736 62726 11792
rect 63314 16768 63370 16824
rect 63130 15272 63186 15328
rect 62946 14864 63002 14920
rect 63038 14048 63094 14104
rect 63038 12552 63094 12608
rect 63038 11872 63094 11928
rect 62946 11464 63002 11520
rect 62854 10920 62910 10976
rect 63038 10648 63094 10704
rect 63314 15544 63370 15600
rect 63222 14456 63278 14512
rect 63222 12960 63278 13016
rect 63314 12144 63370 12200
rect 63590 15020 63646 15056
rect 63590 15000 63592 15020
rect 63592 15000 63644 15020
rect 63644 15000 63646 15020
rect 63498 13776 63554 13832
rect 63590 12552 63646 12608
rect 63406 11756 63462 11792
rect 63406 11736 63408 11756
rect 63408 11736 63460 11756
rect 63460 11736 63462 11756
rect 63774 15272 63830 15328
rect 64510 17584 64566 17640
rect 64694 16904 64750 16960
rect 64050 14356 64052 14376
rect 64052 14356 64104 14376
rect 64104 14356 64106 14376
rect 64050 14320 64106 14356
rect 64050 14048 64106 14104
rect 63774 12552 63830 12608
rect 63682 12416 63738 12472
rect 63590 12144 63646 12200
rect 63590 11636 63592 11656
rect 63592 11636 63644 11656
rect 63644 11636 63646 11656
rect 63590 11600 63646 11636
rect 63590 11464 63646 11520
rect 63406 10784 63462 10840
rect 63406 10668 63462 10704
rect 63406 10648 63408 10668
rect 63408 10648 63460 10668
rect 63460 10648 63462 10668
rect 63498 10240 63554 10296
rect 63774 11872 63830 11928
rect 63774 10512 63830 10568
rect 64050 13096 64106 13152
rect 64050 11756 64106 11792
rect 64050 11736 64052 11756
rect 64052 11736 64104 11756
rect 64104 11736 64106 11756
rect 64418 14184 64474 14240
rect 64694 15136 64750 15192
rect 64970 15136 65026 15192
rect 64510 13232 64566 13288
rect 64326 11192 64382 11248
rect 64510 11092 64512 11112
rect 64512 11092 64564 11112
rect 64564 11092 64566 11112
rect 64510 11056 64566 11092
rect 64878 12280 64934 12336
rect 64878 11056 64934 11112
rect 66800 27226 66856 27228
rect 66880 27226 66936 27228
rect 66960 27226 67016 27228
rect 67040 27226 67096 27228
rect 66800 27174 66846 27226
rect 66846 27174 66856 27226
rect 66880 27174 66910 27226
rect 66910 27174 66922 27226
rect 66922 27174 66936 27226
rect 66960 27174 66974 27226
rect 66974 27174 66986 27226
rect 66986 27174 67016 27226
rect 67040 27174 67050 27226
rect 67050 27174 67096 27226
rect 66800 27172 66856 27174
rect 66880 27172 66936 27174
rect 66960 27172 67016 27174
rect 67040 27172 67096 27174
rect 66800 26138 66856 26140
rect 66880 26138 66936 26140
rect 66960 26138 67016 26140
rect 67040 26138 67096 26140
rect 66800 26086 66846 26138
rect 66846 26086 66856 26138
rect 66880 26086 66910 26138
rect 66910 26086 66922 26138
rect 66922 26086 66936 26138
rect 66960 26086 66974 26138
rect 66974 26086 66986 26138
rect 66986 26086 67016 26138
rect 67040 26086 67050 26138
rect 67050 26086 67096 26138
rect 66800 26084 66856 26086
rect 66880 26084 66936 26086
rect 66960 26084 67016 26086
rect 67040 26084 67096 26086
rect 66800 25050 66856 25052
rect 66880 25050 66936 25052
rect 66960 25050 67016 25052
rect 67040 25050 67096 25052
rect 66800 24998 66846 25050
rect 66846 24998 66856 25050
rect 66880 24998 66910 25050
rect 66910 24998 66922 25050
rect 66922 24998 66936 25050
rect 66960 24998 66974 25050
rect 66974 24998 66986 25050
rect 66986 24998 67016 25050
rect 67040 24998 67050 25050
rect 67050 24998 67096 25050
rect 66800 24996 66856 24998
rect 66880 24996 66936 24998
rect 66960 24996 67016 24998
rect 67040 24996 67096 24998
rect 66800 23962 66856 23964
rect 66880 23962 66936 23964
rect 66960 23962 67016 23964
rect 67040 23962 67096 23964
rect 66800 23910 66846 23962
rect 66846 23910 66856 23962
rect 66880 23910 66910 23962
rect 66910 23910 66922 23962
rect 66922 23910 66936 23962
rect 66960 23910 66974 23962
rect 66974 23910 66986 23962
rect 66986 23910 67016 23962
rect 67040 23910 67050 23962
rect 67050 23910 67096 23962
rect 66800 23908 66856 23910
rect 66880 23908 66936 23910
rect 66960 23908 67016 23910
rect 67040 23908 67096 23910
rect 66800 22874 66856 22876
rect 66880 22874 66936 22876
rect 66960 22874 67016 22876
rect 67040 22874 67096 22876
rect 66800 22822 66846 22874
rect 66846 22822 66856 22874
rect 66880 22822 66910 22874
rect 66910 22822 66922 22874
rect 66922 22822 66936 22874
rect 66960 22822 66974 22874
rect 66974 22822 66986 22874
rect 66986 22822 67016 22874
rect 67040 22822 67050 22874
rect 67050 22822 67096 22874
rect 66800 22820 66856 22822
rect 66880 22820 66936 22822
rect 66960 22820 67016 22822
rect 67040 22820 67096 22822
rect 66800 21786 66856 21788
rect 66880 21786 66936 21788
rect 66960 21786 67016 21788
rect 67040 21786 67096 21788
rect 66800 21734 66846 21786
rect 66846 21734 66856 21786
rect 66880 21734 66910 21786
rect 66910 21734 66922 21786
rect 66922 21734 66936 21786
rect 66960 21734 66974 21786
rect 66974 21734 66986 21786
rect 66986 21734 67016 21786
rect 67040 21734 67050 21786
rect 67050 21734 67096 21786
rect 66800 21732 66856 21734
rect 66880 21732 66936 21734
rect 66960 21732 67016 21734
rect 67040 21732 67096 21734
rect 66800 20698 66856 20700
rect 66880 20698 66936 20700
rect 66960 20698 67016 20700
rect 67040 20698 67096 20700
rect 66800 20646 66846 20698
rect 66846 20646 66856 20698
rect 66880 20646 66910 20698
rect 66910 20646 66922 20698
rect 66922 20646 66936 20698
rect 66960 20646 66974 20698
rect 66974 20646 66986 20698
rect 66986 20646 67016 20698
rect 67040 20646 67050 20698
rect 67050 20646 67096 20698
rect 66800 20644 66856 20646
rect 66880 20644 66936 20646
rect 66960 20644 67016 20646
rect 67040 20644 67096 20646
rect 66800 19610 66856 19612
rect 66880 19610 66936 19612
rect 66960 19610 67016 19612
rect 67040 19610 67096 19612
rect 66800 19558 66846 19610
rect 66846 19558 66856 19610
rect 66880 19558 66910 19610
rect 66910 19558 66922 19610
rect 66922 19558 66936 19610
rect 66960 19558 66974 19610
rect 66974 19558 66986 19610
rect 66986 19558 67016 19610
rect 67040 19558 67050 19610
rect 67050 19558 67096 19610
rect 66800 19556 66856 19558
rect 66880 19556 66936 19558
rect 66960 19556 67016 19558
rect 67040 19556 67096 19558
rect 66800 18522 66856 18524
rect 66880 18522 66936 18524
rect 66960 18522 67016 18524
rect 67040 18522 67096 18524
rect 66800 18470 66846 18522
rect 66846 18470 66856 18522
rect 66880 18470 66910 18522
rect 66910 18470 66922 18522
rect 66922 18470 66936 18522
rect 66960 18470 66974 18522
rect 66974 18470 66986 18522
rect 66986 18470 67016 18522
rect 67040 18470 67050 18522
rect 67050 18470 67096 18522
rect 66800 18468 66856 18470
rect 66880 18468 66936 18470
rect 66960 18468 67016 18470
rect 67040 18468 67096 18470
rect 66534 17312 66590 17368
rect 66800 17434 66856 17436
rect 66880 17434 66936 17436
rect 66960 17434 67016 17436
rect 67040 17434 67096 17436
rect 66800 17382 66846 17434
rect 66846 17382 66856 17434
rect 66880 17382 66910 17434
rect 66910 17382 66922 17434
rect 66922 17382 66936 17434
rect 66960 17382 66974 17434
rect 66974 17382 66986 17434
rect 66986 17382 67016 17434
rect 67040 17382 67050 17434
rect 67050 17382 67096 17434
rect 66800 17380 66856 17382
rect 66880 17380 66936 17382
rect 66960 17380 67016 17382
rect 67040 17380 67096 17382
rect 66994 17196 67050 17232
rect 66994 17176 66996 17196
rect 66996 17176 67048 17196
rect 67048 17176 67050 17196
rect 66442 17076 66444 17096
rect 66444 17076 66496 17096
rect 66496 17076 66498 17096
rect 66442 17040 66498 17076
rect 66258 16904 66314 16960
rect 66442 16496 66498 16552
rect 66800 16346 66856 16348
rect 66880 16346 66936 16348
rect 66960 16346 67016 16348
rect 67040 16346 67096 16348
rect 66800 16294 66846 16346
rect 66846 16294 66856 16346
rect 66880 16294 66910 16346
rect 66910 16294 66922 16346
rect 66922 16294 66936 16346
rect 66960 16294 66974 16346
rect 66974 16294 66986 16346
rect 66986 16294 67016 16346
rect 67040 16294 67050 16346
rect 67050 16294 67096 16346
rect 66800 16292 66856 16294
rect 66880 16292 66936 16294
rect 66960 16292 67016 16294
rect 67040 16292 67096 16294
rect 66074 16088 66130 16144
rect 65706 15020 65762 15056
rect 65706 15000 65708 15020
rect 65708 15000 65760 15020
rect 65760 15000 65762 15020
rect 66800 15258 66856 15260
rect 66880 15258 66936 15260
rect 66960 15258 67016 15260
rect 67040 15258 67096 15260
rect 66800 15206 66846 15258
rect 66846 15206 66856 15258
rect 66880 15206 66910 15258
rect 66910 15206 66922 15258
rect 66922 15206 66936 15258
rect 66960 15206 66974 15258
rect 66974 15206 66986 15258
rect 66986 15206 67016 15258
rect 67040 15206 67050 15258
rect 67050 15206 67096 15258
rect 66800 15204 66856 15206
rect 66880 15204 66936 15206
rect 66960 15204 67016 15206
rect 67040 15204 67096 15206
rect 65246 14864 65302 14920
rect 66718 14728 66774 14784
rect 65798 14048 65854 14104
rect 65154 13640 65210 13696
rect 66350 13504 66406 13560
rect 65982 12280 66038 12336
rect 66166 12008 66222 12064
rect 66800 14170 66856 14172
rect 66880 14170 66936 14172
rect 66960 14170 67016 14172
rect 67040 14170 67096 14172
rect 66800 14118 66846 14170
rect 66846 14118 66856 14170
rect 66880 14118 66910 14170
rect 66910 14118 66922 14170
rect 66922 14118 66936 14170
rect 66960 14118 66974 14170
rect 66974 14118 66986 14170
rect 66986 14118 67016 14170
rect 67040 14118 67050 14170
rect 67050 14118 67096 14170
rect 66800 14116 66856 14118
rect 66880 14116 66936 14118
rect 66960 14116 67016 14118
rect 67040 14116 67096 14118
rect 66800 13082 66856 13084
rect 66880 13082 66936 13084
rect 66960 13082 67016 13084
rect 67040 13082 67096 13084
rect 66800 13030 66846 13082
rect 66846 13030 66856 13082
rect 66880 13030 66910 13082
rect 66910 13030 66922 13082
rect 66922 13030 66936 13082
rect 66960 13030 66974 13082
rect 66974 13030 66986 13082
rect 66986 13030 67016 13082
rect 67040 13030 67050 13082
rect 67050 13030 67096 13082
rect 66800 13028 66856 13030
rect 66880 13028 66936 13030
rect 66960 13028 67016 13030
rect 67040 13028 67096 13030
rect 66626 12960 66682 13016
rect 67454 14320 67510 14376
rect 67822 14320 67878 14376
rect 67454 14184 67510 14240
rect 67730 14068 67786 14104
rect 67730 14048 67732 14068
rect 67732 14048 67784 14068
rect 67784 14048 67786 14068
rect 67454 13776 67510 13832
rect 67730 13096 67786 13152
rect 66800 11994 66856 11996
rect 66880 11994 66936 11996
rect 66960 11994 67016 11996
rect 67040 11994 67096 11996
rect 66800 11942 66846 11994
rect 66846 11942 66856 11994
rect 66880 11942 66910 11994
rect 66910 11942 66922 11994
rect 66922 11942 66936 11994
rect 66960 11942 66974 11994
rect 66974 11942 66986 11994
rect 66986 11942 67016 11994
rect 67040 11942 67050 11994
rect 67050 11942 67096 11994
rect 66800 11940 66856 11942
rect 66880 11940 66936 11942
rect 66960 11940 67016 11942
rect 67040 11940 67096 11942
rect 66994 11772 66996 11792
rect 66996 11772 67048 11792
rect 67048 11772 67050 11792
rect 66994 11736 67050 11772
rect 66810 11600 66866 11656
rect 67638 12416 67694 12472
rect 66534 11192 66590 11248
rect 66800 10906 66856 10908
rect 66880 10906 66936 10908
rect 66960 10906 67016 10908
rect 67040 10906 67096 10908
rect 66800 10854 66846 10906
rect 66846 10854 66856 10906
rect 66880 10854 66910 10906
rect 66910 10854 66922 10906
rect 66922 10854 66936 10906
rect 66960 10854 66974 10906
rect 66974 10854 66986 10906
rect 66986 10854 67016 10906
rect 67040 10854 67050 10906
rect 67050 10854 67096 10906
rect 66800 10852 66856 10854
rect 66880 10852 66936 10854
rect 66960 10852 67016 10854
rect 67040 10852 67096 10854
rect 66800 9818 66856 9820
rect 66880 9818 66936 9820
rect 66960 9818 67016 9820
rect 67040 9818 67096 9820
rect 66800 9766 66846 9818
rect 66846 9766 66856 9818
rect 66880 9766 66910 9818
rect 66910 9766 66922 9818
rect 66922 9766 66936 9818
rect 66960 9766 66974 9818
rect 66974 9766 66986 9818
rect 66986 9766 67016 9818
rect 67040 9766 67050 9818
rect 67050 9766 67096 9818
rect 66800 9764 66856 9766
rect 66880 9764 66936 9766
rect 66960 9764 67016 9766
rect 67040 9764 67096 9766
rect 67822 11328 67878 11384
rect 67546 11228 67548 11248
rect 67548 11228 67600 11248
rect 67600 11228 67602 11248
rect 67546 11192 67602 11228
rect 67730 11192 67786 11248
rect 67454 10376 67510 10432
rect 68926 25744 68982 25800
rect 68650 15136 68706 15192
rect 68650 14456 68706 14512
rect 69110 17584 69166 17640
rect 69294 17040 69350 17096
rect 69570 16904 69626 16960
rect 68926 14048 68982 14104
rect 69202 14340 69258 14376
rect 69202 14320 69204 14340
rect 69204 14320 69256 14340
rect 69256 14320 69258 14340
rect 69110 14184 69166 14240
rect 69938 14592 69994 14648
rect 70858 15156 70914 15192
rect 70858 15136 70860 15156
rect 70860 15136 70912 15156
rect 70912 15136 70914 15156
rect 70398 14492 70400 14512
rect 70400 14492 70452 14512
rect 70452 14492 70454 14512
rect 70398 14456 70454 14492
rect 69386 13524 69442 13560
rect 69386 13504 69388 13524
rect 69388 13504 69440 13524
rect 69440 13504 69442 13524
rect 69294 12960 69350 13016
rect 69478 13096 69534 13152
rect 68834 12552 68890 12608
rect 69846 13096 69902 13152
rect 69754 12144 69810 12200
rect 70306 13504 70362 13560
rect 70766 13096 70822 13152
rect 70214 12280 70270 12336
rect 69018 11600 69074 11656
rect 68742 11464 68798 11520
rect 69202 11328 69258 11384
rect 69386 11228 69388 11248
rect 69388 11228 69440 11248
rect 69440 11228 69442 11248
rect 69386 11192 69442 11228
rect 69294 11056 69350 11112
rect 66800 8730 66856 8732
rect 66880 8730 66936 8732
rect 66960 8730 67016 8732
rect 67040 8730 67096 8732
rect 66800 8678 66846 8730
rect 66846 8678 66856 8730
rect 66880 8678 66910 8730
rect 66910 8678 66922 8730
rect 66922 8678 66936 8730
rect 66960 8678 66974 8730
rect 66974 8678 66986 8730
rect 66986 8678 67016 8730
rect 67040 8678 67050 8730
rect 67050 8678 67096 8730
rect 66800 8676 66856 8678
rect 66880 8676 66936 8678
rect 66960 8676 67016 8678
rect 67040 8676 67096 8678
rect 66800 7642 66856 7644
rect 66880 7642 66936 7644
rect 66960 7642 67016 7644
rect 67040 7642 67096 7644
rect 66800 7590 66846 7642
rect 66846 7590 66856 7642
rect 66880 7590 66910 7642
rect 66910 7590 66922 7642
rect 66922 7590 66936 7642
rect 66960 7590 66974 7642
rect 66974 7590 66986 7642
rect 66986 7590 67016 7642
rect 67040 7590 67050 7642
rect 67050 7590 67096 7642
rect 66800 7588 66856 7590
rect 66880 7588 66936 7590
rect 66960 7588 67016 7590
rect 67040 7588 67096 7590
rect 66800 6554 66856 6556
rect 66880 6554 66936 6556
rect 66960 6554 67016 6556
rect 67040 6554 67096 6556
rect 66800 6502 66846 6554
rect 66846 6502 66856 6554
rect 66880 6502 66910 6554
rect 66910 6502 66922 6554
rect 66922 6502 66936 6554
rect 66960 6502 66974 6554
rect 66974 6502 66986 6554
rect 66986 6502 67016 6554
rect 67040 6502 67050 6554
rect 67050 6502 67096 6554
rect 66800 6500 66856 6502
rect 66880 6500 66936 6502
rect 66960 6500 67016 6502
rect 67040 6500 67096 6502
rect 66800 5466 66856 5468
rect 66880 5466 66936 5468
rect 66960 5466 67016 5468
rect 67040 5466 67096 5468
rect 66800 5414 66846 5466
rect 66846 5414 66856 5466
rect 66880 5414 66910 5466
rect 66910 5414 66922 5466
rect 66922 5414 66936 5466
rect 66960 5414 66974 5466
rect 66974 5414 66986 5466
rect 66986 5414 67016 5466
rect 67040 5414 67050 5466
rect 67050 5414 67096 5466
rect 66800 5412 66856 5414
rect 66880 5412 66936 5414
rect 66960 5412 67016 5414
rect 67040 5412 67096 5414
rect 66800 4378 66856 4380
rect 66880 4378 66936 4380
rect 66960 4378 67016 4380
rect 67040 4378 67096 4380
rect 66800 4326 66846 4378
rect 66846 4326 66856 4378
rect 66880 4326 66910 4378
rect 66910 4326 66922 4378
rect 66922 4326 66936 4378
rect 66960 4326 66974 4378
rect 66974 4326 66986 4378
rect 66986 4326 67016 4378
rect 67040 4326 67050 4378
rect 67050 4326 67096 4378
rect 66800 4324 66856 4326
rect 66880 4324 66936 4326
rect 66960 4324 67016 4326
rect 67040 4324 67096 4326
rect 66800 3290 66856 3292
rect 66880 3290 66936 3292
rect 66960 3290 67016 3292
rect 67040 3290 67096 3292
rect 66800 3238 66846 3290
rect 66846 3238 66856 3290
rect 66880 3238 66910 3290
rect 66910 3238 66922 3290
rect 66922 3238 66936 3290
rect 66960 3238 66974 3290
rect 66974 3238 66986 3290
rect 66986 3238 67016 3290
rect 67040 3238 67050 3290
rect 67050 3238 67096 3290
rect 66800 3236 66856 3238
rect 66880 3236 66936 3238
rect 66960 3236 67016 3238
rect 67040 3236 67096 3238
rect 70858 11772 70860 11792
rect 70860 11772 70912 11792
rect 70912 11772 70914 11792
rect 70858 11736 70914 11772
rect 71686 12960 71742 13016
rect 72422 12588 72424 12608
rect 72424 12588 72476 12608
rect 72476 12588 72478 12608
rect 72422 12552 72478 12588
rect 77774 27770 77830 27772
rect 77854 27770 77910 27772
rect 77934 27770 77990 27772
rect 78014 27770 78070 27772
rect 77774 27718 77820 27770
rect 77820 27718 77830 27770
rect 77854 27718 77884 27770
rect 77884 27718 77896 27770
rect 77896 27718 77910 27770
rect 77934 27718 77948 27770
rect 77948 27718 77960 27770
rect 77960 27718 77990 27770
rect 78014 27718 78024 27770
rect 78024 27718 78070 27770
rect 77774 27716 77830 27718
rect 77854 27716 77910 27718
rect 77934 27716 77990 27718
rect 78014 27716 78070 27718
rect 77774 26682 77830 26684
rect 77854 26682 77910 26684
rect 77934 26682 77990 26684
rect 78014 26682 78070 26684
rect 77774 26630 77820 26682
rect 77820 26630 77830 26682
rect 77854 26630 77884 26682
rect 77884 26630 77896 26682
rect 77896 26630 77910 26682
rect 77934 26630 77948 26682
rect 77948 26630 77960 26682
rect 77960 26630 77990 26682
rect 78014 26630 78024 26682
rect 78024 26630 78070 26682
rect 77774 26628 77830 26630
rect 77854 26628 77910 26630
rect 77934 26628 77990 26630
rect 78014 26628 78070 26630
rect 77774 25594 77830 25596
rect 77854 25594 77910 25596
rect 77934 25594 77990 25596
rect 78014 25594 78070 25596
rect 77774 25542 77820 25594
rect 77820 25542 77830 25594
rect 77854 25542 77884 25594
rect 77884 25542 77896 25594
rect 77896 25542 77910 25594
rect 77934 25542 77948 25594
rect 77948 25542 77960 25594
rect 77960 25542 77990 25594
rect 78014 25542 78024 25594
rect 78024 25542 78070 25594
rect 77774 25540 77830 25542
rect 77854 25540 77910 25542
rect 77934 25540 77990 25542
rect 78014 25540 78070 25542
rect 77774 24506 77830 24508
rect 77854 24506 77910 24508
rect 77934 24506 77990 24508
rect 78014 24506 78070 24508
rect 77774 24454 77820 24506
rect 77820 24454 77830 24506
rect 77854 24454 77884 24506
rect 77884 24454 77896 24506
rect 77896 24454 77910 24506
rect 77934 24454 77948 24506
rect 77948 24454 77960 24506
rect 77960 24454 77990 24506
rect 78014 24454 78024 24506
rect 78024 24454 78070 24506
rect 77774 24452 77830 24454
rect 77854 24452 77910 24454
rect 77934 24452 77990 24454
rect 78014 24452 78070 24454
rect 77774 23418 77830 23420
rect 77854 23418 77910 23420
rect 77934 23418 77990 23420
rect 78014 23418 78070 23420
rect 77774 23366 77820 23418
rect 77820 23366 77830 23418
rect 77854 23366 77884 23418
rect 77884 23366 77896 23418
rect 77896 23366 77910 23418
rect 77934 23366 77948 23418
rect 77948 23366 77960 23418
rect 77960 23366 77990 23418
rect 78014 23366 78024 23418
rect 78024 23366 78070 23418
rect 77774 23364 77830 23366
rect 77854 23364 77910 23366
rect 77934 23364 77990 23366
rect 78014 23364 78070 23366
rect 77774 22330 77830 22332
rect 77854 22330 77910 22332
rect 77934 22330 77990 22332
rect 78014 22330 78070 22332
rect 77774 22278 77820 22330
rect 77820 22278 77830 22330
rect 77854 22278 77884 22330
rect 77884 22278 77896 22330
rect 77896 22278 77910 22330
rect 77934 22278 77948 22330
rect 77948 22278 77960 22330
rect 77960 22278 77990 22330
rect 78014 22278 78024 22330
rect 78024 22278 78070 22330
rect 77774 22276 77830 22278
rect 77854 22276 77910 22278
rect 77934 22276 77990 22278
rect 78014 22276 78070 22278
rect 77774 21242 77830 21244
rect 77854 21242 77910 21244
rect 77934 21242 77990 21244
rect 78014 21242 78070 21244
rect 77774 21190 77820 21242
rect 77820 21190 77830 21242
rect 77854 21190 77884 21242
rect 77884 21190 77896 21242
rect 77896 21190 77910 21242
rect 77934 21190 77948 21242
rect 77948 21190 77960 21242
rect 77960 21190 77990 21242
rect 78014 21190 78024 21242
rect 78024 21190 78070 21242
rect 77774 21188 77830 21190
rect 77854 21188 77910 21190
rect 77934 21188 77990 21190
rect 78014 21188 78070 21190
rect 77774 20154 77830 20156
rect 77854 20154 77910 20156
rect 77934 20154 77990 20156
rect 78014 20154 78070 20156
rect 77774 20102 77820 20154
rect 77820 20102 77830 20154
rect 77854 20102 77884 20154
rect 77884 20102 77896 20154
rect 77896 20102 77910 20154
rect 77934 20102 77948 20154
rect 77948 20102 77960 20154
rect 77960 20102 77990 20154
rect 78014 20102 78024 20154
rect 78024 20102 78070 20154
rect 77774 20100 77830 20102
rect 77854 20100 77910 20102
rect 77934 20100 77990 20102
rect 78014 20100 78070 20102
rect 77774 19066 77830 19068
rect 77854 19066 77910 19068
rect 77934 19066 77990 19068
rect 78014 19066 78070 19068
rect 77774 19014 77820 19066
rect 77820 19014 77830 19066
rect 77854 19014 77884 19066
rect 77884 19014 77896 19066
rect 77896 19014 77910 19066
rect 77934 19014 77948 19066
rect 77948 19014 77960 19066
rect 77960 19014 77990 19066
rect 78014 19014 78024 19066
rect 78024 19014 78070 19066
rect 77774 19012 77830 19014
rect 77854 19012 77910 19014
rect 77934 19012 77990 19014
rect 78014 19012 78070 19014
rect 77774 17978 77830 17980
rect 77854 17978 77910 17980
rect 77934 17978 77990 17980
rect 78014 17978 78070 17980
rect 77774 17926 77820 17978
rect 77820 17926 77830 17978
rect 77854 17926 77884 17978
rect 77884 17926 77896 17978
rect 77896 17926 77910 17978
rect 77934 17926 77948 17978
rect 77948 17926 77960 17978
rect 77960 17926 77990 17978
rect 78014 17926 78024 17978
rect 78024 17926 78070 17978
rect 77774 17924 77830 17926
rect 77854 17924 77910 17926
rect 77934 17924 77990 17926
rect 78014 17924 78070 17926
rect 77774 16890 77830 16892
rect 77854 16890 77910 16892
rect 77934 16890 77990 16892
rect 78014 16890 78070 16892
rect 77774 16838 77820 16890
rect 77820 16838 77830 16890
rect 77854 16838 77884 16890
rect 77884 16838 77896 16890
rect 77896 16838 77910 16890
rect 77934 16838 77948 16890
rect 77948 16838 77960 16890
rect 77960 16838 77990 16890
rect 78014 16838 78024 16890
rect 78024 16838 78070 16890
rect 77774 16836 77830 16838
rect 77854 16836 77910 16838
rect 77934 16836 77990 16838
rect 78014 16836 78070 16838
rect 66800 2202 66856 2204
rect 66880 2202 66936 2204
rect 66960 2202 67016 2204
rect 67040 2202 67096 2204
rect 66800 2150 66846 2202
rect 66846 2150 66856 2202
rect 66880 2150 66910 2202
rect 66910 2150 66922 2202
rect 66922 2150 66936 2202
rect 66960 2150 66974 2202
rect 66974 2150 66986 2202
rect 66986 2150 67016 2202
rect 67040 2150 67050 2202
rect 67050 2150 67096 2202
rect 66800 2148 66856 2150
rect 66880 2148 66936 2150
rect 66960 2148 67016 2150
rect 67040 2148 67096 2150
rect 77774 15802 77830 15804
rect 77854 15802 77910 15804
rect 77934 15802 77990 15804
rect 78014 15802 78070 15804
rect 77774 15750 77820 15802
rect 77820 15750 77830 15802
rect 77854 15750 77884 15802
rect 77884 15750 77896 15802
rect 77896 15750 77910 15802
rect 77934 15750 77948 15802
rect 77948 15750 77960 15802
rect 77960 15750 77990 15802
rect 78014 15750 78024 15802
rect 78024 15750 78070 15802
rect 77774 15748 77830 15750
rect 77854 15748 77910 15750
rect 77934 15748 77990 15750
rect 78014 15748 78070 15750
rect 77774 14714 77830 14716
rect 77854 14714 77910 14716
rect 77934 14714 77990 14716
rect 78014 14714 78070 14716
rect 77774 14662 77820 14714
rect 77820 14662 77830 14714
rect 77854 14662 77884 14714
rect 77884 14662 77896 14714
rect 77896 14662 77910 14714
rect 77934 14662 77948 14714
rect 77948 14662 77960 14714
rect 77960 14662 77990 14714
rect 78014 14662 78024 14714
rect 78024 14662 78070 14714
rect 77774 14660 77830 14662
rect 77854 14660 77910 14662
rect 77934 14660 77990 14662
rect 78014 14660 78070 14662
rect 77774 13626 77830 13628
rect 77854 13626 77910 13628
rect 77934 13626 77990 13628
rect 78014 13626 78070 13628
rect 77774 13574 77820 13626
rect 77820 13574 77830 13626
rect 77854 13574 77884 13626
rect 77884 13574 77896 13626
rect 77896 13574 77910 13626
rect 77934 13574 77948 13626
rect 77948 13574 77960 13626
rect 77960 13574 77990 13626
rect 78014 13574 78024 13626
rect 78024 13574 78070 13626
rect 77774 13572 77830 13574
rect 77854 13572 77910 13574
rect 77934 13572 77990 13574
rect 78014 13572 78070 13574
rect 80242 24112 80298 24168
rect 79598 13368 79654 13424
rect 77774 12538 77830 12540
rect 77854 12538 77910 12540
rect 77934 12538 77990 12540
rect 78014 12538 78070 12540
rect 77774 12486 77820 12538
rect 77820 12486 77830 12538
rect 77854 12486 77884 12538
rect 77884 12486 77896 12538
rect 77896 12486 77910 12538
rect 77934 12486 77948 12538
rect 77948 12486 77960 12538
rect 77960 12486 77990 12538
rect 78014 12486 78024 12538
rect 78024 12486 78070 12538
rect 77774 12484 77830 12486
rect 77854 12484 77910 12486
rect 77934 12484 77990 12486
rect 78014 12484 78070 12486
rect 86314 29280 86370 29336
rect 77774 11450 77830 11452
rect 77854 11450 77910 11452
rect 77934 11450 77990 11452
rect 78014 11450 78070 11452
rect 77774 11398 77820 11450
rect 77820 11398 77830 11450
rect 77854 11398 77884 11450
rect 77884 11398 77896 11450
rect 77896 11398 77910 11450
rect 77934 11398 77948 11450
rect 77948 11398 77960 11450
rect 77960 11398 77990 11450
rect 78014 11398 78024 11450
rect 78024 11398 78070 11450
rect 77774 11396 77830 11398
rect 77854 11396 77910 11398
rect 77934 11396 77990 11398
rect 78014 11396 78070 11398
rect 77774 10362 77830 10364
rect 77854 10362 77910 10364
rect 77934 10362 77990 10364
rect 78014 10362 78070 10364
rect 77774 10310 77820 10362
rect 77820 10310 77830 10362
rect 77854 10310 77884 10362
rect 77884 10310 77896 10362
rect 77896 10310 77910 10362
rect 77934 10310 77948 10362
rect 77948 10310 77960 10362
rect 77960 10310 77990 10362
rect 78014 10310 78024 10362
rect 78024 10310 78070 10362
rect 77774 10308 77830 10310
rect 77854 10308 77910 10310
rect 77934 10308 77990 10310
rect 78014 10308 78070 10310
rect 77774 9274 77830 9276
rect 77854 9274 77910 9276
rect 77934 9274 77990 9276
rect 78014 9274 78070 9276
rect 77774 9222 77820 9274
rect 77820 9222 77830 9274
rect 77854 9222 77884 9274
rect 77884 9222 77896 9274
rect 77896 9222 77910 9274
rect 77934 9222 77948 9274
rect 77948 9222 77960 9274
rect 77960 9222 77990 9274
rect 78014 9222 78024 9274
rect 78024 9222 78070 9274
rect 77774 9220 77830 9222
rect 77854 9220 77910 9222
rect 77934 9220 77990 9222
rect 78014 9220 78070 9222
rect 77774 8186 77830 8188
rect 77854 8186 77910 8188
rect 77934 8186 77990 8188
rect 78014 8186 78070 8188
rect 77774 8134 77820 8186
rect 77820 8134 77830 8186
rect 77854 8134 77884 8186
rect 77884 8134 77896 8186
rect 77896 8134 77910 8186
rect 77934 8134 77948 8186
rect 77948 8134 77960 8186
rect 77960 8134 77990 8186
rect 78014 8134 78024 8186
rect 78024 8134 78070 8186
rect 77774 8132 77830 8134
rect 77854 8132 77910 8134
rect 77934 8132 77990 8134
rect 78014 8132 78070 8134
rect 77774 7098 77830 7100
rect 77854 7098 77910 7100
rect 77934 7098 77990 7100
rect 78014 7098 78070 7100
rect 77774 7046 77820 7098
rect 77820 7046 77830 7098
rect 77854 7046 77884 7098
rect 77884 7046 77896 7098
rect 77896 7046 77910 7098
rect 77934 7046 77948 7098
rect 77948 7046 77960 7098
rect 77960 7046 77990 7098
rect 78014 7046 78024 7098
rect 78024 7046 78070 7098
rect 77774 7044 77830 7046
rect 77854 7044 77910 7046
rect 77934 7044 77990 7046
rect 78014 7044 78070 7046
rect 77774 6010 77830 6012
rect 77854 6010 77910 6012
rect 77934 6010 77990 6012
rect 78014 6010 78070 6012
rect 77774 5958 77820 6010
rect 77820 5958 77830 6010
rect 77854 5958 77884 6010
rect 77884 5958 77896 6010
rect 77896 5958 77910 6010
rect 77934 5958 77948 6010
rect 77948 5958 77960 6010
rect 77960 5958 77990 6010
rect 78014 5958 78024 6010
rect 78024 5958 78070 6010
rect 77774 5956 77830 5958
rect 77854 5956 77910 5958
rect 77934 5956 77990 5958
rect 78014 5956 78070 5958
rect 77774 4922 77830 4924
rect 77854 4922 77910 4924
rect 77934 4922 77990 4924
rect 78014 4922 78070 4924
rect 77774 4870 77820 4922
rect 77820 4870 77830 4922
rect 77854 4870 77884 4922
rect 77884 4870 77896 4922
rect 77896 4870 77910 4922
rect 77934 4870 77948 4922
rect 77948 4870 77960 4922
rect 77960 4870 77990 4922
rect 78014 4870 78024 4922
rect 78024 4870 78070 4922
rect 77774 4868 77830 4870
rect 77854 4868 77910 4870
rect 77934 4868 77990 4870
rect 78014 4868 78070 4870
rect 77774 3834 77830 3836
rect 77854 3834 77910 3836
rect 77934 3834 77990 3836
rect 78014 3834 78070 3836
rect 77774 3782 77820 3834
rect 77820 3782 77830 3834
rect 77854 3782 77884 3834
rect 77884 3782 77896 3834
rect 77896 3782 77910 3834
rect 77934 3782 77948 3834
rect 77948 3782 77960 3834
rect 77960 3782 77990 3834
rect 78014 3782 78024 3834
rect 78024 3782 78070 3834
rect 77774 3780 77830 3782
rect 77854 3780 77910 3782
rect 77934 3780 77990 3782
rect 78014 3780 78070 3782
rect 77774 2746 77830 2748
rect 77854 2746 77910 2748
rect 77934 2746 77990 2748
rect 78014 2746 78070 2748
rect 77774 2694 77820 2746
rect 77820 2694 77830 2746
rect 77854 2694 77884 2746
rect 77884 2694 77896 2746
rect 77896 2694 77910 2746
rect 77934 2694 77948 2746
rect 77948 2694 77960 2746
rect 77960 2694 77990 2746
rect 78014 2694 78024 2746
rect 78024 2694 78070 2746
rect 77774 2692 77830 2694
rect 77854 2692 77910 2694
rect 77934 2692 77990 2694
rect 78014 2692 78070 2694
rect 80794 2524 80796 2544
rect 80796 2524 80848 2544
rect 80848 2524 80850 2544
rect 80794 2488 80850 2524
rect 87510 27920 87566 27976
rect 86958 12688 87014 12744
rect 87418 26560 87474 26616
rect 87694 28600 87750 28656
rect 87970 27240 88026 27296
rect 87418 20440 87474 20496
rect 87878 25220 87934 25256
rect 87878 25200 87880 25220
rect 87880 25200 87932 25220
rect 87932 25200 87934 25220
rect 87786 12824 87842 12880
rect 87418 10920 87474 10976
rect 87418 8916 87420 8936
rect 87420 8916 87472 8936
rect 87472 8916 87474 8936
rect 87418 8880 87474 8916
rect 86866 856 86922 912
rect 87418 6196 87420 6216
rect 87420 6196 87472 6216
rect 87472 6196 87474 6216
rect 87418 6160 87474 6196
rect 88062 24556 88064 24576
rect 88064 24556 88116 24576
rect 88116 24556 88118 24576
rect 88062 24520 88118 24556
rect 88062 23840 88118 23896
rect 88062 23160 88118 23216
rect 88062 22480 88118 22536
rect 88062 21836 88064 21856
rect 88064 21836 88116 21856
rect 88116 21836 88118 21856
rect 88062 21800 88118 21836
rect 88062 21120 88118 21176
rect 88062 19760 88118 19816
rect 88062 19116 88064 19136
rect 88064 19116 88116 19136
rect 88116 19116 88118 19136
rect 88062 19080 88118 19116
rect 88246 18400 88302 18456
rect 88062 17060 88118 17096
rect 88062 17040 88064 17060
rect 88064 17040 88116 17060
rect 88116 17040 88118 17060
rect 88062 16396 88064 16416
rect 88064 16396 88116 16416
rect 88116 16396 88118 16416
rect 88062 16360 88118 16396
rect 88062 15680 88118 15736
rect 88062 15000 88118 15056
rect 88062 14340 88118 14376
rect 88062 14320 88064 14340
rect 88064 14320 88116 14340
rect 88116 14320 88118 14340
rect 87970 13912 88026 13968
rect 88062 13676 88064 13696
rect 88064 13676 88116 13696
rect 88116 13676 88118 13696
rect 88062 13640 88118 13676
rect 88062 12960 88118 13016
rect 88062 12280 88118 12336
rect 88062 11620 88118 11656
rect 88062 11600 88064 11620
rect 88064 11600 88116 11620
rect 88116 11600 88118 11620
rect 88062 10240 88118 10296
rect 88246 8200 88302 8256
rect 88062 7520 88118 7576
rect 88062 6840 88118 6896
rect 87970 5480 88026 5536
rect 88062 4800 88118 4856
rect 88062 4120 88118 4176
rect 88062 2760 88118 2816
rect 88154 2080 88210 2136
rect 88338 3440 88394 3496
rect 86682 40 86738 96
<< metal3 >>
rect 0 29338 800 29368
rect 86309 29338 86375 29341
rect 89200 29338 90000 29368
rect 0 29278 1456 29338
rect 0 29248 800 29278
rect 1396 29202 1456 29278
rect 86309 29336 90000 29338
rect 86309 29280 86314 29336
rect 86370 29280 90000 29336
rect 86309 29278 90000 29280
rect 86309 29275 86375 29278
rect 89200 29248 90000 29278
rect 2773 29202 2839 29205
rect 1396 29200 2839 29202
rect 1396 29144 2778 29200
rect 2834 29144 2839 29200
rect 1396 29142 2839 29144
rect 2773 29139 2839 29142
rect 0 28658 800 28688
rect 1761 28658 1827 28661
rect 0 28656 1827 28658
rect 0 28600 1766 28656
rect 1822 28600 1827 28656
rect 0 28598 1827 28600
rect 0 28568 800 28598
rect 1761 28595 1827 28598
rect 87689 28658 87755 28661
rect 89200 28658 90000 28688
rect 87689 28656 90000 28658
rect 87689 28600 87694 28656
rect 87750 28600 90000 28656
rect 87689 28598 90000 28600
rect 87689 28595 87755 28598
rect 89200 28568 90000 28598
rect 0 27978 800 28008
rect 1485 27978 1551 27981
rect 0 27976 1551 27978
rect 0 27920 1490 27976
rect 1546 27920 1551 27976
rect 0 27918 1551 27920
rect 0 27888 800 27918
rect 1485 27915 1551 27918
rect 87505 27978 87571 27981
rect 89200 27978 90000 28008
rect 87505 27976 90000 27978
rect 87505 27920 87510 27976
rect 87566 27920 90000 27976
rect 87505 27918 90000 27920
rect 87505 27915 87571 27918
rect 89200 27888 90000 27918
rect 11920 27776 12236 27777
rect 11920 27712 11926 27776
rect 11990 27712 12006 27776
rect 12070 27712 12086 27776
rect 12150 27712 12166 27776
rect 12230 27712 12236 27776
rect 11920 27711 12236 27712
rect 33868 27776 34184 27777
rect 33868 27712 33874 27776
rect 33938 27712 33954 27776
rect 34018 27712 34034 27776
rect 34098 27712 34114 27776
rect 34178 27712 34184 27776
rect 33868 27711 34184 27712
rect 55816 27776 56132 27777
rect 55816 27712 55822 27776
rect 55886 27712 55902 27776
rect 55966 27712 55982 27776
rect 56046 27712 56062 27776
rect 56126 27712 56132 27776
rect 55816 27711 56132 27712
rect 77764 27776 78080 27777
rect 77764 27712 77770 27776
rect 77834 27712 77850 27776
rect 77914 27712 77930 27776
rect 77994 27712 78010 27776
rect 78074 27712 78080 27776
rect 77764 27711 78080 27712
rect 25405 27434 25471 27437
rect 31201 27434 31267 27437
rect 25405 27432 31267 27434
rect 25405 27376 25410 27432
rect 25466 27376 31206 27432
rect 31262 27376 31267 27432
rect 25405 27374 31267 27376
rect 25405 27371 25471 27374
rect 31201 27371 31267 27374
rect 42609 27434 42675 27437
rect 46749 27434 46815 27437
rect 42609 27432 46815 27434
rect 42609 27376 42614 27432
rect 42670 27376 46754 27432
rect 46810 27376 46815 27432
rect 42609 27374 46815 27376
rect 42609 27371 42675 27374
rect 46749 27371 46815 27374
rect 0 27298 800 27328
rect 3049 27298 3115 27301
rect 0 27296 3115 27298
rect 0 27240 3054 27296
rect 3110 27240 3115 27296
rect 0 27238 3115 27240
rect 0 27208 800 27238
rect 3049 27235 3115 27238
rect 87965 27298 88031 27301
rect 89200 27298 90000 27328
rect 87965 27296 90000 27298
rect 87965 27240 87970 27296
rect 88026 27240 90000 27296
rect 87965 27238 90000 27240
rect 87965 27235 88031 27238
rect 22894 27232 23210 27233
rect 22894 27168 22900 27232
rect 22964 27168 22980 27232
rect 23044 27168 23060 27232
rect 23124 27168 23140 27232
rect 23204 27168 23210 27232
rect 22894 27167 23210 27168
rect 44842 27232 45158 27233
rect 44842 27168 44848 27232
rect 44912 27168 44928 27232
rect 44992 27168 45008 27232
rect 45072 27168 45088 27232
rect 45152 27168 45158 27232
rect 44842 27167 45158 27168
rect 66790 27232 67106 27233
rect 66790 27168 66796 27232
rect 66860 27168 66876 27232
rect 66940 27168 66956 27232
rect 67020 27168 67036 27232
rect 67100 27168 67106 27232
rect 89200 27208 90000 27238
rect 66790 27167 67106 27168
rect 40677 27026 40743 27029
rect 41781 27026 41847 27029
rect 40677 27024 41847 27026
rect 40677 26968 40682 27024
rect 40738 26968 41786 27024
rect 41842 26968 41847 27024
rect 40677 26966 41847 26968
rect 40677 26963 40743 26966
rect 41781 26963 41847 26966
rect 42701 27026 42767 27029
rect 44817 27026 44883 27029
rect 42701 27024 44883 27026
rect 42701 26968 42706 27024
rect 42762 26968 44822 27024
rect 44878 26968 44883 27024
rect 42701 26966 44883 26968
rect 42701 26963 42767 26966
rect 44817 26963 44883 26966
rect 29361 26890 29427 26893
rect 38193 26890 38259 26893
rect 29361 26888 38259 26890
rect 29361 26832 29366 26888
rect 29422 26832 38198 26888
rect 38254 26832 38259 26888
rect 29361 26830 38259 26832
rect 29361 26827 29427 26830
rect 38193 26827 38259 26830
rect 23381 26754 23447 26757
rect 27797 26754 27863 26757
rect 23381 26752 27863 26754
rect 23381 26696 23386 26752
rect 23442 26696 27802 26752
rect 27858 26696 27863 26752
rect 23381 26694 27863 26696
rect 23381 26691 23447 26694
rect 27797 26691 27863 26694
rect 11920 26688 12236 26689
rect 0 26618 800 26648
rect 11920 26624 11926 26688
rect 11990 26624 12006 26688
rect 12070 26624 12086 26688
rect 12150 26624 12166 26688
rect 12230 26624 12236 26688
rect 11920 26623 12236 26624
rect 33868 26688 34184 26689
rect 33868 26624 33874 26688
rect 33938 26624 33954 26688
rect 34018 26624 34034 26688
rect 34098 26624 34114 26688
rect 34178 26624 34184 26688
rect 33868 26623 34184 26624
rect 55816 26688 56132 26689
rect 55816 26624 55822 26688
rect 55886 26624 55902 26688
rect 55966 26624 55982 26688
rect 56046 26624 56062 26688
rect 56126 26624 56132 26688
rect 55816 26623 56132 26624
rect 77764 26688 78080 26689
rect 77764 26624 77770 26688
rect 77834 26624 77850 26688
rect 77914 26624 77930 26688
rect 77994 26624 78010 26688
rect 78074 26624 78080 26688
rect 77764 26623 78080 26624
rect 1669 26618 1735 26621
rect 0 26616 1735 26618
rect 0 26560 1674 26616
rect 1730 26560 1735 26616
rect 0 26558 1735 26560
rect 0 26528 800 26558
rect 1669 26555 1735 26558
rect 26417 26618 26483 26621
rect 27337 26618 27403 26621
rect 29637 26618 29703 26621
rect 26417 26616 29703 26618
rect 26417 26560 26422 26616
rect 26478 26560 27342 26616
rect 27398 26560 29642 26616
rect 29698 26560 29703 26616
rect 26417 26558 29703 26560
rect 26417 26555 26483 26558
rect 27337 26555 27403 26558
rect 29637 26555 29703 26558
rect 87413 26618 87479 26621
rect 89200 26618 90000 26648
rect 87413 26616 90000 26618
rect 87413 26560 87418 26616
rect 87474 26560 90000 26616
rect 87413 26558 90000 26560
rect 87413 26555 87479 26558
rect 89200 26528 90000 26558
rect 27521 26482 27587 26485
rect 33041 26482 33107 26485
rect 27521 26480 33107 26482
rect 27521 26424 27526 26480
rect 27582 26424 33046 26480
rect 33102 26424 33107 26480
rect 27521 26422 33107 26424
rect 27521 26419 27587 26422
rect 33041 26419 33107 26422
rect 40677 26346 40743 26349
rect 41689 26346 41755 26349
rect 40677 26344 41755 26346
rect 40677 26288 40682 26344
rect 40738 26288 41694 26344
rect 41750 26288 41755 26344
rect 40677 26286 41755 26288
rect 40677 26283 40743 26286
rect 41689 26283 41755 26286
rect 22894 26144 23210 26145
rect 22894 26080 22900 26144
rect 22964 26080 22980 26144
rect 23044 26080 23060 26144
rect 23124 26080 23140 26144
rect 23204 26080 23210 26144
rect 22894 26079 23210 26080
rect 44842 26144 45158 26145
rect 44842 26080 44848 26144
rect 44912 26080 44928 26144
rect 44992 26080 45008 26144
rect 45072 26080 45088 26144
rect 45152 26080 45158 26144
rect 44842 26079 45158 26080
rect 66790 26144 67106 26145
rect 66790 26080 66796 26144
rect 66860 26080 66876 26144
rect 66940 26080 66956 26144
rect 67020 26080 67036 26144
rect 67100 26080 67106 26144
rect 66790 26079 67106 26080
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 28022 25740 28028 25804
rect 28092 25802 28098 25804
rect 68921 25802 68987 25805
rect 28092 25800 68987 25802
rect 28092 25744 68926 25800
rect 68982 25744 68987 25800
rect 28092 25742 68987 25744
rect 28092 25740 28098 25742
rect 68921 25739 68987 25742
rect 11920 25600 12236 25601
rect 11920 25536 11926 25600
rect 11990 25536 12006 25600
rect 12070 25536 12086 25600
rect 12150 25536 12166 25600
rect 12230 25536 12236 25600
rect 11920 25535 12236 25536
rect 33868 25600 34184 25601
rect 33868 25536 33874 25600
rect 33938 25536 33954 25600
rect 34018 25536 34034 25600
rect 34098 25536 34114 25600
rect 34178 25536 34184 25600
rect 33868 25535 34184 25536
rect 55816 25600 56132 25601
rect 55816 25536 55822 25600
rect 55886 25536 55902 25600
rect 55966 25536 55982 25600
rect 56046 25536 56062 25600
rect 56126 25536 56132 25600
rect 55816 25535 56132 25536
rect 77764 25600 78080 25601
rect 77764 25536 77770 25600
rect 77834 25536 77850 25600
rect 77914 25536 77930 25600
rect 77994 25536 78010 25600
rect 78074 25536 78080 25600
rect 77764 25535 78080 25536
rect 0 25258 800 25288
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25168 800 25198
rect 1393 25195 1459 25198
rect 87873 25258 87939 25261
rect 89200 25258 90000 25288
rect 87873 25256 90000 25258
rect 87873 25200 87878 25256
rect 87934 25200 90000 25256
rect 87873 25198 90000 25200
rect 87873 25195 87939 25198
rect 89200 25168 90000 25198
rect 22894 25056 23210 25057
rect 22894 24992 22900 25056
rect 22964 24992 22980 25056
rect 23044 24992 23060 25056
rect 23124 24992 23140 25056
rect 23204 24992 23210 25056
rect 22894 24991 23210 24992
rect 44842 25056 45158 25057
rect 44842 24992 44848 25056
rect 44912 24992 44928 25056
rect 44992 24992 45008 25056
rect 45072 24992 45088 25056
rect 45152 24992 45158 25056
rect 44842 24991 45158 24992
rect 66790 25056 67106 25057
rect 66790 24992 66796 25056
rect 66860 24992 66876 25056
rect 66940 24992 66956 25056
rect 67020 24992 67036 25056
rect 67100 24992 67106 25056
rect 66790 24991 67106 24992
rect 0 24578 800 24608
rect 1393 24578 1459 24581
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 800 24518
rect 1393 24515 1459 24518
rect 88057 24578 88123 24581
rect 89200 24578 90000 24608
rect 88057 24576 90000 24578
rect 88057 24520 88062 24576
rect 88118 24520 90000 24576
rect 88057 24518 90000 24520
rect 88057 24515 88123 24518
rect 11920 24512 12236 24513
rect 11920 24448 11926 24512
rect 11990 24448 12006 24512
rect 12070 24448 12086 24512
rect 12150 24448 12166 24512
rect 12230 24448 12236 24512
rect 11920 24447 12236 24448
rect 33868 24512 34184 24513
rect 33868 24448 33874 24512
rect 33938 24448 33954 24512
rect 34018 24448 34034 24512
rect 34098 24448 34114 24512
rect 34178 24448 34184 24512
rect 33868 24447 34184 24448
rect 55816 24512 56132 24513
rect 55816 24448 55822 24512
rect 55886 24448 55902 24512
rect 55966 24448 55982 24512
rect 56046 24448 56062 24512
rect 56126 24448 56132 24512
rect 55816 24447 56132 24448
rect 77764 24512 78080 24513
rect 77764 24448 77770 24512
rect 77834 24448 77850 24512
rect 77914 24448 77930 24512
rect 77994 24448 78010 24512
rect 78074 24448 78080 24512
rect 89200 24488 90000 24518
rect 77764 24447 78080 24448
rect 27470 24108 27476 24172
rect 27540 24170 27546 24172
rect 80237 24170 80303 24173
rect 27540 24168 80303 24170
rect 27540 24112 80242 24168
rect 80298 24112 80303 24168
rect 27540 24110 80303 24112
rect 27540 24108 27546 24110
rect 80237 24107 80303 24110
rect 22894 23968 23210 23969
rect 22894 23904 22900 23968
rect 22964 23904 22980 23968
rect 23044 23904 23060 23968
rect 23124 23904 23140 23968
rect 23204 23904 23210 23968
rect 22894 23903 23210 23904
rect 44842 23968 45158 23969
rect 44842 23904 44848 23968
rect 44912 23904 44928 23968
rect 44992 23904 45008 23968
rect 45072 23904 45088 23968
rect 45152 23904 45158 23968
rect 44842 23903 45158 23904
rect 66790 23968 67106 23969
rect 66790 23904 66796 23968
rect 66860 23904 66876 23968
rect 66940 23904 66956 23968
rect 67020 23904 67036 23968
rect 67100 23904 67106 23968
rect 66790 23903 67106 23904
rect 88057 23898 88123 23901
rect 89200 23898 90000 23928
rect 88057 23896 90000 23898
rect 88057 23840 88062 23896
rect 88118 23840 90000 23896
rect 88057 23838 90000 23840
rect 88057 23835 88123 23838
rect 89200 23808 90000 23838
rect 11920 23424 12236 23425
rect 11920 23360 11926 23424
rect 11990 23360 12006 23424
rect 12070 23360 12086 23424
rect 12150 23360 12166 23424
rect 12230 23360 12236 23424
rect 11920 23359 12236 23360
rect 33868 23424 34184 23425
rect 33868 23360 33874 23424
rect 33938 23360 33954 23424
rect 34018 23360 34034 23424
rect 34098 23360 34114 23424
rect 34178 23360 34184 23424
rect 33868 23359 34184 23360
rect 55816 23424 56132 23425
rect 55816 23360 55822 23424
rect 55886 23360 55902 23424
rect 55966 23360 55982 23424
rect 56046 23360 56062 23424
rect 56126 23360 56132 23424
rect 55816 23359 56132 23360
rect 77764 23424 78080 23425
rect 77764 23360 77770 23424
rect 77834 23360 77850 23424
rect 77914 23360 77930 23424
rect 77994 23360 78010 23424
rect 78074 23360 78080 23424
rect 77764 23359 78080 23360
rect 0 23218 800 23248
rect 1761 23218 1827 23221
rect 0 23216 1827 23218
rect 0 23160 1766 23216
rect 1822 23160 1827 23216
rect 0 23158 1827 23160
rect 0 23128 800 23158
rect 1761 23155 1827 23158
rect 88057 23218 88123 23221
rect 89200 23218 90000 23248
rect 88057 23216 90000 23218
rect 88057 23160 88062 23216
rect 88118 23160 90000 23216
rect 88057 23158 90000 23160
rect 88057 23155 88123 23158
rect 89200 23128 90000 23158
rect 22894 22880 23210 22881
rect 22894 22816 22900 22880
rect 22964 22816 22980 22880
rect 23044 22816 23060 22880
rect 23124 22816 23140 22880
rect 23204 22816 23210 22880
rect 22894 22815 23210 22816
rect 44842 22880 45158 22881
rect 44842 22816 44848 22880
rect 44912 22816 44928 22880
rect 44992 22816 45008 22880
rect 45072 22816 45088 22880
rect 45152 22816 45158 22880
rect 44842 22815 45158 22816
rect 66790 22880 67106 22881
rect 66790 22816 66796 22880
rect 66860 22816 66876 22880
rect 66940 22816 66956 22880
rect 67020 22816 67036 22880
rect 67100 22816 67106 22880
rect 66790 22815 67106 22816
rect 31109 22674 31175 22677
rect 42149 22674 42215 22677
rect 31109 22672 42215 22674
rect 31109 22616 31114 22672
rect 31170 22616 42154 22672
rect 42210 22616 42215 22672
rect 31109 22614 42215 22616
rect 31109 22611 31175 22614
rect 42149 22611 42215 22614
rect 0 22538 800 22568
rect 1577 22538 1643 22541
rect 0 22536 1643 22538
rect 0 22480 1582 22536
rect 1638 22480 1643 22536
rect 0 22478 1643 22480
rect 0 22448 800 22478
rect 1577 22475 1643 22478
rect 88057 22538 88123 22541
rect 89200 22538 90000 22568
rect 88057 22536 90000 22538
rect 88057 22480 88062 22536
rect 88118 22480 90000 22536
rect 88057 22478 90000 22480
rect 88057 22475 88123 22478
rect 89200 22448 90000 22478
rect 11920 22336 12236 22337
rect 11920 22272 11926 22336
rect 11990 22272 12006 22336
rect 12070 22272 12086 22336
rect 12150 22272 12166 22336
rect 12230 22272 12236 22336
rect 11920 22271 12236 22272
rect 33868 22336 34184 22337
rect 33868 22272 33874 22336
rect 33938 22272 33954 22336
rect 34018 22272 34034 22336
rect 34098 22272 34114 22336
rect 34178 22272 34184 22336
rect 33868 22271 34184 22272
rect 55816 22336 56132 22337
rect 55816 22272 55822 22336
rect 55886 22272 55902 22336
rect 55966 22272 55982 22336
rect 56046 22272 56062 22336
rect 56126 22272 56132 22336
rect 55816 22271 56132 22272
rect 77764 22336 78080 22337
rect 77764 22272 77770 22336
rect 77834 22272 77850 22336
rect 77914 22272 77930 22336
rect 77994 22272 78010 22336
rect 78074 22272 78080 22336
rect 77764 22271 78080 22272
rect 0 21858 800 21888
rect 1393 21858 1459 21861
rect 0 21856 1459 21858
rect 0 21800 1398 21856
rect 1454 21800 1459 21856
rect 0 21798 1459 21800
rect 0 21768 800 21798
rect 1393 21795 1459 21798
rect 88057 21858 88123 21861
rect 89200 21858 90000 21888
rect 88057 21856 90000 21858
rect 88057 21800 88062 21856
rect 88118 21800 90000 21856
rect 88057 21798 90000 21800
rect 88057 21795 88123 21798
rect 22894 21792 23210 21793
rect 22894 21728 22900 21792
rect 22964 21728 22980 21792
rect 23044 21728 23060 21792
rect 23124 21728 23140 21792
rect 23204 21728 23210 21792
rect 22894 21727 23210 21728
rect 44842 21792 45158 21793
rect 44842 21728 44848 21792
rect 44912 21728 44928 21792
rect 44992 21728 45008 21792
rect 45072 21728 45088 21792
rect 45152 21728 45158 21792
rect 44842 21727 45158 21728
rect 66790 21792 67106 21793
rect 66790 21728 66796 21792
rect 66860 21728 66876 21792
rect 66940 21728 66956 21792
rect 67020 21728 67036 21792
rect 67100 21728 67106 21792
rect 89200 21768 90000 21798
rect 66790 21727 67106 21728
rect 26550 21388 26556 21452
rect 26620 21450 26626 21452
rect 59261 21450 59327 21453
rect 26620 21448 59327 21450
rect 26620 21392 59266 21448
rect 59322 21392 59327 21448
rect 26620 21390 59327 21392
rect 26620 21388 26626 21390
rect 59261 21387 59327 21390
rect 11920 21248 12236 21249
rect 0 21178 800 21208
rect 11920 21184 11926 21248
rect 11990 21184 12006 21248
rect 12070 21184 12086 21248
rect 12150 21184 12166 21248
rect 12230 21184 12236 21248
rect 11920 21183 12236 21184
rect 33868 21248 34184 21249
rect 33868 21184 33874 21248
rect 33938 21184 33954 21248
rect 34018 21184 34034 21248
rect 34098 21184 34114 21248
rect 34178 21184 34184 21248
rect 33868 21183 34184 21184
rect 55816 21248 56132 21249
rect 55816 21184 55822 21248
rect 55886 21184 55902 21248
rect 55966 21184 55982 21248
rect 56046 21184 56062 21248
rect 56126 21184 56132 21248
rect 55816 21183 56132 21184
rect 77764 21248 78080 21249
rect 77764 21184 77770 21248
rect 77834 21184 77850 21248
rect 77914 21184 77930 21248
rect 77994 21184 78010 21248
rect 78074 21184 78080 21248
rect 77764 21183 78080 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 800 21118
rect 1393 21115 1459 21118
rect 88057 21178 88123 21181
rect 89200 21178 90000 21208
rect 88057 21176 90000 21178
rect 88057 21120 88062 21176
rect 88118 21120 90000 21176
rect 88057 21118 90000 21120
rect 88057 21115 88123 21118
rect 89200 21088 90000 21118
rect 22894 20704 23210 20705
rect 22894 20640 22900 20704
rect 22964 20640 22980 20704
rect 23044 20640 23060 20704
rect 23124 20640 23140 20704
rect 23204 20640 23210 20704
rect 22894 20639 23210 20640
rect 44842 20704 45158 20705
rect 44842 20640 44848 20704
rect 44912 20640 44928 20704
rect 44992 20640 45008 20704
rect 45072 20640 45088 20704
rect 45152 20640 45158 20704
rect 44842 20639 45158 20640
rect 66790 20704 67106 20705
rect 66790 20640 66796 20704
rect 66860 20640 66876 20704
rect 66940 20640 66956 20704
rect 67020 20640 67036 20704
rect 67100 20640 67106 20704
rect 66790 20639 67106 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 87413 20498 87479 20501
rect 89200 20498 90000 20528
rect 87413 20496 90000 20498
rect 87413 20440 87418 20496
rect 87474 20440 90000 20496
rect 87413 20438 90000 20440
rect 87413 20435 87479 20438
rect 89200 20408 90000 20438
rect 11920 20160 12236 20161
rect 11920 20096 11926 20160
rect 11990 20096 12006 20160
rect 12070 20096 12086 20160
rect 12150 20096 12166 20160
rect 12230 20096 12236 20160
rect 11920 20095 12236 20096
rect 33868 20160 34184 20161
rect 33868 20096 33874 20160
rect 33938 20096 33954 20160
rect 34018 20096 34034 20160
rect 34098 20096 34114 20160
rect 34178 20096 34184 20160
rect 33868 20095 34184 20096
rect 55816 20160 56132 20161
rect 55816 20096 55822 20160
rect 55886 20096 55902 20160
rect 55966 20096 55982 20160
rect 56046 20096 56062 20160
rect 56126 20096 56132 20160
rect 55816 20095 56132 20096
rect 77764 20160 78080 20161
rect 77764 20096 77770 20160
rect 77834 20096 77850 20160
rect 77914 20096 77930 20160
rect 77994 20096 78010 20160
rect 78074 20096 78080 20160
rect 77764 20095 78080 20096
rect 0 19818 800 19848
rect 1393 19818 1459 19821
rect 0 19816 1459 19818
rect 0 19760 1398 19816
rect 1454 19760 1459 19816
rect 0 19758 1459 19760
rect 0 19728 800 19758
rect 1393 19755 1459 19758
rect 88057 19818 88123 19821
rect 89200 19818 90000 19848
rect 88057 19816 90000 19818
rect 88057 19760 88062 19816
rect 88118 19760 90000 19816
rect 88057 19758 90000 19760
rect 88057 19755 88123 19758
rect 89200 19728 90000 19758
rect 22894 19616 23210 19617
rect 22894 19552 22900 19616
rect 22964 19552 22980 19616
rect 23044 19552 23060 19616
rect 23124 19552 23140 19616
rect 23204 19552 23210 19616
rect 22894 19551 23210 19552
rect 44842 19616 45158 19617
rect 44842 19552 44848 19616
rect 44912 19552 44928 19616
rect 44992 19552 45008 19616
rect 45072 19552 45088 19616
rect 45152 19552 45158 19616
rect 44842 19551 45158 19552
rect 66790 19616 67106 19617
rect 66790 19552 66796 19616
rect 66860 19552 66876 19616
rect 66940 19552 66956 19616
rect 67020 19552 67036 19616
rect 67100 19552 67106 19616
rect 66790 19551 67106 19552
rect 0 19138 800 19168
rect 1761 19138 1827 19141
rect 0 19136 1827 19138
rect 0 19080 1766 19136
rect 1822 19080 1827 19136
rect 0 19078 1827 19080
rect 0 19048 800 19078
rect 1761 19075 1827 19078
rect 88057 19138 88123 19141
rect 89200 19138 90000 19168
rect 88057 19136 90000 19138
rect 88057 19080 88062 19136
rect 88118 19080 90000 19136
rect 88057 19078 90000 19080
rect 88057 19075 88123 19078
rect 11920 19072 12236 19073
rect 11920 19008 11926 19072
rect 11990 19008 12006 19072
rect 12070 19008 12086 19072
rect 12150 19008 12166 19072
rect 12230 19008 12236 19072
rect 11920 19007 12236 19008
rect 33868 19072 34184 19073
rect 33868 19008 33874 19072
rect 33938 19008 33954 19072
rect 34018 19008 34034 19072
rect 34098 19008 34114 19072
rect 34178 19008 34184 19072
rect 33868 19007 34184 19008
rect 55816 19072 56132 19073
rect 55816 19008 55822 19072
rect 55886 19008 55902 19072
rect 55966 19008 55982 19072
rect 56046 19008 56062 19072
rect 56126 19008 56132 19072
rect 55816 19007 56132 19008
rect 77764 19072 78080 19073
rect 77764 19008 77770 19072
rect 77834 19008 77850 19072
rect 77914 19008 77930 19072
rect 77994 19008 78010 19072
rect 78074 19008 78080 19072
rect 89200 19048 90000 19078
rect 77764 19007 78080 19008
rect 22894 18528 23210 18529
rect 0 18458 800 18488
rect 22894 18464 22900 18528
rect 22964 18464 22980 18528
rect 23044 18464 23060 18528
rect 23124 18464 23140 18528
rect 23204 18464 23210 18528
rect 22894 18463 23210 18464
rect 44842 18528 45158 18529
rect 44842 18464 44848 18528
rect 44912 18464 44928 18528
rect 44992 18464 45008 18528
rect 45072 18464 45088 18528
rect 45152 18464 45158 18528
rect 44842 18463 45158 18464
rect 66790 18528 67106 18529
rect 66790 18464 66796 18528
rect 66860 18464 66876 18528
rect 66940 18464 66956 18528
rect 67020 18464 67036 18528
rect 67100 18464 67106 18528
rect 66790 18463 67106 18464
rect 1393 18458 1459 18461
rect 0 18456 1459 18458
rect 0 18400 1398 18456
rect 1454 18400 1459 18456
rect 0 18398 1459 18400
rect 0 18368 800 18398
rect 1393 18395 1459 18398
rect 88241 18458 88307 18461
rect 89200 18458 90000 18488
rect 88241 18456 90000 18458
rect 88241 18400 88246 18456
rect 88302 18400 90000 18456
rect 88241 18398 90000 18400
rect 88241 18395 88307 18398
rect 89200 18368 90000 18398
rect 12249 18322 12315 18325
rect 36445 18322 36511 18325
rect 56317 18324 56383 18325
rect 56317 18322 56364 18324
rect 12249 18320 36511 18322
rect 12249 18264 12254 18320
rect 12310 18264 36450 18320
rect 36506 18264 36511 18320
rect 12249 18262 36511 18264
rect 56272 18320 56364 18322
rect 56272 18264 56322 18320
rect 56272 18262 56364 18264
rect 12249 18259 12315 18262
rect 36445 18259 36511 18262
rect 56317 18260 56364 18262
rect 56428 18260 56434 18324
rect 56317 18259 56383 18260
rect 50521 18186 50587 18189
rect 56409 18186 56475 18189
rect 50521 18184 56475 18186
rect 50521 18128 50526 18184
rect 50582 18128 56414 18184
rect 56470 18128 56475 18184
rect 50521 18126 56475 18128
rect 50521 18123 50587 18126
rect 56409 18123 56475 18126
rect 11920 17984 12236 17985
rect 11920 17920 11926 17984
rect 11990 17920 12006 17984
rect 12070 17920 12086 17984
rect 12150 17920 12166 17984
rect 12230 17920 12236 17984
rect 11920 17919 12236 17920
rect 33868 17984 34184 17985
rect 33868 17920 33874 17984
rect 33938 17920 33954 17984
rect 34018 17920 34034 17984
rect 34098 17920 34114 17984
rect 34178 17920 34184 17984
rect 33868 17919 34184 17920
rect 55816 17984 56132 17985
rect 55816 17920 55822 17984
rect 55886 17920 55902 17984
rect 55966 17920 55982 17984
rect 56046 17920 56062 17984
rect 56126 17920 56132 17984
rect 55816 17919 56132 17920
rect 77764 17984 78080 17985
rect 77764 17920 77770 17984
rect 77834 17920 77850 17984
rect 77914 17920 77930 17984
rect 77994 17920 78010 17984
rect 78074 17920 78080 17984
rect 77764 17919 78080 17920
rect 40677 17914 40743 17917
rect 45645 17914 45711 17917
rect 40677 17912 45711 17914
rect 40677 17856 40682 17912
rect 40738 17856 45650 17912
rect 45706 17856 45711 17912
rect 40677 17854 45711 17856
rect 40677 17851 40743 17854
rect 45645 17851 45711 17854
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 27153 17778 27219 17781
rect 28993 17778 29059 17781
rect 27153 17776 29059 17778
rect 27153 17720 27158 17776
rect 27214 17720 28998 17776
rect 29054 17720 29059 17776
rect 27153 17718 29059 17720
rect 27153 17715 27219 17718
rect 28993 17715 29059 17718
rect 41505 17778 41571 17781
rect 42241 17778 42307 17781
rect 41505 17776 42307 17778
rect 41505 17720 41510 17776
rect 41566 17720 42246 17776
rect 42302 17720 42307 17776
rect 41505 17718 42307 17720
rect 41505 17715 41571 17718
rect 42241 17715 42307 17718
rect 43437 17778 43503 17781
rect 46289 17778 46355 17781
rect 43437 17776 46355 17778
rect 43437 17720 43442 17776
rect 43498 17720 46294 17776
rect 46350 17720 46355 17776
rect 43437 17718 46355 17720
rect 43437 17715 43503 17718
rect 46289 17715 46355 17718
rect 55305 17778 55371 17781
rect 58617 17778 58683 17781
rect 55305 17776 58683 17778
rect 55305 17720 55310 17776
rect 55366 17720 58622 17776
rect 58678 17720 58683 17776
rect 55305 17718 58683 17720
rect 55305 17715 55371 17718
rect 58617 17715 58683 17718
rect 60457 17778 60523 17781
rect 60825 17778 60891 17781
rect 60457 17776 60891 17778
rect 60457 17720 60462 17776
rect 60518 17720 60830 17776
rect 60886 17720 60891 17776
rect 60457 17718 60891 17720
rect 60457 17715 60523 17718
rect 60825 17715 60891 17718
rect 22369 17642 22435 17645
rect 28441 17642 28507 17645
rect 46289 17642 46355 17645
rect 22369 17640 28507 17642
rect 22369 17584 22374 17640
rect 22430 17584 28446 17640
rect 28502 17584 28507 17640
rect 22369 17582 28507 17584
rect 22369 17579 22435 17582
rect 28441 17579 28507 17582
rect 38610 17640 46355 17642
rect 38610 17584 46294 17640
rect 46350 17584 46355 17640
rect 38610 17582 46355 17584
rect 24577 17506 24643 17509
rect 26325 17506 26391 17509
rect 24577 17504 26391 17506
rect 24577 17448 24582 17504
rect 24638 17448 26330 17504
rect 26386 17448 26391 17504
rect 24577 17446 26391 17448
rect 24577 17443 24643 17446
rect 26325 17443 26391 17446
rect 31109 17506 31175 17509
rect 32765 17506 32831 17509
rect 31109 17504 32831 17506
rect 31109 17448 31114 17504
rect 31170 17448 32770 17504
rect 32826 17448 32831 17504
rect 31109 17446 32831 17448
rect 31109 17443 31175 17446
rect 32765 17443 32831 17446
rect 22894 17440 23210 17441
rect 22894 17376 22900 17440
rect 22964 17376 22980 17440
rect 23044 17376 23060 17440
rect 23124 17376 23140 17440
rect 23204 17376 23210 17440
rect 22894 17375 23210 17376
rect 31753 17370 31819 17373
rect 38610 17370 38670 17582
rect 46289 17579 46355 17582
rect 46749 17642 46815 17645
rect 48129 17642 48195 17645
rect 46749 17640 48195 17642
rect 46749 17584 46754 17640
rect 46810 17584 48134 17640
rect 48190 17584 48195 17640
rect 46749 17582 48195 17584
rect 46749 17579 46815 17582
rect 48129 17579 48195 17582
rect 53005 17642 53071 17645
rect 56869 17642 56935 17645
rect 53005 17640 56935 17642
rect 53005 17584 53010 17640
rect 53066 17584 56874 17640
rect 56930 17584 56935 17640
rect 53005 17582 56935 17584
rect 53005 17579 53071 17582
rect 56869 17579 56935 17582
rect 64505 17642 64571 17645
rect 69105 17642 69171 17645
rect 64505 17640 69171 17642
rect 64505 17584 64510 17640
rect 64566 17584 69110 17640
rect 69166 17584 69171 17640
rect 64505 17582 69171 17584
rect 64505 17579 64571 17582
rect 69105 17579 69171 17582
rect 41321 17506 41387 17509
rect 41689 17506 41755 17509
rect 41321 17504 41755 17506
rect 41321 17448 41326 17504
rect 41382 17448 41694 17504
rect 41750 17448 41755 17504
rect 41321 17446 41755 17448
rect 41321 17443 41387 17446
rect 41689 17443 41755 17446
rect 48865 17506 48931 17509
rect 57881 17506 57947 17509
rect 48865 17504 57947 17506
rect 48865 17448 48870 17504
rect 48926 17448 57886 17504
rect 57942 17448 57947 17504
rect 48865 17446 57947 17448
rect 48865 17443 48931 17446
rect 57881 17443 57947 17446
rect 59077 17506 59143 17509
rect 62573 17506 62639 17509
rect 59077 17504 62639 17506
rect 59077 17448 59082 17504
rect 59138 17448 62578 17504
rect 62634 17448 62639 17504
rect 59077 17446 62639 17448
rect 59077 17443 59143 17446
rect 62573 17443 62639 17446
rect 44842 17440 45158 17441
rect 44842 17376 44848 17440
rect 44912 17376 44928 17440
rect 44992 17376 45008 17440
rect 45072 17376 45088 17440
rect 45152 17376 45158 17440
rect 44842 17375 45158 17376
rect 66790 17440 67106 17441
rect 66790 17376 66796 17440
rect 66860 17376 66876 17440
rect 66940 17376 66956 17440
rect 67020 17376 67036 17440
rect 67100 17376 67106 17440
rect 66790 17375 67106 17376
rect 31753 17368 38670 17370
rect 31753 17312 31758 17368
rect 31814 17312 38670 17368
rect 31753 17310 38670 17312
rect 45645 17370 45711 17373
rect 48681 17370 48747 17373
rect 49693 17370 49759 17373
rect 45645 17368 49759 17370
rect 45645 17312 45650 17368
rect 45706 17312 48686 17368
rect 48742 17312 49698 17368
rect 49754 17312 49759 17368
rect 45645 17310 49759 17312
rect 31753 17307 31819 17310
rect 45645 17307 45711 17310
rect 48681 17307 48747 17310
rect 49693 17307 49759 17310
rect 50061 17370 50127 17373
rect 54477 17370 54543 17373
rect 50061 17368 54543 17370
rect 50061 17312 50066 17368
rect 50122 17312 54482 17368
rect 54538 17312 54543 17368
rect 50061 17310 54543 17312
rect 50061 17307 50127 17310
rect 54477 17307 54543 17310
rect 60273 17370 60339 17373
rect 66529 17370 66595 17373
rect 60273 17368 66595 17370
rect 60273 17312 60278 17368
rect 60334 17312 66534 17368
rect 66590 17312 66595 17368
rect 60273 17310 66595 17312
rect 60273 17307 60339 17310
rect 66529 17307 66595 17310
rect 33593 17234 33659 17237
rect 35065 17234 35131 17237
rect 37641 17234 37707 17237
rect 33593 17232 37707 17234
rect 33593 17176 33598 17232
rect 33654 17176 35070 17232
rect 35126 17176 37646 17232
rect 37702 17176 37707 17232
rect 33593 17174 37707 17176
rect 33593 17171 33659 17174
rect 35065 17171 35131 17174
rect 37641 17171 37707 17174
rect 40493 17234 40559 17237
rect 47853 17234 47919 17237
rect 40493 17232 47919 17234
rect 40493 17176 40498 17232
rect 40554 17176 47858 17232
rect 47914 17176 47919 17232
rect 40493 17174 47919 17176
rect 40493 17171 40559 17174
rect 47853 17171 47919 17174
rect 49417 17234 49483 17237
rect 56777 17234 56843 17237
rect 49417 17232 56843 17234
rect 49417 17176 49422 17232
rect 49478 17176 56782 17232
rect 56838 17176 56843 17232
rect 49417 17174 56843 17176
rect 49417 17171 49483 17174
rect 56777 17171 56843 17174
rect 58617 17234 58683 17237
rect 66989 17234 67055 17237
rect 58617 17232 67055 17234
rect 58617 17176 58622 17232
rect 58678 17176 66994 17232
rect 67050 17176 67055 17232
rect 58617 17174 67055 17176
rect 58617 17171 58683 17174
rect 66989 17171 67055 17174
rect 0 17098 800 17128
rect 1761 17098 1827 17101
rect 0 17096 1827 17098
rect 0 17040 1766 17096
rect 1822 17040 1827 17096
rect 0 17038 1827 17040
rect 0 17008 800 17038
rect 1761 17035 1827 17038
rect 24669 17098 24735 17101
rect 28349 17098 28415 17101
rect 24669 17096 28415 17098
rect 24669 17040 24674 17096
rect 24730 17040 28354 17096
rect 28410 17040 28415 17096
rect 24669 17038 28415 17040
rect 24669 17035 24735 17038
rect 28349 17035 28415 17038
rect 42333 17098 42399 17101
rect 49969 17098 50035 17101
rect 42333 17096 50035 17098
rect 42333 17040 42338 17096
rect 42394 17040 49974 17096
rect 50030 17040 50035 17096
rect 42333 17038 50035 17040
rect 42333 17035 42399 17038
rect 49969 17035 50035 17038
rect 58801 17098 58867 17101
rect 60641 17098 60707 17101
rect 58801 17096 60707 17098
rect 58801 17040 58806 17096
rect 58862 17040 60646 17096
rect 60702 17040 60707 17096
rect 58801 17038 60707 17040
rect 58801 17035 58867 17038
rect 60641 17035 60707 17038
rect 66437 17098 66503 17101
rect 69289 17098 69355 17101
rect 66437 17096 69355 17098
rect 66437 17040 66442 17096
rect 66498 17040 69294 17096
rect 69350 17040 69355 17096
rect 66437 17038 69355 17040
rect 66437 17035 66503 17038
rect 69289 17035 69355 17038
rect 88057 17098 88123 17101
rect 89200 17098 90000 17128
rect 88057 17096 90000 17098
rect 88057 17040 88062 17096
rect 88118 17040 90000 17096
rect 88057 17038 90000 17040
rect 88057 17035 88123 17038
rect 89200 17008 90000 17038
rect 21817 16962 21883 16965
rect 28257 16962 28323 16965
rect 28533 16962 28599 16965
rect 21817 16960 28599 16962
rect 21817 16904 21822 16960
rect 21878 16904 28262 16960
rect 28318 16904 28538 16960
rect 28594 16904 28599 16960
rect 21817 16902 28599 16904
rect 21817 16899 21883 16902
rect 28257 16899 28323 16902
rect 28533 16899 28599 16902
rect 45921 16962 45987 16965
rect 50981 16962 51047 16965
rect 45921 16960 51047 16962
rect 45921 16904 45926 16960
rect 45982 16904 50986 16960
rect 51042 16904 51047 16960
rect 45921 16902 51047 16904
rect 45921 16899 45987 16902
rect 50981 16899 51047 16902
rect 53465 16962 53531 16965
rect 54661 16962 54727 16965
rect 53465 16960 54727 16962
rect 53465 16904 53470 16960
rect 53526 16904 54666 16960
rect 54722 16904 54727 16960
rect 53465 16902 54727 16904
rect 53465 16899 53531 16902
rect 54661 16899 54727 16902
rect 64689 16962 64755 16965
rect 66253 16962 66319 16965
rect 69565 16962 69631 16965
rect 64689 16960 69631 16962
rect 64689 16904 64694 16960
rect 64750 16904 66258 16960
rect 66314 16904 69570 16960
rect 69626 16904 69631 16960
rect 64689 16902 69631 16904
rect 64689 16899 64755 16902
rect 66253 16899 66319 16902
rect 69565 16899 69631 16902
rect 11920 16896 12236 16897
rect 11920 16832 11926 16896
rect 11990 16832 12006 16896
rect 12070 16832 12086 16896
rect 12150 16832 12166 16896
rect 12230 16832 12236 16896
rect 11920 16831 12236 16832
rect 33868 16896 34184 16897
rect 33868 16832 33874 16896
rect 33938 16832 33954 16896
rect 34018 16832 34034 16896
rect 34098 16832 34114 16896
rect 34178 16832 34184 16896
rect 33868 16831 34184 16832
rect 55816 16896 56132 16897
rect 55816 16832 55822 16896
rect 55886 16832 55902 16896
rect 55966 16832 55982 16896
rect 56046 16832 56062 16896
rect 56126 16832 56132 16896
rect 55816 16831 56132 16832
rect 77764 16896 78080 16897
rect 77764 16832 77770 16896
rect 77834 16832 77850 16896
rect 77914 16832 77930 16896
rect 77994 16832 78010 16896
rect 78074 16832 78080 16896
rect 77764 16831 78080 16832
rect 25865 16826 25931 16829
rect 28073 16826 28139 16829
rect 25865 16824 28139 16826
rect 25865 16768 25870 16824
rect 25926 16768 28078 16824
rect 28134 16768 28139 16824
rect 25865 16766 28139 16768
rect 25865 16763 25931 16766
rect 28073 16763 28139 16766
rect 39573 16826 39639 16829
rect 42333 16826 42399 16829
rect 39573 16824 42399 16826
rect 39573 16768 39578 16824
rect 39634 16768 42338 16824
rect 42394 16768 42399 16824
rect 39573 16766 42399 16768
rect 39573 16763 39639 16766
rect 42333 16763 42399 16766
rect 48129 16826 48195 16829
rect 50245 16826 50311 16829
rect 51901 16826 51967 16829
rect 55397 16826 55463 16829
rect 48129 16824 48882 16826
rect 48129 16768 48134 16824
rect 48190 16768 48882 16824
rect 48129 16766 48882 16768
rect 48129 16763 48195 16766
rect 38745 16690 38811 16693
rect 42977 16690 43043 16693
rect 38745 16688 43043 16690
rect 38745 16632 38750 16688
rect 38806 16632 42982 16688
rect 43038 16632 43043 16688
rect 38745 16630 43043 16632
rect 38745 16627 38811 16630
rect 42977 16627 43043 16630
rect 44725 16690 44791 16693
rect 48405 16690 48471 16693
rect 44725 16688 48471 16690
rect 44725 16632 44730 16688
rect 44786 16632 48410 16688
rect 48466 16632 48471 16688
rect 44725 16630 48471 16632
rect 48822 16690 48882 16766
rect 50245 16824 51967 16826
rect 50245 16768 50250 16824
rect 50306 16768 51906 16824
rect 51962 16768 51967 16824
rect 50245 16766 51967 16768
rect 50245 16763 50311 16766
rect 51901 16763 51967 16766
rect 52088 16824 55463 16826
rect 52088 16768 55402 16824
rect 55458 16768 55463 16824
rect 52088 16766 55463 16768
rect 50613 16690 50679 16693
rect 48822 16688 50679 16690
rect 48822 16632 50618 16688
rect 50674 16632 50679 16688
rect 48822 16630 50679 16632
rect 44725 16627 44791 16630
rect 48405 16627 48471 16630
rect 50613 16627 50679 16630
rect 34329 16554 34395 16557
rect 47577 16554 47643 16557
rect 34329 16552 47643 16554
rect 34329 16496 34334 16552
rect 34390 16496 47582 16552
rect 47638 16496 47643 16552
rect 34329 16494 47643 16496
rect 34329 16491 34395 16494
rect 47577 16491 47643 16494
rect 48129 16554 48195 16557
rect 52088 16554 52148 16766
rect 55397 16763 55463 16766
rect 58893 16826 58959 16829
rect 63309 16826 63375 16829
rect 58893 16824 63375 16826
rect 58893 16768 58898 16824
rect 58954 16768 63314 16824
rect 63370 16768 63375 16824
rect 58893 16766 63375 16768
rect 58893 16763 58959 16766
rect 63309 16763 63375 16766
rect 57421 16690 57487 16693
rect 48129 16552 52148 16554
rect 48129 16496 48134 16552
rect 48190 16496 52148 16552
rect 48129 16494 52148 16496
rect 52640 16688 57487 16690
rect 52640 16632 57426 16688
rect 57482 16632 57487 16688
rect 52640 16630 57487 16632
rect 48129 16491 48195 16494
rect 0 16418 800 16448
rect 1393 16418 1459 16421
rect 0 16416 1459 16418
rect 0 16360 1398 16416
rect 1454 16360 1459 16416
rect 0 16358 1459 16360
rect 0 16328 800 16358
rect 1393 16355 1459 16358
rect 46197 16418 46263 16421
rect 48037 16418 48103 16421
rect 46197 16416 48103 16418
rect 46197 16360 46202 16416
rect 46258 16360 48042 16416
rect 48098 16360 48103 16416
rect 46197 16358 48103 16360
rect 46197 16355 46263 16358
rect 48037 16355 48103 16358
rect 51349 16418 51415 16421
rect 52640 16418 52700 16630
rect 57421 16627 57487 16630
rect 59537 16690 59603 16693
rect 63033 16690 63099 16693
rect 59537 16688 63099 16690
rect 59537 16632 59542 16688
rect 59598 16632 63038 16688
rect 63094 16632 63099 16688
rect 59537 16630 63099 16632
rect 59537 16627 59603 16630
rect 63033 16627 63099 16630
rect 52821 16554 52887 16557
rect 57513 16554 57579 16557
rect 52821 16552 57579 16554
rect 52821 16496 52826 16552
rect 52882 16496 57518 16552
rect 57574 16496 57579 16552
rect 52821 16494 57579 16496
rect 52821 16491 52887 16494
rect 57513 16491 57579 16494
rect 58893 16554 58959 16557
rect 66437 16554 66503 16557
rect 58893 16552 66503 16554
rect 58893 16496 58898 16552
rect 58954 16496 66442 16552
rect 66498 16496 66503 16552
rect 58893 16494 66503 16496
rect 58893 16491 58959 16494
rect 66437 16491 66503 16494
rect 51349 16416 52700 16418
rect 51349 16360 51354 16416
rect 51410 16360 52700 16416
rect 51349 16358 52700 16360
rect 54477 16418 54543 16421
rect 60733 16418 60799 16421
rect 54477 16416 60799 16418
rect 54477 16360 54482 16416
rect 54538 16360 60738 16416
rect 60794 16360 60799 16416
rect 54477 16358 60799 16360
rect 51349 16355 51415 16358
rect 54477 16355 54543 16358
rect 60733 16355 60799 16358
rect 88057 16418 88123 16421
rect 89200 16418 90000 16448
rect 88057 16416 90000 16418
rect 88057 16360 88062 16416
rect 88118 16360 90000 16416
rect 88057 16358 90000 16360
rect 88057 16355 88123 16358
rect 22894 16352 23210 16353
rect 22894 16288 22900 16352
rect 22964 16288 22980 16352
rect 23044 16288 23060 16352
rect 23124 16288 23140 16352
rect 23204 16288 23210 16352
rect 22894 16287 23210 16288
rect 44842 16352 45158 16353
rect 44842 16288 44848 16352
rect 44912 16288 44928 16352
rect 44992 16288 45008 16352
rect 45072 16288 45088 16352
rect 45152 16288 45158 16352
rect 44842 16287 45158 16288
rect 66790 16352 67106 16353
rect 66790 16288 66796 16352
rect 66860 16288 66876 16352
rect 66940 16288 66956 16352
rect 67020 16288 67036 16352
rect 67100 16288 67106 16352
rect 89200 16328 90000 16358
rect 66790 16287 67106 16288
rect 25037 16282 25103 16285
rect 25773 16282 25839 16285
rect 26141 16282 26207 16285
rect 26969 16282 27035 16285
rect 28257 16282 28323 16285
rect 25037 16280 28323 16282
rect 25037 16224 25042 16280
rect 25098 16224 25778 16280
rect 25834 16224 26146 16280
rect 26202 16224 26974 16280
rect 27030 16224 28262 16280
rect 28318 16224 28323 16280
rect 25037 16222 28323 16224
rect 25037 16219 25103 16222
rect 25773 16219 25839 16222
rect 26141 16219 26207 16222
rect 26969 16219 27035 16222
rect 28257 16219 28323 16222
rect 46657 16282 46723 16285
rect 48221 16282 48287 16285
rect 46657 16280 48287 16282
rect 46657 16224 46662 16280
rect 46718 16224 48226 16280
rect 48282 16224 48287 16280
rect 46657 16222 48287 16224
rect 46657 16219 46723 16222
rect 48221 16219 48287 16222
rect 49601 16282 49667 16285
rect 53189 16282 53255 16285
rect 49601 16280 53255 16282
rect 49601 16224 49606 16280
rect 49662 16224 53194 16280
rect 53250 16224 53255 16280
rect 49601 16222 53255 16224
rect 49601 16219 49667 16222
rect 53189 16219 53255 16222
rect 53741 16282 53807 16285
rect 58617 16282 58683 16285
rect 53741 16280 58683 16282
rect 53741 16224 53746 16280
rect 53802 16224 58622 16280
rect 58678 16224 58683 16280
rect 53741 16222 58683 16224
rect 53741 16219 53807 16222
rect 58617 16219 58683 16222
rect 26049 16146 26115 16149
rect 46381 16146 46447 16149
rect 55489 16146 55555 16149
rect 26049 16144 46447 16146
rect 26049 16088 26054 16144
rect 26110 16088 46386 16144
rect 46442 16088 46447 16144
rect 26049 16086 46447 16088
rect 26049 16083 26115 16086
rect 46381 16083 46447 16086
rect 51030 16144 55555 16146
rect 51030 16088 55494 16144
rect 55550 16088 55555 16144
rect 51030 16086 55555 16088
rect 27337 16010 27403 16013
rect 27705 16010 27771 16013
rect 27337 16008 27771 16010
rect 27337 15952 27342 16008
rect 27398 15952 27710 16008
rect 27766 15952 27771 16008
rect 27337 15950 27771 15952
rect 27337 15947 27403 15950
rect 27705 15947 27771 15950
rect 29177 16010 29243 16013
rect 51030 16010 51090 16086
rect 55489 16083 55555 16086
rect 55622 16084 55628 16148
rect 55692 16146 55698 16148
rect 57973 16146 58039 16149
rect 55692 16144 58039 16146
rect 55692 16088 57978 16144
rect 58034 16088 58039 16144
rect 55692 16086 58039 16088
rect 55692 16084 55698 16086
rect 57973 16083 58039 16086
rect 58249 16146 58315 16149
rect 66069 16146 66135 16149
rect 58249 16144 66135 16146
rect 58249 16088 58254 16144
rect 58310 16088 66074 16144
rect 66130 16088 66135 16144
rect 58249 16086 66135 16088
rect 58249 16083 58315 16086
rect 66069 16083 66135 16086
rect 29177 16008 51090 16010
rect 29177 15952 29182 16008
rect 29238 15952 51090 16008
rect 29177 15950 51090 15952
rect 51165 16010 51231 16013
rect 52821 16010 52887 16013
rect 51165 16008 52887 16010
rect 51165 15952 51170 16008
rect 51226 15952 52826 16008
rect 52882 15952 52887 16008
rect 51165 15950 52887 15952
rect 29177 15947 29243 15950
rect 51165 15947 51231 15950
rect 52821 15947 52887 15950
rect 53925 16010 53991 16013
rect 55673 16010 55739 16013
rect 56593 16010 56659 16013
rect 53925 16008 56659 16010
rect 53925 15952 53930 16008
rect 53986 15952 55678 16008
rect 55734 15952 56598 16008
rect 56654 15952 56659 16008
rect 53925 15950 56659 15952
rect 53925 15947 53991 15950
rect 55673 15947 55739 15950
rect 56593 15947 56659 15950
rect 57973 16010 58039 16013
rect 59261 16010 59327 16013
rect 57973 16008 59327 16010
rect 57973 15952 57978 16008
rect 58034 15952 59266 16008
rect 59322 15952 59327 16008
rect 57973 15950 59327 15952
rect 57973 15947 58039 15950
rect 59261 15947 59327 15950
rect 25405 15874 25471 15877
rect 27797 15874 27863 15877
rect 25405 15872 27863 15874
rect 25405 15816 25410 15872
rect 25466 15816 27802 15872
rect 27858 15816 27863 15872
rect 25405 15814 27863 15816
rect 25405 15811 25471 15814
rect 27797 15811 27863 15814
rect 30557 15874 30623 15877
rect 33133 15874 33199 15877
rect 30557 15872 33199 15874
rect 30557 15816 30562 15872
rect 30618 15816 33138 15872
rect 33194 15816 33199 15872
rect 30557 15814 33199 15816
rect 30557 15811 30623 15814
rect 33133 15811 33199 15814
rect 42885 15874 42951 15877
rect 43897 15874 43963 15877
rect 46841 15874 46907 15877
rect 49417 15874 49483 15877
rect 42885 15872 49483 15874
rect 42885 15816 42890 15872
rect 42946 15816 43902 15872
rect 43958 15816 46846 15872
rect 46902 15816 49422 15872
rect 49478 15816 49483 15872
rect 42885 15814 49483 15816
rect 42885 15811 42951 15814
rect 43897 15811 43963 15814
rect 46841 15811 46907 15814
rect 49417 15811 49483 15814
rect 50153 15874 50219 15877
rect 54937 15874 55003 15877
rect 50153 15872 55003 15874
rect 50153 15816 50158 15872
rect 50214 15816 54942 15872
rect 54998 15816 55003 15872
rect 50153 15814 55003 15816
rect 50153 15811 50219 15814
rect 54937 15811 55003 15814
rect 11920 15808 12236 15809
rect 11920 15744 11926 15808
rect 11990 15744 12006 15808
rect 12070 15744 12086 15808
rect 12150 15744 12166 15808
rect 12230 15744 12236 15808
rect 11920 15743 12236 15744
rect 33868 15808 34184 15809
rect 33868 15744 33874 15808
rect 33938 15744 33954 15808
rect 34018 15744 34034 15808
rect 34098 15744 34114 15808
rect 34178 15744 34184 15808
rect 33868 15743 34184 15744
rect 55816 15808 56132 15809
rect 55816 15744 55822 15808
rect 55886 15744 55902 15808
rect 55966 15744 55982 15808
rect 56046 15744 56062 15808
rect 56126 15744 56132 15808
rect 55816 15743 56132 15744
rect 77764 15808 78080 15809
rect 77764 15744 77770 15808
rect 77834 15744 77850 15808
rect 77914 15744 77930 15808
rect 77994 15744 78010 15808
rect 78074 15744 78080 15808
rect 77764 15743 78080 15744
rect 24209 15738 24275 15741
rect 27429 15738 27495 15741
rect 33593 15738 33659 15741
rect 24209 15736 33659 15738
rect 24209 15680 24214 15736
rect 24270 15680 27434 15736
rect 27490 15680 33598 15736
rect 33654 15680 33659 15736
rect 24209 15678 33659 15680
rect 24209 15675 24275 15678
rect 27429 15675 27495 15678
rect 33593 15675 33659 15678
rect 42609 15738 42675 15741
rect 48221 15738 48287 15741
rect 42609 15736 48287 15738
rect 42609 15680 42614 15736
rect 42670 15680 48226 15736
rect 48282 15680 48287 15736
rect 42609 15678 48287 15680
rect 42609 15675 42675 15678
rect 48221 15675 48287 15678
rect 48497 15738 48563 15741
rect 53465 15738 53531 15741
rect 54753 15738 54819 15741
rect 48497 15736 54819 15738
rect 48497 15680 48502 15736
rect 48558 15680 53470 15736
rect 53526 15680 54758 15736
rect 54814 15680 54819 15736
rect 48497 15678 54819 15680
rect 48497 15675 48563 15678
rect 53465 15675 53531 15678
rect 54753 15675 54819 15678
rect 88057 15738 88123 15741
rect 89200 15738 90000 15768
rect 88057 15736 90000 15738
rect 88057 15680 88062 15736
rect 88118 15680 90000 15736
rect 88057 15678 90000 15680
rect 88057 15675 88123 15678
rect 89200 15648 90000 15678
rect 27889 15602 27955 15605
rect 28022 15602 28028 15604
rect 27889 15600 28028 15602
rect 27889 15544 27894 15600
rect 27950 15544 28028 15600
rect 27889 15542 28028 15544
rect 27889 15539 27955 15542
rect 28022 15540 28028 15542
rect 28092 15540 28098 15604
rect 31937 15602 32003 15605
rect 32489 15602 32555 15605
rect 31937 15600 32555 15602
rect 31937 15544 31942 15600
rect 31998 15544 32494 15600
rect 32550 15544 32555 15600
rect 31937 15542 32555 15544
rect 31937 15539 32003 15542
rect 32489 15539 32555 15542
rect 44265 15602 44331 15605
rect 48037 15602 48103 15605
rect 44265 15600 48103 15602
rect 44265 15544 44270 15600
rect 44326 15544 48042 15600
rect 48098 15544 48103 15600
rect 44265 15542 48103 15544
rect 44265 15539 44331 15542
rect 48037 15539 48103 15542
rect 49969 15602 50035 15605
rect 51993 15602 52059 15605
rect 49969 15600 52059 15602
rect 49969 15544 49974 15600
rect 50030 15544 51998 15600
rect 52054 15544 52059 15600
rect 49969 15542 52059 15544
rect 49969 15539 50035 15542
rect 51993 15539 52059 15542
rect 52269 15602 52335 15605
rect 56317 15602 56383 15605
rect 52269 15600 56383 15602
rect 52269 15544 52274 15600
rect 52330 15544 56322 15600
rect 56378 15544 56383 15600
rect 52269 15542 56383 15544
rect 52269 15539 52335 15542
rect 56317 15539 56383 15542
rect 58617 15602 58683 15605
rect 62205 15602 62271 15605
rect 62665 15602 62731 15605
rect 58617 15600 62731 15602
rect 58617 15544 58622 15600
rect 58678 15544 62210 15600
rect 62266 15544 62670 15600
rect 62726 15544 62731 15600
rect 58617 15542 62731 15544
rect 58617 15539 58683 15542
rect 62205 15539 62271 15542
rect 62665 15539 62731 15542
rect 63309 15600 63375 15605
rect 63309 15544 63314 15600
rect 63370 15544 63375 15600
rect 63309 15539 63375 15544
rect 15101 15466 15167 15469
rect 61837 15466 61903 15469
rect 15101 15464 61903 15466
rect 15101 15408 15106 15464
rect 15162 15408 61842 15464
rect 61898 15408 61903 15464
rect 15101 15406 61903 15408
rect 15101 15403 15167 15406
rect 61837 15403 61903 15406
rect 23381 15330 23447 15333
rect 28901 15330 28967 15333
rect 23381 15328 28967 15330
rect 23381 15272 23386 15328
rect 23442 15272 28906 15328
rect 28962 15272 28967 15328
rect 23381 15270 28967 15272
rect 23381 15267 23447 15270
rect 28901 15267 28967 15270
rect 48313 15330 48379 15333
rect 48773 15330 48839 15333
rect 51073 15330 51139 15333
rect 48313 15328 51139 15330
rect 48313 15272 48318 15328
rect 48374 15272 48778 15328
rect 48834 15272 51078 15328
rect 51134 15272 51139 15328
rect 48313 15270 51139 15272
rect 48313 15267 48379 15270
rect 48773 15267 48839 15270
rect 51073 15267 51139 15270
rect 51441 15330 51507 15333
rect 52545 15330 52611 15333
rect 51441 15328 52611 15330
rect 51441 15272 51446 15328
rect 51502 15272 52550 15328
rect 52606 15272 52611 15328
rect 51441 15270 52611 15272
rect 51441 15267 51507 15270
rect 52545 15267 52611 15270
rect 60549 15330 60615 15333
rect 63125 15330 63191 15333
rect 60549 15328 63191 15330
rect 60549 15272 60554 15328
rect 60610 15272 63130 15328
rect 63186 15272 63191 15328
rect 60549 15270 63191 15272
rect 63312 15330 63372 15539
rect 63769 15330 63835 15333
rect 63312 15328 63835 15330
rect 63312 15272 63774 15328
rect 63830 15272 63835 15328
rect 63312 15270 63835 15272
rect 60549 15267 60615 15270
rect 63125 15267 63191 15270
rect 63769 15267 63835 15270
rect 22894 15264 23210 15265
rect 22894 15200 22900 15264
rect 22964 15200 22980 15264
rect 23044 15200 23060 15264
rect 23124 15200 23140 15264
rect 23204 15200 23210 15264
rect 22894 15199 23210 15200
rect 44842 15264 45158 15265
rect 44842 15200 44848 15264
rect 44912 15200 44928 15264
rect 44992 15200 45008 15264
rect 45072 15200 45088 15264
rect 45152 15200 45158 15264
rect 44842 15199 45158 15200
rect 66790 15264 67106 15265
rect 66790 15200 66796 15264
rect 66860 15200 66876 15264
rect 66940 15200 66956 15264
rect 67020 15200 67036 15264
rect 67100 15200 67106 15264
rect 66790 15199 67106 15200
rect 27337 15194 27403 15197
rect 27470 15194 27476 15196
rect 27337 15192 27476 15194
rect 27337 15136 27342 15192
rect 27398 15136 27476 15192
rect 27337 15134 27476 15136
rect 27337 15131 27403 15134
rect 27470 15132 27476 15134
rect 27540 15132 27546 15196
rect 31477 15194 31543 15197
rect 36169 15194 36235 15197
rect 31477 15192 36235 15194
rect 31477 15136 31482 15192
rect 31538 15136 36174 15192
rect 36230 15136 36235 15192
rect 31477 15134 36235 15136
rect 31477 15131 31543 15134
rect 36169 15131 36235 15134
rect 39297 15194 39363 15197
rect 40769 15194 40835 15197
rect 44633 15194 44699 15197
rect 39297 15192 44699 15194
rect 39297 15136 39302 15192
rect 39358 15136 40774 15192
rect 40830 15136 44638 15192
rect 44694 15136 44699 15192
rect 39297 15134 44699 15136
rect 39297 15131 39363 15134
rect 40769 15131 40835 15134
rect 44633 15131 44699 15134
rect 46841 15194 46907 15197
rect 50981 15194 51047 15197
rect 46841 15192 51047 15194
rect 46841 15136 46846 15192
rect 46902 15136 50986 15192
rect 51042 15136 51047 15192
rect 46841 15134 51047 15136
rect 46841 15131 46907 15134
rect 50981 15131 51047 15134
rect 53189 15194 53255 15197
rect 56869 15194 56935 15197
rect 53189 15192 56935 15194
rect 53189 15136 53194 15192
rect 53250 15136 56874 15192
rect 56930 15136 56935 15192
rect 53189 15134 56935 15136
rect 53189 15131 53255 15134
rect 56869 15131 56935 15134
rect 59905 15194 59971 15197
rect 62297 15194 62363 15197
rect 64689 15194 64755 15197
rect 64965 15194 65031 15197
rect 59905 15192 65031 15194
rect 59905 15136 59910 15192
rect 59966 15136 62302 15192
rect 62358 15136 64694 15192
rect 64750 15136 64970 15192
rect 65026 15136 65031 15192
rect 59905 15134 65031 15136
rect 59905 15131 59971 15134
rect 62297 15131 62363 15134
rect 64689 15131 64755 15134
rect 64965 15131 65031 15134
rect 68645 15194 68711 15197
rect 70853 15194 70919 15197
rect 68645 15192 70919 15194
rect 68645 15136 68650 15192
rect 68706 15136 70858 15192
rect 70914 15136 70919 15192
rect 68645 15134 70919 15136
rect 68645 15131 68711 15134
rect 70853 15131 70919 15134
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 1577 15058 1643 15061
rect 62389 15058 62455 15061
rect 1577 15056 62455 15058
rect 1577 15000 1582 15056
rect 1638 15000 62394 15056
rect 62450 15000 62455 15056
rect 1577 14998 62455 15000
rect 1577 14995 1643 14998
rect 62389 14995 62455 14998
rect 62573 15058 62639 15061
rect 63585 15058 63651 15061
rect 65701 15058 65767 15061
rect 62573 15056 65767 15058
rect 62573 15000 62578 15056
rect 62634 15000 63590 15056
rect 63646 15000 65706 15056
rect 65762 15000 65767 15056
rect 62573 14998 65767 15000
rect 62573 14995 62639 14998
rect 63585 14995 63651 14998
rect 65701 14995 65767 14998
rect 88057 15058 88123 15061
rect 89200 15058 90000 15088
rect 88057 15056 90000 15058
rect 88057 15000 88062 15056
rect 88118 15000 90000 15056
rect 88057 14998 90000 15000
rect 88057 14995 88123 14998
rect 89200 14968 90000 14998
rect 22001 14922 22067 14925
rect 28533 14922 28599 14925
rect 22001 14920 28599 14922
rect 22001 14864 22006 14920
rect 22062 14864 28538 14920
rect 28594 14864 28599 14920
rect 22001 14862 28599 14864
rect 22001 14859 22067 14862
rect 28533 14859 28599 14862
rect 30281 14922 30347 14925
rect 33317 14922 33383 14925
rect 30281 14920 33383 14922
rect 30281 14864 30286 14920
rect 30342 14864 33322 14920
rect 33378 14864 33383 14920
rect 30281 14862 33383 14864
rect 30281 14859 30347 14862
rect 33317 14859 33383 14862
rect 33961 14922 34027 14925
rect 36261 14922 36327 14925
rect 37365 14922 37431 14925
rect 33961 14920 34530 14922
rect 33961 14864 33966 14920
rect 34022 14864 34530 14920
rect 33961 14862 34530 14864
rect 33961 14859 34027 14862
rect 23105 14786 23171 14789
rect 28533 14786 28599 14789
rect 23105 14784 28599 14786
rect 23105 14728 23110 14784
rect 23166 14728 28538 14784
rect 28594 14728 28599 14784
rect 23105 14726 28599 14728
rect 23105 14723 23171 14726
rect 28533 14723 28599 14726
rect 32397 14786 32463 14789
rect 33501 14786 33567 14789
rect 32397 14784 33567 14786
rect 32397 14728 32402 14784
rect 32458 14728 33506 14784
rect 33562 14728 33567 14784
rect 32397 14726 33567 14728
rect 32397 14723 32463 14726
rect 33501 14723 33567 14726
rect 11920 14720 12236 14721
rect 11920 14656 11926 14720
rect 11990 14656 12006 14720
rect 12070 14656 12086 14720
rect 12150 14656 12166 14720
rect 12230 14656 12236 14720
rect 11920 14655 12236 14656
rect 33868 14720 34184 14721
rect 33868 14656 33874 14720
rect 33938 14656 33954 14720
rect 34018 14656 34034 14720
rect 34098 14656 34114 14720
rect 34178 14656 34184 14720
rect 33868 14655 34184 14656
rect 24117 14650 24183 14653
rect 28165 14650 28231 14653
rect 24117 14648 28231 14650
rect 24117 14592 24122 14648
rect 24178 14592 28170 14648
rect 28226 14592 28231 14648
rect 24117 14590 28231 14592
rect 34470 14650 34530 14862
rect 36261 14920 37431 14922
rect 36261 14864 36266 14920
rect 36322 14864 37370 14920
rect 37426 14864 37431 14920
rect 36261 14862 37431 14864
rect 36261 14859 36327 14862
rect 37365 14859 37431 14862
rect 37917 14922 37983 14925
rect 42793 14922 42859 14925
rect 46933 14922 46999 14925
rect 37917 14920 42626 14922
rect 37917 14864 37922 14920
rect 37978 14864 42626 14920
rect 37917 14862 42626 14864
rect 37917 14859 37983 14862
rect 41597 14650 41663 14653
rect 34470 14648 41663 14650
rect 34470 14592 41602 14648
rect 41658 14592 41663 14648
rect 34470 14590 41663 14592
rect 42566 14650 42626 14862
rect 42793 14920 46999 14922
rect 42793 14864 42798 14920
rect 42854 14864 46938 14920
rect 46994 14864 46999 14920
rect 42793 14862 46999 14864
rect 42793 14859 42859 14862
rect 46933 14859 46999 14862
rect 48865 14922 48931 14925
rect 52269 14922 52335 14925
rect 48865 14920 52335 14922
rect 48865 14864 48870 14920
rect 48926 14864 52274 14920
rect 52330 14864 52335 14920
rect 48865 14862 52335 14864
rect 48865 14859 48931 14862
rect 52269 14859 52335 14862
rect 53097 14922 53163 14925
rect 54293 14922 54359 14925
rect 53097 14920 54359 14922
rect 53097 14864 53102 14920
rect 53158 14864 54298 14920
rect 54354 14864 54359 14920
rect 53097 14862 54359 14864
rect 53097 14859 53163 14862
rect 54293 14859 54359 14862
rect 56961 14922 57027 14925
rect 60825 14922 60891 14925
rect 56961 14920 60891 14922
rect 56961 14864 56966 14920
rect 57022 14864 60830 14920
rect 60886 14864 60891 14920
rect 56961 14862 60891 14864
rect 56961 14859 57027 14862
rect 60825 14859 60891 14862
rect 62941 14922 63007 14925
rect 65241 14922 65307 14925
rect 62941 14920 65307 14922
rect 62941 14864 62946 14920
rect 63002 14864 65246 14920
rect 65302 14864 65307 14920
rect 62941 14862 65307 14864
rect 62941 14859 63007 14862
rect 65241 14859 65307 14862
rect 42885 14786 42951 14789
rect 46657 14786 46723 14789
rect 42885 14784 46723 14786
rect 42885 14728 42890 14784
rect 42946 14728 46662 14784
rect 46718 14728 46723 14784
rect 42885 14726 46723 14728
rect 42885 14723 42951 14726
rect 46657 14723 46723 14726
rect 48405 14786 48471 14789
rect 54201 14786 54267 14789
rect 56869 14788 56935 14789
rect 56869 14786 56916 14788
rect 48405 14784 54267 14786
rect 48405 14728 48410 14784
rect 48466 14728 54206 14784
rect 54262 14728 54267 14784
rect 48405 14726 54267 14728
rect 56824 14784 56916 14786
rect 56824 14728 56874 14784
rect 56824 14726 56916 14728
rect 48405 14723 48471 14726
rect 54201 14723 54267 14726
rect 56869 14724 56916 14726
rect 56980 14724 56986 14788
rect 59997 14786 60063 14789
rect 66713 14786 66779 14789
rect 59997 14784 66779 14786
rect 59997 14728 60002 14784
rect 60058 14728 66718 14784
rect 66774 14728 66779 14784
rect 59997 14726 66779 14728
rect 56869 14723 56935 14724
rect 59997 14723 60063 14726
rect 66713 14723 66779 14726
rect 55816 14720 56132 14721
rect 55816 14656 55822 14720
rect 55886 14656 55902 14720
rect 55966 14656 55982 14720
rect 56046 14656 56062 14720
rect 56126 14656 56132 14720
rect 55816 14655 56132 14656
rect 77764 14720 78080 14721
rect 77764 14656 77770 14720
rect 77834 14656 77850 14720
rect 77914 14656 77930 14720
rect 77994 14656 78010 14720
rect 78074 14656 78080 14720
rect 77764 14655 78080 14656
rect 43897 14650 43963 14653
rect 50613 14650 50679 14653
rect 42566 14648 50679 14650
rect 42566 14592 43902 14648
rect 43958 14592 50618 14648
rect 50674 14592 50679 14648
rect 42566 14590 50679 14592
rect 24117 14587 24183 14590
rect 28165 14587 28231 14590
rect 41597 14587 41663 14590
rect 43897 14587 43963 14590
rect 50613 14587 50679 14590
rect 50889 14650 50955 14653
rect 51349 14650 51415 14653
rect 50889 14648 51415 14650
rect 50889 14592 50894 14648
rect 50950 14592 51354 14648
rect 51410 14592 51415 14648
rect 50889 14590 51415 14592
rect 50889 14587 50955 14590
rect 51349 14587 51415 14590
rect 51533 14650 51599 14653
rect 57973 14650 58039 14653
rect 69933 14650 69999 14653
rect 51533 14648 54586 14650
rect 51533 14592 51538 14648
rect 51594 14592 54586 14648
rect 51533 14590 54586 14592
rect 51533 14587 51599 14590
rect 22829 14514 22895 14517
rect 25589 14514 25655 14517
rect 27061 14514 27127 14517
rect 22829 14512 25376 14514
rect 22829 14456 22834 14512
rect 22890 14456 25376 14512
rect 22829 14454 25376 14456
rect 22829 14451 22895 14454
rect 0 14378 800 14408
rect 1577 14378 1643 14381
rect 0 14376 1643 14378
rect 0 14320 1582 14376
rect 1638 14320 1643 14376
rect 0 14318 1643 14320
rect 0 14288 800 14318
rect 1577 14315 1643 14318
rect 21909 14378 21975 14381
rect 23289 14378 23355 14381
rect 21909 14376 23355 14378
rect 21909 14320 21914 14376
rect 21970 14320 23294 14376
rect 23350 14320 23355 14376
rect 21909 14318 23355 14320
rect 25316 14378 25376 14454
rect 25589 14512 27127 14514
rect 25589 14456 25594 14512
rect 25650 14456 27066 14512
rect 27122 14456 27127 14512
rect 25589 14454 27127 14456
rect 25589 14451 25655 14454
rect 27061 14451 27127 14454
rect 31845 14514 31911 14517
rect 34237 14514 34303 14517
rect 39941 14514 40007 14517
rect 31845 14512 40007 14514
rect 31845 14456 31850 14512
rect 31906 14456 34242 14512
rect 34298 14456 39946 14512
rect 40002 14456 40007 14512
rect 31845 14454 40007 14456
rect 31845 14451 31911 14454
rect 34237 14451 34303 14454
rect 39941 14451 40007 14454
rect 41781 14514 41847 14517
rect 47669 14514 47735 14517
rect 51625 14514 51691 14517
rect 41781 14512 51691 14514
rect 41781 14456 41786 14512
rect 41842 14456 47674 14512
rect 47730 14456 51630 14512
rect 51686 14456 51691 14512
rect 41781 14454 51691 14456
rect 41781 14451 41847 14454
rect 47669 14451 47735 14454
rect 51625 14451 51691 14454
rect 52821 14514 52887 14517
rect 54385 14514 54451 14517
rect 52821 14512 54451 14514
rect 52821 14456 52826 14512
rect 52882 14456 54390 14512
rect 54446 14456 54451 14512
rect 52821 14454 54451 14456
rect 54526 14514 54586 14590
rect 57973 14648 69999 14650
rect 57973 14592 57978 14648
rect 58034 14592 69938 14648
rect 69994 14592 69999 14648
rect 57973 14590 69999 14592
rect 57973 14587 58039 14590
rect 69933 14587 69999 14590
rect 57605 14514 57671 14517
rect 58525 14514 58591 14517
rect 54526 14512 58591 14514
rect 54526 14456 57610 14512
rect 57666 14456 58530 14512
rect 58586 14456 58591 14512
rect 54526 14454 58591 14456
rect 52821 14451 52887 14454
rect 54385 14451 54451 14454
rect 57605 14451 57671 14454
rect 58525 14451 58591 14454
rect 62113 14514 62179 14517
rect 63217 14514 63283 14517
rect 62113 14512 63283 14514
rect 62113 14456 62118 14512
rect 62174 14456 63222 14512
rect 63278 14456 63283 14512
rect 62113 14454 63283 14456
rect 62113 14451 62179 14454
rect 63217 14451 63283 14454
rect 68645 14514 68711 14517
rect 70393 14514 70459 14517
rect 68645 14512 70459 14514
rect 68645 14456 68650 14512
rect 68706 14456 70398 14512
rect 70454 14456 70459 14512
rect 68645 14454 70459 14456
rect 68645 14451 68711 14454
rect 70393 14451 70459 14454
rect 25865 14378 25931 14381
rect 25316 14376 25931 14378
rect 25316 14320 25870 14376
rect 25926 14320 25931 14376
rect 25316 14318 25931 14320
rect 21909 14315 21975 14318
rect 23289 14315 23355 14318
rect 25865 14315 25931 14318
rect 26141 14378 26207 14381
rect 26693 14378 26759 14381
rect 26141 14376 26759 14378
rect 26141 14320 26146 14376
rect 26202 14320 26698 14376
rect 26754 14320 26759 14376
rect 26141 14318 26759 14320
rect 26141 14315 26207 14318
rect 26693 14315 26759 14318
rect 34973 14378 35039 14381
rect 36629 14378 36695 14381
rect 38285 14378 38351 14381
rect 46473 14378 46539 14381
rect 34973 14376 36695 14378
rect 34973 14320 34978 14376
rect 35034 14320 36634 14376
rect 36690 14320 36695 14376
rect 34973 14318 36695 14320
rect 34973 14315 35039 14318
rect 36629 14315 36695 14318
rect 36862 14376 46539 14378
rect 36862 14320 38290 14376
rect 38346 14320 46478 14376
rect 46534 14320 46539 14376
rect 36862 14318 46539 14320
rect 23933 14242 23999 14245
rect 28809 14242 28875 14245
rect 23933 14240 28875 14242
rect 23933 14184 23938 14240
rect 23994 14184 28814 14240
rect 28870 14184 28875 14240
rect 23933 14182 28875 14184
rect 23933 14179 23999 14182
rect 28809 14179 28875 14182
rect 30833 14242 30899 14245
rect 33317 14242 33383 14245
rect 36862 14242 36922 14318
rect 38285 14315 38351 14318
rect 46473 14315 46539 14318
rect 50429 14378 50495 14381
rect 52177 14378 52243 14381
rect 50429 14376 52243 14378
rect 50429 14320 50434 14376
rect 50490 14320 52182 14376
rect 52238 14320 52243 14376
rect 50429 14318 52243 14320
rect 50429 14315 50495 14318
rect 52177 14315 52243 14318
rect 52453 14378 52519 14381
rect 57789 14378 57855 14381
rect 52453 14376 57855 14378
rect 52453 14320 52458 14376
rect 52514 14320 57794 14376
rect 57850 14320 57855 14376
rect 52453 14318 57855 14320
rect 52453 14315 52519 14318
rect 57789 14315 57855 14318
rect 63902 14316 63908 14380
rect 63972 14378 63978 14380
rect 64045 14378 64111 14381
rect 67449 14378 67515 14381
rect 63972 14376 67515 14378
rect 63972 14320 64050 14376
rect 64106 14320 67454 14376
rect 67510 14320 67515 14376
rect 63972 14318 67515 14320
rect 63972 14316 63978 14318
rect 64045 14315 64111 14318
rect 67449 14315 67515 14318
rect 67817 14378 67883 14381
rect 69197 14378 69263 14381
rect 67817 14376 69263 14378
rect 67817 14320 67822 14376
rect 67878 14320 69202 14376
rect 69258 14320 69263 14376
rect 67817 14318 69263 14320
rect 67817 14315 67883 14318
rect 69197 14315 69263 14318
rect 88057 14378 88123 14381
rect 89200 14378 90000 14408
rect 88057 14376 90000 14378
rect 88057 14320 88062 14376
rect 88118 14320 90000 14376
rect 88057 14318 90000 14320
rect 88057 14315 88123 14318
rect 89200 14288 90000 14318
rect 30833 14240 36922 14242
rect 30833 14184 30838 14240
rect 30894 14184 33322 14240
rect 33378 14184 36922 14240
rect 30833 14182 36922 14184
rect 36997 14242 37063 14245
rect 37365 14242 37431 14245
rect 41413 14242 41479 14245
rect 44541 14242 44607 14245
rect 36997 14240 40970 14242
rect 36997 14184 37002 14240
rect 37058 14184 37370 14240
rect 37426 14184 40970 14240
rect 36997 14182 40970 14184
rect 30833 14179 30899 14182
rect 33317 14179 33383 14182
rect 36997 14179 37063 14182
rect 37365 14179 37431 14182
rect 22894 14176 23210 14177
rect 22894 14112 22900 14176
rect 22964 14112 22980 14176
rect 23044 14112 23060 14176
rect 23124 14112 23140 14176
rect 23204 14112 23210 14176
rect 22894 14111 23210 14112
rect 33869 14106 33935 14109
rect 35249 14106 35315 14109
rect 35801 14106 35867 14109
rect 37273 14106 37339 14109
rect 33869 14104 37339 14106
rect 33869 14048 33874 14104
rect 33930 14048 35254 14104
rect 35310 14048 35806 14104
rect 35862 14048 37278 14104
rect 37334 14048 37339 14104
rect 33869 14046 37339 14048
rect 40910 14106 40970 14182
rect 41413 14240 44607 14242
rect 41413 14184 41418 14240
rect 41474 14184 44546 14240
rect 44602 14184 44607 14240
rect 41413 14182 44607 14184
rect 41413 14179 41479 14182
rect 44541 14179 44607 14182
rect 47485 14242 47551 14245
rect 50613 14242 50679 14245
rect 47485 14240 50679 14242
rect 47485 14184 47490 14240
rect 47546 14184 50618 14240
rect 50674 14184 50679 14240
rect 47485 14182 50679 14184
rect 47485 14179 47551 14182
rect 50613 14179 50679 14182
rect 50797 14242 50863 14245
rect 54937 14242 55003 14245
rect 50797 14240 55003 14242
rect 50797 14184 50802 14240
rect 50858 14184 54942 14240
rect 54998 14184 55003 14240
rect 50797 14182 55003 14184
rect 50797 14179 50863 14182
rect 54937 14179 55003 14182
rect 55121 14242 55187 14245
rect 60273 14242 60339 14245
rect 55121 14240 60339 14242
rect 55121 14184 55126 14240
rect 55182 14184 60278 14240
rect 60334 14184 60339 14240
rect 55121 14182 60339 14184
rect 55121 14179 55187 14182
rect 60273 14179 60339 14182
rect 60549 14242 60615 14245
rect 64413 14242 64479 14245
rect 60549 14240 64479 14242
rect 60549 14184 60554 14240
rect 60610 14184 64418 14240
rect 64474 14184 64479 14240
rect 60549 14182 64479 14184
rect 60549 14179 60615 14182
rect 64413 14179 64479 14182
rect 67449 14242 67515 14245
rect 69105 14242 69171 14245
rect 67449 14240 69171 14242
rect 67449 14184 67454 14240
rect 67510 14184 69110 14240
rect 69166 14184 69171 14240
rect 67449 14182 69171 14184
rect 67449 14179 67515 14182
rect 69105 14179 69171 14182
rect 44842 14176 45158 14177
rect 44842 14112 44848 14176
rect 44912 14112 44928 14176
rect 44992 14112 45008 14176
rect 45072 14112 45088 14176
rect 45152 14112 45158 14176
rect 44842 14111 45158 14112
rect 66790 14176 67106 14177
rect 66790 14112 66796 14176
rect 66860 14112 66876 14176
rect 66940 14112 66956 14176
rect 67020 14112 67036 14176
rect 67100 14112 67106 14176
rect 66790 14111 67106 14112
rect 41505 14106 41571 14109
rect 40910 14104 41571 14106
rect 40910 14048 41510 14104
rect 41566 14048 41571 14104
rect 40910 14046 41571 14048
rect 33869 14043 33935 14046
rect 35249 14043 35315 14046
rect 35801 14043 35867 14046
rect 37273 14043 37339 14046
rect 41505 14043 41571 14046
rect 45277 14106 45343 14109
rect 50337 14106 50403 14109
rect 45277 14104 50403 14106
rect 45277 14048 45282 14104
rect 45338 14048 50342 14104
rect 50398 14048 50403 14104
rect 45277 14046 50403 14048
rect 45277 14043 45343 14046
rect 50337 14043 50403 14046
rect 52269 14106 52335 14109
rect 57053 14106 57119 14109
rect 52269 14104 57119 14106
rect 52269 14048 52274 14104
rect 52330 14048 57058 14104
rect 57114 14048 57119 14104
rect 52269 14046 57119 14048
rect 52269 14043 52335 14046
rect 57053 14043 57119 14046
rect 57237 14106 57303 14109
rect 61561 14106 61627 14109
rect 57237 14104 61627 14106
rect 57237 14048 57242 14104
rect 57298 14048 61566 14104
rect 61622 14048 61627 14104
rect 57237 14046 61627 14048
rect 57237 14043 57303 14046
rect 61561 14043 61627 14046
rect 61837 14106 61903 14109
rect 63033 14106 63099 14109
rect 61837 14104 63099 14106
rect 61837 14048 61842 14104
rect 61898 14048 63038 14104
rect 63094 14048 63099 14104
rect 61837 14046 63099 14048
rect 61837 14043 61903 14046
rect 63033 14043 63099 14046
rect 64045 14106 64111 14109
rect 65793 14106 65859 14109
rect 64045 14104 65859 14106
rect 64045 14048 64050 14104
rect 64106 14048 65798 14104
rect 65854 14048 65859 14104
rect 64045 14046 65859 14048
rect 64045 14043 64111 14046
rect 65793 14043 65859 14046
rect 67725 14106 67791 14109
rect 68921 14106 68987 14109
rect 67725 14104 68987 14106
rect 67725 14048 67730 14104
rect 67786 14048 68926 14104
rect 68982 14048 68987 14104
rect 67725 14046 68987 14048
rect 67725 14043 67791 14046
rect 68921 14043 68987 14046
rect 22093 13970 22159 13973
rect 22829 13970 22895 13973
rect 27797 13970 27863 13973
rect 22093 13968 27863 13970
rect 22093 13912 22098 13968
rect 22154 13912 22834 13968
rect 22890 13912 27802 13968
rect 27858 13912 27863 13968
rect 22093 13910 27863 13912
rect 22093 13907 22159 13910
rect 22829 13907 22895 13910
rect 27797 13907 27863 13910
rect 28073 13970 28139 13973
rect 87965 13970 88031 13973
rect 28073 13968 88031 13970
rect 28073 13912 28078 13968
rect 28134 13912 87970 13968
rect 88026 13912 88031 13968
rect 28073 13910 88031 13912
rect 28073 13907 28139 13910
rect 87965 13907 88031 13910
rect 22093 13834 22159 13837
rect 30925 13834 30991 13837
rect 22093 13832 30991 13834
rect 22093 13776 22098 13832
rect 22154 13776 30930 13832
rect 30986 13776 30991 13832
rect 22093 13774 30991 13776
rect 22093 13771 22159 13774
rect 30925 13771 30991 13774
rect 31109 13834 31175 13837
rect 33409 13834 33475 13837
rect 36997 13834 37063 13837
rect 31109 13832 33475 13834
rect 31109 13776 31114 13832
rect 31170 13776 33414 13832
rect 33470 13776 33475 13832
rect 31109 13774 33475 13776
rect 31109 13771 31175 13774
rect 33409 13771 33475 13774
rect 33734 13832 37063 13834
rect 33734 13776 37002 13832
rect 37058 13776 37063 13832
rect 33734 13774 37063 13776
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 19885 13698 19951 13701
rect 26785 13698 26851 13701
rect 19885 13696 26851 13698
rect 19885 13640 19890 13696
rect 19946 13640 26790 13696
rect 26846 13640 26851 13696
rect 19885 13638 26851 13640
rect 19885 13635 19951 13638
rect 26785 13635 26851 13638
rect 32857 13698 32923 13701
rect 33734 13698 33794 13774
rect 36997 13771 37063 13774
rect 37549 13834 37615 13837
rect 40125 13834 40191 13837
rect 37549 13832 40191 13834
rect 37549 13776 37554 13832
rect 37610 13776 40130 13832
rect 40186 13776 40191 13832
rect 37549 13774 40191 13776
rect 37549 13771 37615 13774
rect 40125 13771 40191 13774
rect 40309 13834 40375 13837
rect 41689 13834 41755 13837
rect 47853 13834 47919 13837
rect 40309 13832 41755 13834
rect 40309 13776 40314 13832
rect 40370 13776 41694 13832
rect 41750 13776 41755 13832
rect 40309 13774 41755 13776
rect 40309 13771 40375 13774
rect 41689 13771 41755 13774
rect 41830 13832 47919 13834
rect 41830 13776 47858 13832
rect 47914 13776 47919 13832
rect 41830 13774 47919 13776
rect 32857 13696 33794 13698
rect 32857 13640 32862 13696
rect 32918 13640 33794 13696
rect 32857 13638 33794 13640
rect 34881 13698 34947 13701
rect 36445 13698 36511 13701
rect 34881 13696 36511 13698
rect 34881 13640 34886 13696
rect 34942 13640 36450 13696
rect 36506 13640 36511 13696
rect 34881 13638 36511 13640
rect 32857 13635 32923 13638
rect 34881 13635 34947 13638
rect 36445 13635 36511 13638
rect 39389 13698 39455 13701
rect 40953 13698 41019 13701
rect 39389 13696 41019 13698
rect 39389 13640 39394 13696
rect 39450 13640 40958 13696
rect 41014 13640 41019 13696
rect 39389 13638 41019 13640
rect 39389 13635 39455 13638
rect 40953 13635 41019 13638
rect 41321 13698 41387 13701
rect 41830 13698 41890 13774
rect 47853 13771 47919 13774
rect 48313 13834 48379 13837
rect 52361 13834 52427 13837
rect 48313 13832 52427 13834
rect 48313 13776 48318 13832
rect 48374 13776 52366 13832
rect 52422 13776 52427 13832
rect 48313 13774 52427 13776
rect 48313 13771 48379 13774
rect 52361 13771 52427 13774
rect 52913 13834 52979 13837
rect 56869 13834 56935 13837
rect 59997 13834 60063 13837
rect 52913 13832 60063 13834
rect 52913 13776 52918 13832
rect 52974 13776 56874 13832
rect 56930 13776 60002 13832
rect 60058 13776 60063 13832
rect 52913 13774 60063 13776
rect 52913 13771 52979 13774
rect 56869 13771 56935 13774
rect 59997 13771 60063 13774
rect 60641 13834 60707 13837
rect 60825 13834 60891 13837
rect 60641 13832 60891 13834
rect 60641 13776 60646 13832
rect 60702 13776 60830 13832
rect 60886 13776 60891 13832
rect 60641 13774 60891 13776
rect 60641 13771 60707 13774
rect 60825 13771 60891 13774
rect 61009 13834 61075 13837
rect 63493 13834 63559 13837
rect 67449 13834 67515 13837
rect 61009 13832 67515 13834
rect 61009 13776 61014 13832
rect 61070 13776 63498 13832
rect 63554 13776 67454 13832
rect 67510 13776 67515 13832
rect 61009 13774 67515 13776
rect 61009 13771 61075 13774
rect 63493 13771 63559 13774
rect 67449 13771 67515 13774
rect 41321 13696 41890 13698
rect 41321 13640 41326 13696
rect 41382 13640 41890 13696
rect 41321 13638 41890 13640
rect 43805 13698 43871 13701
rect 46013 13698 46079 13701
rect 43805 13696 46079 13698
rect 43805 13640 43810 13696
rect 43866 13640 46018 13696
rect 46074 13640 46079 13696
rect 43805 13638 46079 13640
rect 41321 13635 41387 13638
rect 43805 13635 43871 13638
rect 46013 13635 46079 13638
rect 49233 13698 49299 13701
rect 55673 13698 55739 13701
rect 49233 13696 55739 13698
rect 49233 13640 49238 13696
rect 49294 13640 55678 13696
rect 55734 13640 55739 13696
rect 49233 13638 55739 13640
rect 49233 13635 49299 13638
rect 55673 13635 55739 13638
rect 57421 13698 57487 13701
rect 61377 13698 61443 13701
rect 57421 13696 61443 13698
rect 57421 13640 57426 13696
rect 57482 13640 61382 13696
rect 61438 13640 61443 13696
rect 57421 13638 61443 13640
rect 57421 13635 57487 13638
rect 61377 13635 61443 13638
rect 62113 13698 62179 13701
rect 65149 13698 65215 13701
rect 62113 13696 65215 13698
rect 62113 13640 62118 13696
rect 62174 13640 65154 13696
rect 65210 13640 65215 13696
rect 62113 13638 65215 13640
rect 62113 13635 62179 13638
rect 65149 13635 65215 13638
rect 88057 13698 88123 13701
rect 89200 13698 90000 13728
rect 88057 13696 90000 13698
rect 88057 13640 88062 13696
rect 88118 13640 90000 13696
rect 88057 13638 90000 13640
rect 88057 13635 88123 13638
rect 11920 13632 12236 13633
rect 11920 13568 11926 13632
rect 11990 13568 12006 13632
rect 12070 13568 12086 13632
rect 12150 13568 12166 13632
rect 12230 13568 12236 13632
rect 11920 13567 12236 13568
rect 33868 13632 34184 13633
rect 33868 13568 33874 13632
rect 33938 13568 33954 13632
rect 34018 13568 34034 13632
rect 34098 13568 34114 13632
rect 34178 13568 34184 13632
rect 33868 13567 34184 13568
rect 55816 13632 56132 13633
rect 55816 13568 55822 13632
rect 55886 13568 55902 13632
rect 55966 13568 55982 13632
rect 56046 13568 56062 13632
rect 56126 13568 56132 13632
rect 55816 13567 56132 13568
rect 77764 13632 78080 13633
rect 77764 13568 77770 13632
rect 77834 13568 77850 13632
rect 77914 13568 77930 13632
rect 77994 13568 78010 13632
rect 78074 13568 78080 13632
rect 89200 13608 90000 13638
rect 77764 13567 78080 13568
rect 20069 13562 20135 13565
rect 26877 13562 26943 13565
rect 20069 13560 26943 13562
rect 20069 13504 20074 13560
rect 20130 13504 26882 13560
rect 26938 13504 26943 13560
rect 20069 13502 26943 13504
rect 20069 13499 20135 13502
rect 26877 13499 26943 13502
rect 34605 13562 34671 13565
rect 35709 13562 35775 13565
rect 34605 13560 35775 13562
rect 34605 13504 34610 13560
rect 34666 13504 35714 13560
rect 35770 13504 35775 13560
rect 34605 13502 35775 13504
rect 34605 13499 34671 13502
rect 35709 13499 35775 13502
rect 38745 13562 38811 13565
rect 39389 13562 39455 13565
rect 42885 13562 42951 13565
rect 38745 13560 42951 13562
rect 38745 13504 38750 13560
rect 38806 13504 39394 13560
rect 39450 13504 42890 13560
rect 42946 13504 42951 13560
rect 38745 13502 42951 13504
rect 38745 13499 38811 13502
rect 39389 13499 39455 13502
rect 42885 13499 42951 13502
rect 44081 13562 44147 13565
rect 44725 13562 44791 13565
rect 44081 13560 44791 13562
rect 44081 13504 44086 13560
rect 44142 13504 44730 13560
rect 44786 13504 44791 13560
rect 44081 13502 44791 13504
rect 44081 13499 44147 13502
rect 44725 13499 44791 13502
rect 45553 13562 45619 13565
rect 48221 13562 48287 13565
rect 45553 13560 48287 13562
rect 45553 13504 45558 13560
rect 45614 13504 48226 13560
rect 48282 13504 48287 13560
rect 45553 13502 48287 13504
rect 45553 13499 45619 13502
rect 48221 13499 48287 13502
rect 48865 13562 48931 13565
rect 49233 13562 49299 13565
rect 48865 13560 49299 13562
rect 48865 13504 48870 13560
rect 48926 13504 49238 13560
rect 49294 13504 49299 13560
rect 48865 13502 49299 13504
rect 48865 13499 48931 13502
rect 49233 13499 49299 13502
rect 50153 13562 50219 13565
rect 50981 13562 51047 13565
rect 50153 13560 51047 13562
rect 50153 13504 50158 13560
rect 50214 13504 50986 13560
rect 51042 13504 51047 13560
rect 50153 13502 51047 13504
rect 50153 13499 50219 13502
rect 50981 13499 51047 13502
rect 51165 13562 51231 13565
rect 55622 13562 55628 13564
rect 51165 13560 55628 13562
rect 51165 13504 51170 13560
rect 51226 13504 55628 13560
rect 51165 13502 55628 13504
rect 51165 13499 51231 13502
rect 55622 13500 55628 13502
rect 55692 13500 55698 13564
rect 57053 13562 57119 13565
rect 60273 13562 60339 13565
rect 57053 13560 60339 13562
rect 57053 13504 57058 13560
rect 57114 13504 60278 13560
rect 60334 13504 60339 13560
rect 57053 13502 60339 13504
rect 57053 13499 57119 13502
rect 60273 13499 60339 13502
rect 60549 13562 60615 13565
rect 62297 13562 62363 13565
rect 66345 13562 66411 13565
rect 60549 13560 66411 13562
rect 60549 13504 60554 13560
rect 60610 13504 62302 13560
rect 62358 13504 66350 13560
rect 66406 13504 66411 13560
rect 60549 13502 66411 13504
rect 60549 13499 60615 13502
rect 62297 13499 62363 13502
rect 66345 13499 66411 13502
rect 69381 13562 69447 13565
rect 70301 13562 70367 13565
rect 69381 13560 70367 13562
rect 69381 13504 69386 13560
rect 69442 13504 70306 13560
rect 70362 13504 70367 13560
rect 69381 13502 70367 13504
rect 69381 13499 69447 13502
rect 70301 13499 70367 13502
rect 25037 13426 25103 13429
rect 27889 13426 27955 13429
rect 79593 13426 79659 13429
rect 25037 13424 79659 13426
rect 25037 13368 25042 13424
rect 25098 13368 27894 13424
rect 27950 13368 79598 13424
rect 79654 13368 79659 13424
rect 25037 13366 79659 13368
rect 25037 13363 25103 13366
rect 27889 13363 27955 13366
rect 79593 13363 79659 13366
rect 21173 13290 21239 13293
rect 26049 13290 26115 13293
rect 21173 13288 26115 13290
rect 21173 13232 21178 13288
rect 21234 13232 26054 13288
rect 26110 13232 26115 13288
rect 21173 13230 26115 13232
rect 21173 13227 21239 13230
rect 26049 13227 26115 13230
rect 29637 13290 29703 13293
rect 51165 13290 51231 13293
rect 29637 13288 51231 13290
rect 29637 13232 29642 13288
rect 29698 13232 51170 13288
rect 51226 13232 51231 13288
rect 29637 13230 51231 13232
rect 29637 13227 29703 13230
rect 51165 13227 51231 13230
rect 51533 13290 51599 13293
rect 58065 13290 58131 13293
rect 58341 13290 58407 13293
rect 51533 13288 58407 13290
rect 51533 13232 51538 13288
rect 51594 13232 58070 13288
rect 58126 13232 58346 13288
rect 58402 13232 58407 13288
rect 51533 13230 58407 13232
rect 51533 13227 51599 13230
rect 58065 13227 58131 13230
rect 58341 13227 58407 13230
rect 59445 13290 59511 13293
rect 60549 13290 60615 13293
rect 59445 13288 60615 13290
rect 59445 13232 59450 13288
rect 59506 13232 60554 13288
rect 60610 13232 60615 13288
rect 59445 13230 60615 13232
rect 59445 13227 59511 13230
rect 60549 13227 60615 13230
rect 60733 13290 60799 13293
rect 64505 13290 64571 13293
rect 60733 13288 64571 13290
rect 60733 13232 60738 13288
rect 60794 13232 64510 13288
rect 64566 13232 64571 13288
rect 60733 13230 64571 13232
rect 60733 13227 60799 13230
rect 64505 13227 64571 13230
rect 23933 13154 23999 13157
rect 26325 13154 26391 13157
rect 23933 13152 26391 13154
rect 23933 13096 23938 13152
rect 23994 13096 26330 13152
rect 26386 13096 26391 13152
rect 23933 13094 26391 13096
rect 23933 13091 23999 13094
rect 26325 13091 26391 13094
rect 34145 13154 34211 13157
rect 36905 13154 36971 13157
rect 34145 13152 36971 13154
rect 34145 13096 34150 13152
rect 34206 13096 36910 13152
rect 36966 13096 36971 13152
rect 34145 13094 36971 13096
rect 34145 13091 34211 13094
rect 36905 13091 36971 13094
rect 37273 13154 37339 13157
rect 40585 13154 40651 13157
rect 37273 13152 40651 13154
rect 37273 13096 37278 13152
rect 37334 13096 40590 13152
rect 40646 13096 40651 13152
rect 37273 13094 40651 13096
rect 37273 13091 37339 13094
rect 40585 13091 40651 13094
rect 40953 13154 41019 13157
rect 43897 13154 43963 13157
rect 40953 13152 43963 13154
rect 40953 13096 40958 13152
rect 41014 13096 43902 13152
rect 43958 13096 43963 13152
rect 40953 13094 43963 13096
rect 40953 13091 41019 13094
rect 43897 13091 43963 13094
rect 45829 13154 45895 13157
rect 49417 13154 49483 13157
rect 45829 13152 49483 13154
rect 45829 13096 45834 13152
rect 45890 13096 49422 13152
rect 49478 13096 49483 13152
rect 45829 13094 49483 13096
rect 45829 13091 45895 13094
rect 49417 13091 49483 13094
rect 49601 13154 49667 13157
rect 55673 13154 55739 13157
rect 60825 13154 60891 13157
rect 64045 13154 64111 13157
rect 49601 13152 55552 13154
rect 49601 13096 49606 13152
rect 49662 13096 55552 13152
rect 49601 13094 55552 13096
rect 49601 13091 49667 13094
rect 22894 13088 23210 13089
rect 0 13018 800 13048
rect 22894 13024 22900 13088
rect 22964 13024 22980 13088
rect 23044 13024 23060 13088
rect 23124 13024 23140 13088
rect 23204 13024 23210 13088
rect 22894 13023 23210 13024
rect 44842 13088 45158 13089
rect 44842 13024 44848 13088
rect 44912 13024 44928 13088
rect 44992 13024 45008 13088
rect 45072 13024 45088 13088
rect 45152 13024 45158 13088
rect 44842 13023 45158 13024
rect 1577 13018 1643 13021
rect 0 13016 1643 13018
rect 0 12960 1582 13016
rect 1638 12960 1643 13016
rect 0 12958 1643 12960
rect 0 12928 800 12958
rect 1577 12955 1643 12958
rect 24209 13018 24275 13021
rect 26141 13018 26207 13021
rect 43437 13018 43503 13021
rect 24209 13016 26207 13018
rect 24209 12960 24214 13016
rect 24270 12960 26146 13016
rect 26202 12960 26207 13016
rect 24209 12958 26207 12960
rect 24209 12955 24275 12958
rect 26141 12955 26207 12958
rect 38610 13016 43503 13018
rect 38610 12960 43442 13016
rect 43498 12960 43503 13016
rect 38610 12958 43503 12960
rect 24025 12882 24091 12885
rect 26509 12884 26575 12885
rect 26509 12882 26556 12884
rect 24025 12880 26556 12882
rect 24025 12824 24030 12880
rect 24086 12824 26514 12880
rect 24025 12822 26556 12824
rect 24025 12819 24091 12822
rect 26509 12820 26556 12822
rect 26620 12820 26626 12884
rect 35525 12882 35591 12885
rect 38610 12882 38670 12958
rect 43437 12955 43503 12958
rect 45461 13018 45527 13021
rect 46841 13018 46907 13021
rect 49509 13018 49575 13021
rect 45461 13016 49575 13018
rect 45461 12960 45466 13016
rect 45522 12960 46846 13016
rect 46902 12960 49514 13016
rect 49570 12960 49575 13016
rect 45461 12958 49575 12960
rect 45461 12955 45527 12958
rect 46841 12955 46907 12958
rect 49509 12955 49575 12958
rect 50889 13018 50955 13021
rect 52821 13018 52887 13021
rect 50889 13016 52887 13018
rect 50889 12960 50894 13016
rect 50950 12960 52826 13016
rect 52882 12960 52887 13016
rect 50889 12958 52887 12960
rect 50889 12955 50955 12958
rect 52821 12955 52887 12958
rect 53005 13018 53071 13021
rect 54109 13018 54175 13021
rect 54753 13018 54819 13021
rect 53005 13016 54819 13018
rect 53005 12960 53010 13016
rect 53066 12960 54114 13016
rect 54170 12960 54758 13016
rect 54814 12960 54819 13016
rect 53005 12958 54819 12960
rect 55492 13018 55552 13094
rect 55673 13152 60891 13154
rect 55673 13096 55678 13152
rect 55734 13096 60830 13152
rect 60886 13096 60891 13152
rect 55673 13094 60891 13096
rect 55673 13091 55739 13094
rect 60825 13091 60891 13094
rect 60966 13152 64111 13154
rect 60966 13096 64050 13152
rect 64106 13096 64111 13152
rect 60966 13094 64111 13096
rect 56041 13018 56107 13021
rect 58157 13018 58223 13021
rect 55492 13016 58223 13018
rect 55492 12960 56046 13016
rect 56102 12960 58162 13016
rect 58218 12960 58223 13016
rect 55492 12958 58223 12960
rect 53005 12955 53071 12958
rect 54109 12955 54175 12958
rect 54753 12955 54819 12958
rect 56041 12955 56107 12958
rect 58157 12955 58223 12958
rect 58341 13018 58407 13021
rect 60966 13018 61026 13094
rect 64045 13091 64111 13094
rect 67725 13154 67791 13157
rect 69473 13154 69539 13157
rect 67725 13152 69539 13154
rect 67725 13096 67730 13152
rect 67786 13096 69478 13152
rect 69534 13096 69539 13152
rect 67725 13094 69539 13096
rect 67725 13091 67791 13094
rect 69473 13091 69539 13094
rect 69841 13154 69907 13157
rect 70761 13154 70827 13157
rect 69841 13152 70827 13154
rect 69841 13096 69846 13152
rect 69902 13096 70766 13152
rect 70822 13096 70827 13152
rect 69841 13094 70827 13096
rect 69841 13091 69907 13094
rect 70761 13091 70827 13094
rect 66790 13088 67106 13089
rect 66790 13024 66796 13088
rect 66860 13024 66876 13088
rect 66940 13024 66956 13088
rect 67020 13024 67036 13088
rect 67100 13024 67106 13088
rect 66790 13023 67106 13024
rect 58341 13016 61026 13018
rect 58341 12960 58346 13016
rect 58402 12960 61026 13016
rect 58341 12958 61026 12960
rect 63217 13018 63283 13021
rect 66621 13018 66687 13021
rect 63217 13016 66687 13018
rect 63217 12960 63222 13016
rect 63278 12960 66626 13016
rect 66682 12960 66687 13016
rect 63217 12958 66687 12960
rect 58341 12955 58407 12958
rect 63217 12955 63283 12958
rect 66621 12955 66687 12958
rect 69289 13018 69355 13021
rect 71681 13018 71747 13021
rect 69289 13016 71747 13018
rect 69289 12960 69294 13016
rect 69350 12960 71686 13016
rect 71742 12960 71747 13016
rect 69289 12958 71747 12960
rect 69289 12955 69355 12958
rect 71681 12955 71747 12958
rect 88057 13018 88123 13021
rect 89200 13018 90000 13048
rect 88057 13016 90000 13018
rect 88057 12960 88062 13016
rect 88118 12960 90000 13016
rect 88057 12958 90000 12960
rect 88057 12955 88123 12958
rect 89200 12928 90000 12958
rect 35525 12880 38670 12882
rect 35525 12824 35530 12880
rect 35586 12824 38670 12880
rect 35525 12822 38670 12824
rect 41781 12882 41847 12885
rect 42793 12882 42859 12885
rect 41781 12880 42859 12882
rect 41781 12824 41786 12880
rect 41842 12824 42798 12880
rect 42854 12824 42859 12880
rect 41781 12822 42859 12824
rect 26509 12819 26575 12820
rect 35525 12819 35591 12822
rect 41781 12819 41847 12822
rect 42793 12819 42859 12822
rect 45277 12882 45343 12885
rect 48405 12882 48471 12885
rect 87781 12882 87847 12885
rect 45277 12880 48471 12882
rect 45277 12824 45282 12880
rect 45338 12824 48410 12880
rect 48466 12824 48471 12880
rect 45277 12822 48471 12824
rect 45277 12819 45343 12822
rect 48405 12819 48471 12822
rect 48638 12880 87847 12882
rect 48638 12824 87786 12880
rect 87842 12824 87847 12880
rect 48638 12822 87847 12824
rect 26049 12746 26115 12749
rect 41505 12746 41571 12749
rect 45921 12746 45987 12749
rect 26049 12744 38670 12746
rect 26049 12688 26054 12744
rect 26110 12688 38670 12744
rect 26049 12686 38670 12688
rect 26049 12683 26115 12686
rect 19977 12610 20043 12613
rect 26325 12610 26391 12613
rect 26969 12610 27035 12613
rect 19977 12608 27035 12610
rect 19977 12552 19982 12608
rect 20038 12552 26330 12608
rect 26386 12552 26974 12608
rect 27030 12552 27035 12608
rect 19977 12550 27035 12552
rect 38610 12610 38670 12686
rect 41505 12744 45987 12746
rect 41505 12688 41510 12744
rect 41566 12688 45926 12744
rect 45982 12688 45987 12744
rect 41505 12686 45987 12688
rect 41505 12683 41571 12686
rect 45921 12683 45987 12686
rect 46105 12746 46171 12749
rect 48638 12746 48698 12822
rect 87781 12819 87847 12822
rect 46105 12744 48698 12746
rect 46105 12688 46110 12744
rect 46166 12688 48698 12744
rect 46105 12686 48698 12688
rect 50153 12746 50219 12749
rect 53281 12746 53347 12749
rect 86953 12746 87019 12749
rect 50153 12744 53347 12746
rect 50153 12688 50158 12744
rect 50214 12688 53286 12744
rect 53342 12688 53347 12744
rect 50153 12686 53347 12688
rect 46105 12683 46171 12686
rect 50153 12683 50219 12686
rect 53281 12683 53347 12686
rect 55492 12744 87019 12746
rect 55492 12688 86958 12744
rect 87014 12688 87019 12744
rect 55492 12686 87019 12688
rect 46565 12610 46631 12613
rect 38610 12608 46631 12610
rect 38610 12552 46570 12608
rect 46626 12552 46631 12608
rect 38610 12550 46631 12552
rect 19977 12547 20043 12550
rect 26325 12547 26391 12550
rect 26969 12547 27035 12550
rect 46565 12547 46631 12550
rect 47117 12610 47183 12613
rect 55492 12610 55552 12686
rect 86953 12683 87019 12686
rect 47117 12608 55552 12610
rect 47117 12552 47122 12608
rect 47178 12552 55552 12608
rect 47117 12550 55552 12552
rect 56593 12610 56659 12613
rect 62757 12610 62823 12613
rect 56593 12608 62823 12610
rect 56593 12552 56598 12608
rect 56654 12552 62762 12608
rect 62818 12552 62823 12608
rect 56593 12550 62823 12552
rect 47117 12547 47183 12550
rect 56593 12547 56659 12550
rect 62757 12547 62823 12550
rect 63033 12610 63099 12613
rect 63585 12610 63651 12613
rect 63033 12608 63651 12610
rect 63033 12552 63038 12608
rect 63094 12552 63590 12608
rect 63646 12552 63651 12608
rect 63033 12550 63651 12552
rect 63033 12547 63099 12550
rect 63585 12547 63651 12550
rect 63769 12610 63835 12613
rect 64270 12610 64276 12612
rect 63769 12608 64276 12610
rect 63769 12552 63774 12608
rect 63830 12552 64276 12608
rect 63769 12550 64276 12552
rect 63769 12547 63835 12550
rect 64270 12548 64276 12550
rect 64340 12548 64346 12612
rect 68829 12610 68895 12613
rect 72417 12610 72483 12613
rect 68829 12608 72483 12610
rect 68829 12552 68834 12608
rect 68890 12552 72422 12608
rect 72478 12552 72483 12608
rect 68829 12550 72483 12552
rect 68829 12547 68895 12550
rect 72417 12547 72483 12550
rect 11920 12544 12236 12545
rect 11920 12480 11926 12544
rect 11990 12480 12006 12544
rect 12070 12480 12086 12544
rect 12150 12480 12166 12544
rect 12230 12480 12236 12544
rect 11920 12479 12236 12480
rect 33868 12544 34184 12545
rect 33868 12480 33874 12544
rect 33938 12480 33954 12544
rect 34018 12480 34034 12544
rect 34098 12480 34114 12544
rect 34178 12480 34184 12544
rect 33868 12479 34184 12480
rect 55816 12544 56132 12545
rect 55816 12480 55822 12544
rect 55886 12480 55902 12544
rect 55966 12480 55982 12544
rect 56046 12480 56062 12544
rect 56126 12480 56132 12544
rect 55816 12479 56132 12480
rect 77764 12544 78080 12545
rect 77764 12480 77770 12544
rect 77834 12480 77850 12544
rect 77914 12480 77930 12544
rect 77994 12480 78010 12544
rect 78074 12480 78080 12544
rect 77764 12479 78080 12480
rect 24669 12474 24735 12477
rect 28349 12474 28415 12477
rect 24669 12472 28415 12474
rect 24669 12416 24674 12472
rect 24730 12416 28354 12472
rect 28410 12416 28415 12472
rect 24669 12414 28415 12416
rect 24669 12411 24735 12414
rect 28349 12411 28415 12414
rect 48129 12474 48195 12477
rect 48405 12474 48471 12477
rect 48129 12472 48471 12474
rect 48129 12416 48134 12472
rect 48190 12416 48410 12472
rect 48466 12416 48471 12472
rect 48129 12414 48471 12416
rect 48129 12411 48195 12414
rect 48405 12411 48471 12414
rect 48681 12474 48747 12477
rect 53005 12474 53071 12477
rect 48681 12472 53071 12474
rect 48681 12416 48686 12472
rect 48742 12416 53010 12472
rect 53066 12416 53071 12472
rect 48681 12414 53071 12416
rect 48681 12411 48747 12414
rect 53005 12411 53071 12414
rect 53373 12474 53439 12477
rect 58709 12474 58775 12477
rect 60365 12474 60431 12477
rect 62665 12474 62731 12477
rect 53373 12472 53988 12474
rect 53373 12416 53378 12472
rect 53434 12416 53988 12472
rect 53373 12414 53988 12416
rect 53373 12411 53439 12414
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 25129 12338 25195 12341
rect 27981 12338 28047 12341
rect 25129 12336 28047 12338
rect 25129 12280 25134 12336
rect 25190 12280 27986 12336
rect 28042 12280 28047 12336
rect 25129 12278 28047 12280
rect 25129 12275 25195 12278
rect 27981 12275 28047 12278
rect 28257 12338 28323 12341
rect 28809 12338 28875 12341
rect 28257 12336 28875 12338
rect 28257 12280 28262 12336
rect 28318 12280 28814 12336
rect 28870 12280 28875 12336
rect 28257 12278 28875 12280
rect 28257 12275 28323 12278
rect 28809 12275 28875 12278
rect 33225 12338 33291 12341
rect 38561 12338 38627 12341
rect 33225 12336 38627 12338
rect 33225 12280 33230 12336
rect 33286 12280 38566 12336
rect 38622 12280 38627 12336
rect 33225 12278 38627 12280
rect 33225 12275 33291 12278
rect 38561 12275 38627 12278
rect 38837 12338 38903 12341
rect 43621 12338 43687 12341
rect 49969 12338 50035 12341
rect 38837 12336 41890 12338
rect 38837 12280 38842 12336
rect 38898 12280 41890 12336
rect 38837 12278 41890 12280
rect 38837 12275 38903 12278
rect 25221 12202 25287 12205
rect 30005 12202 30071 12205
rect 25221 12200 30071 12202
rect 25221 12144 25226 12200
rect 25282 12144 30010 12200
rect 30066 12144 30071 12200
rect 25221 12142 30071 12144
rect 25221 12139 25287 12142
rect 30005 12139 30071 12142
rect 35433 12202 35499 12205
rect 37181 12202 37247 12205
rect 35433 12200 37247 12202
rect 35433 12144 35438 12200
rect 35494 12144 37186 12200
rect 37242 12144 37247 12200
rect 35433 12142 37247 12144
rect 35433 12139 35499 12142
rect 37181 12139 37247 12142
rect 40033 12202 40099 12205
rect 41689 12202 41755 12205
rect 40033 12200 41755 12202
rect 40033 12144 40038 12200
rect 40094 12144 41694 12200
rect 41750 12144 41755 12200
rect 40033 12142 41755 12144
rect 41830 12202 41890 12278
rect 43621 12336 50035 12338
rect 43621 12280 43626 12336
rect 43682 12280 49974 12336
rect 50030 12280 50035 12336
rect 43621 12278 50035 12280
rect 43621 12275 43687 12278
rect 49969 12275 50035 12278
rect 50429 12338 50495 12341
rect 53741 12338 53807 12341
rect 50429 12336 53807 12338
rect 50429 12280 50434 12336
rect 50490 12280 53746 12336
rect 53802 12280 53807 12336
rect 50429 12278 53807 12280
rect 53928 12338 53988 12414
rect 58709 12472 60106 12474
rect 58709 12416 58714 12472
rect 58770 12416 60106 12472
rect 58709 12414 60106 12416
rect 58709 12411 58775 12414
rect 59905 12338 59971 12341
rect 53928 12336 59971 12338
rect 53928 12280 59910 12336
rect 59966 12280 59971 12336
rect 53928 12278 59971 12280
rect 50429 12275 50495 12278
rect 53741 12275 53807 12278
rect 59905 12275 59971 12278
rect 46381 12202 46447 12205
rect 41830 12200 46447 12202
rect 41830 12144 46386 12200
rect 46442 12144 46447 12200
rect 41830 12142 46447 12144
rect 40033 12139 40099 12142
rect 41689 12139 41755 12142
rect 46381 12139 46447 12142
rect 52913 12202 52979 12205
rect 60046 12202 60106 12414
rect 60365 12472 62731 12474
rect 60365 12416 60370 12472
rect 60426 12416 62670 12472
rect 62726 12416 62731 12472
rect 60365 12414 62731 12416
rect 60365 12411 60431 12414
rect 62665 12411 62731 12414
rect 63677 12476 63743 12477
rect 63677 12472 63724 12476
rect 63788 12474 63794 12476
rect 67633 12474 67699 12477
rect 63677 12416 63682 12472
rect 63677 12412 63724 12416
rect 63788 12414 63834 12474
rect 64876 12472 67699 12474
rect 64876 12416 67638 12472
rect 67694 12416 67699 12472
rect 64876 12414 67699 12416
rect 63788 12412 63794 12414
rect 63677 12411 63743 12412
rect 64876 12341 64936 12414
rect 67633 12411 67699 12414
rect 60273 12338 60339 12341
rect 61101 12338 61167 12341
rect 60273 12336 61167 12338
rect 60273 12280 60278 12336
rect 60334 12280 61106 12336
rect 61162 12280 61167 12336
rect 60273 12278 61167 12280
rect 60273 12275 60339 12278
rect 61101 12275 61167 12278
rect 62481 12338 62547 12341
rect 64873 12338 64939 12341
rect 62481 12336 64939 12338
rect 62481 12280 62486 12336
rect 62542 12280 64878 12336
rect 64934 12280 64939 12336
rect 62481 12278 64939 12280
rect 62481 12275 62547 12278
rect 64873 12275 64939 12278
rect 65977 12338 66043 12341
rect 70209 12338 70275 12341
rect 65977 12336 70275 12338
rect 65977 12280 65982 12336
rect 66038 12280 70214 12336
rect 70270 12280 70275 12336
rect 65977 12278 70275 12280
rect 65977 12275 66043 12278
rect 70209 12275 70275 12278
rect 88057 12338 88123 12341
rect 89200 12338 90000 12368
rect 88057 12336 90000 12338
rect 88057 12280 88062 12336
rect 88118 12280 90000 12336
rect 88057 12278 90000 12280
rect 88057 12275 88123 12278
rect 89200 12248 90000 12278
rect 63309 12202 63375 12205
rect 52913 12200 59738 12202
rect 52913 12144 52918 12200
rect 52974 12144 59738 12200
rect 52913 12142 59738 12144
rect 60046 12200 63375 12202
rect 60046 12144 63314 12200
rect 63370 12144 63375 12200
rect 60046 12142 63375 12144
rect 52913 12139 52979 12142
rect 25313 12066 25379 12069
rect 26417 12066 26483 12069
rect 25313 12064 26483 12066
rect 25313 12008 25318 12064
rect 25374 12008 26422 12064
rect 26478 12008 26483 12064
rect 25313 12006 26483 12008
rect 25313 12003 25379 12006
rect 26417 12003 26483 12006
rect 28349 12066 28415 12069
rect 28901 12066 28967 12069
rect 28349 12064 28967 12066
rect 28349 12008 28354 12064
rect 28410 12008 28906 12064
rect 28962 12008 28967 12064
rect 28349 12006 28967 12008
rect 28349 12003 28415 12006
rect 28901 12003 28967 12006
rect 29545 12066 29611 12069
rect 33317 12066 33383 12069
rect 35065 12066 35131 12069
rect 29545 12064 35131 12066
rect 29545 12008 29550 12064
rect 29606 12008 33322 12064
rect 33378 12008 35070 12064
rect 35126 12008 35131 12064
rect 29545 12006 35131 12008
rect 29545 12003 29611 12006
rect 33317 12003 33383 12006
rect 35065 12003 35131 12006
rect 35249 12066 35315 12069
rect 36261 12066 36327 12069
rect 35249 12064 36327 12066
rect 35249 12008 35254 12064
rect 35310 12008 36266 12064
rect 36322 12008 36327 12064
rect 35249 12006 36327 12008
rect 35249 12003 35315 12006
rect 36261 12003 36327 12006
rect 39021 12066 39087 12069
rect 43989 12066 44055 12069
rect 39021 12064 44055 12066
rect 39021 12008 39026 12064
rect 39082 12008 43994 12064
rect 44050 12008 44055 12064
rect 39021 12006 44055 12008
rect 39021 12003 39087 12006
rect 43989 12003 44055 12006
rect 46749 12066 46815 12069
rect 48037 12066 48103 12069
rect 46749 12064 48103 12066
rect 46749 12008 46754 12064
rect 46810 12008 48042 12064
rect 48098 12008 48103 12064
rect 46749 12006 48103 12008
rect 46749 12003 46815 12006
rect 48037 12003 48103 12006
rect 48405 12066 48471 12069
rect 48865 12066 48931 12069
rect 48405 12064 48931 12066
rect 48405 12008 48410 12064
rect 48466 12008 48870 12064
rect 48926 12008 48931 12064
rect 48405 12006 48931 12008
rect 48405 12003 48471 12006
rect 48865 12003 48931 12006
rect 51349 12066 51415 12069
rect 59678 12066 59738 12142
rect 63309 12139 63375 12142
rect 63585 12202 63651 12205
rect 69749 12202 69815 12205
rect 63585 12200 69815 12202
rect 63585 12144 63590 12200
rect 63646 12144 69754 12200
rect 69810 12144 69815 12200
rect 63585 12142 69815 12144
rect 63585 12139 63651 12142
rect 69749 12139 69815 12142
rect 60457 12066 60523 12069
rect 51349 12064 59554 12066
rect 51349 12008 51354 12064
rect 51410 12008 59554 12064
rect 51349 12006 59554 12008
rect 59678 12064 60523 12066
rect 59678 12008 60462 12064
rect 60518 12008 60523 12064
rect 59678 12006 60523 12008
rect 51349 12003 51415 12006
rect 22894 12000 23210 12001
rect 22894 11936 22900 12000
rect 22964 11936 22980 12000
rect 23044 11936 23060 12000
rect 23124 11936 23140 12000
rect 23204 11936 23210 12000
rect 22894 11935 23210 11936
rect 44842 12000 45158 12001
rect 44842 11936 44848 12000
rect 44912 11936 44928 12000
rect 44992 11936 45008 12000
rect 45072 11936 45088 12000
rect 45152 11936 45158 12000
rect 44842 11935 45158 11936
rect 25037 11930 25103 11933
rect 26509 11930 26575 11933
rect 25037 11928 26575 11930
rect 25037 11872 25042 11928
rect 25098 11872 26514 11928
rect 26570 11872 26575 11928
rect 25037 11870 26575 11872
rect 25037 11867 25103 11870
rect 26509 11867 26575 11870
rect 29821 11930 29887 11933
rect 33869 11930 33935 11933
rect 29821 11928 33935 11930
rect 29821 11872 29826 11928
rect 29882 11872 33874 11928
rect 33930 11872 33935 11928
rect 29821 11870 33935 11872
rect 29821 11867 29887 11870
rect 33869 11867 33935 11870
rect 35801 11930 35867 11933
rect 37733 11930 37799 11933
rect 43345 11930 43411 11933
rect 35801 11928 43411 11930
rect 35801 11872 35806 11928
rect 35862 11872 37738 11928
rect 37794 11872 43350 11928
rect 43406 11872 43411 11928
rect 35801 11870 43411 11872
rect 35801 11867 35867 11870
rect 37733 11867 37799 11870
rect 43345 11867 43411 11870
rect 46749 11930 46815 11933
rect 54385 11930 54451 11933
rect 46749 11928 54451 11930
rect 46749 11872 46754 11928
rect 46810 11872 54390 11928
rect 54446 11872 54451 11928
rect 46749 11870 54451 11872
rect 46749 11867 46815 11870
rect 54385 11867 54451 11870
rect 54661 11930 54727 11933
rect 59261 11930 59327 11933
rect 54661 11928 59327 11930
rect 54661 11872 54666 11928
rect 54722 11872 59266 11928
rect 59322 11872 59327 11928
rect 54661 11870 59327 11872
rect 59494 11930 59554 12006
rect 60457 12003 60523 12006
rect 60641 12066 60707 12069
rect 62297 12066 62363 12069
rect 66161 12066 66227 12069
rect 60641 12064 66227 12066
rect 60641 12008 60646 12064
rect 60702 12008 62302 12064
rect 62358 12008 66166 12064
rect 66222 12008 66227 12064
rect 60641 12006 66227 12008
rect 60641 12003 60707 12006
rect 62297 12003 62363 12006
rect 66161 12003 66227 12006
rect 66790 12000 67106 12001
rect 66790 11936 66796 12000
rect 66860 11936 66876 12000
rect 66940 11936 66956 12000
rect 67020 11936 67036 12000
rect 67100 11936 67106 12000
rect 66790 11935 67106 11936
rect 63033 11930 63099 11933
rect 63769 11932 63835 11933
rect 63718 11930 63724 11932
rect 59494 11928 63099 11930
rect 59494 11872 63038 11928
rect 63094 11872 63099 11928
rect 59494 11870 63099 11872
rect 63678 11870 63724 11930
rect 63788 11928 63835 11932
rect 63830 11872 63835 11928
rect 54661 11867 54727 11870
rect 59261 11867 59327 11870
rect 63033 11867 63099 11870
rect 63718 11868 63724 11870
rect 63788 11868 63835 11872
rect 63769 11867 63835 11868
rect 25681 11794 25747 11797
rect 28809 11794 28875 11797
rect 25681 11792 28875 11794
rect 25681 11736 25686 11792
rect 25742 11736 28814 11792
rect 28870 11736 28875 11792
rect 25681 11734 28875 11736
rect 25681 11731 25747 11734
rect 28809 11731 28875 11734
rect 31753 11794 31819 11797
rect 34329 11794 34395 11797
rect 31753 11792 34395 11794
rect 31753 11736 31758 11792
rect 31814 11736 34334 11792
rect 34390 11736 34395 11792
rect 31753 11734 34395 11736
rect 31753 11731 31819 11734
rect 34329 11731 34395 11734
rect 35433 11794 35499 11797
rect 36721 11794 36787 11797
rect 35433 11792 36787 11794
rect 35433 11736 35438 11792
rect 35494 11736 36726 11792
rect 36782 11736 36787 11792
rect 35433 11734 36787 11736
rect 35433 11731 35499 11734
rect 36721 11731 36787 11734
rect 39389 11794 39455 11797
rect 60958 11794 60964 11796
rect 39389 11792 60964 11794
rect 39389 11736 39394 11792
rect 39450 11736 60964 11792
rect 39389 11734 60964 11736
rect 39389 11731 39455 11734
rect 60958 11732 60964 11734
rect 61028 11732 61034 11796
rect 61101 11794 61167 11797
rect 62665 11794 62731 11797
rect 61101 11792 62731 11794
rect 61101 11736 61106 11792
rect 61162 11736 62670 11792
rect 62726 11736 62731 11792
rect 61101 11734 62731 11736
rect 61101 11731 61167 11734
rect 62665 11731 62731 11734
rect 63401 11794 63467 11797
rect 64045 11794 64111 11797
rect 63401 11792 64111 11794
rect 63401 11736 63406 11792
rect 63462 11736 64050 11792
rect 64106 11736 64111 11792
rect 63401 11734 64111 11736
rect 63401 11731 63467 11734
rect 64045 11731 64111 11734
rect 66989 11794 67055 11797
rect 70853 11794 70919 11797
rect 66989 11792 70919 11794
rect 66989 11736 66994 11792
rect 67050 11736 70858 11792
rect 70914 11736 70919 11792
rect 66989 11734 70919 11736
rect 66989 11731 67055 11734
rect 70853 11731 70919 11734
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 21081 11658 21147 11661
rect 26049 11658 26115 11661
rect 21081 11656 26115 11658
rect 21081 11600 21086 11656
rect 21142 11600 26054 11656
rect 26110 11600 26115 11656
rect 21081 11598 26115 11600
rect 21081 11595 21147 11598
rect 26049 11595 26115 11598
rect 32857 11658 32923 11661
rect 35801 11658 35867 11661
rect 32857 11656 35867 11658
rect 32857 11600 32862 11656
rect 32918 11600 35806 11656
rect 35862 11600 35867 11656
rect 32857 11598 35867 11600
rect 32857 11595 32923 11598
rect 35801 11595 35867 11598
rect 36261 11658 36327 11661
rect 63585 11658 63651 11661
rect 36261 11656 63651 11658
rect 36261 11600 36266 11656
rect 36322 11600 63590 11656
rect 63646 11600 63651 11656
rect 36261 11598 63651 11600
rect 36261 11595 36327 11598
rect 63585 11595 63651 11598
rect 66805 11658 66871 11661
rect 69013 11658 69079 11661
rect 66805 11656 69079 11658
rect 66805 11600 66810 11656
rect 66866 11600 69018 11656
rect 69074 11600 69079 11656
rect 66805 11598 69079 11600
rect 66805 11595 66871 11598
rect 69013 11595 69079 11598
rect 88057 11658 88123 11661
rect 89200 11658 90000 11688
rect 88057 11656 90000 11658
rect 88057 11600 88062 11656
rect 88118 11600 90000 11656
rect 88057 11598 90000 11600
rect 88057 11595 88123 11598
rect 89200 11568 90000 11598
rect 25589 11522 25655 11525
rect 26325 11522 26391 11525
rect 25589 11520 26391 11522
rect 25589 11464 25594 11520
rect 25650 11464 26330 11520
rect 26386 11464 26391 11520
rect 25589 11462 26391 11464
rect 25589 11459 25655 11462
rect 26325 11459 26391 11462
rect 43713 11522 43779 11525
rect 48497 11522 48563 11525
rect 43713 11520 48563 11522
rect 43713 11464 43718 11520
rect 43774 11464 48502 11520
rect 48558 11464 48563 11520
rect 43713 11462 48563 11464
rect 43713 11459 43779 11462
rect 48497 11459 48563 11462
rect 49233 11522 49299 11525
rect 51349 11522 51415 11525
rect 49233 11520 51415 11522
rect 49233 11464 49238 11520
rect 49294 11464 51354 11520
rect 51410 11464 51415 11520
rect 49233 11462 51415 11464
rect 49233 11459 49299 11462
rect 51349 11459 51415 11462
rect 53833 11522 53899 11525
rect 55213 11522 55279 11525
rect 56409 11524 56475 11525
rect 56358 11522 56364 11524
rect 53833 11520 55279 11522
rect 53833 11464 53838 11520
rect 53894 11464 55218 11520
rect 55274 11464 55279 11520
rect 53833 11462 55279 11464
rect 56318 11462 56364 11522
rect 56428 11520 56475 11524
rect 56470 11464 56475 11520
rect 53833 11459 53899 11462
rect 55213 11459 55279 11462
rect 56358 11460 56364 11462
rect 56428 11460 56475 11464
rect 56409 11459 56475 11460
rect 56593 11522 56659 11525
rect 57513 11522 57579 11525
rect 56593 11520 57579 11522
rect 56593 11464 56598 11520
rect 56654 11464 57518 11520
rect 57574 11464 57579 11520
rect 56593 11462 57579 11464
rect 56593 11459 56659 11462
rect 57513 11459 57579 11462
rect 58341 11522 58407 11525
rect 60273 11522 60339 11525
rect 58341 11520 60339 11522
rect 58341 11464 58346 11520
rect 58402 11464 60278 11520
rect 60334 11464 60339 11520
rect 58341 11462 60339 11464
rect 58341 11459 58407 11462
rect 60273 11459 60339 11462
rect 60549 11522 60615 11525
rect 62941 11522 63007 11525
rect 60549 11520 63007 11522
rect 60549 11464 60554 11520
rect 60610 11464 62946 11520
rect 63002 11464 63007 11520
rect 60549 11462 63007 11464
rect 60549 11459 60615 11462
rect 62941 11459 63007 11462
rect 63585 11522 63651 11525
rect 63902 11522 63908 11524
rect 63585 11520 63908 11522
rect 63585 11464 63590 11520
rect 63646 11464 63908 11520
rect 63585 11462 63908 11464
rect 63585 11459 63651 11462
rect 63902 11460 63908 11462
rect 63972 11460 63978 11524
rect 68737 11522 68803 11525
rect 67590 11520 68803 11522
rect 67590 11464 68742 11520
rect 68798 11464 68803 11520
rect 67590 11462 68803 11464
rect 11920 11456 12236 11457
rect 11920 11392 11926 11456
rect 11990 11392 12006 11456
rect 12070 11392 12086 11456
rect 12150 11392 12166 11456
rect 12230 11392 12236 11456
rect 11920 11391 12236 11392
rect 33868 11456 34184 11457
rect 33868 11392 33874 11456
rect 33938 11392 33954 11456
rect 34018 11392 34034 11456
rect 34098 11392 34114 11456
rect 34178 11392 34184 11456
rect 33868 11391 34184 11392
rect 55816 11456 56132 11457
rect 55816 11392 55822 11456
rect 55886 11392 55902 11456
rect 55966 11392 55982 11456
rect 56046 11392 56062 11456
rect 56126 11392 56132 11456
rect 55816 11391 56132 11392
rect 14457 11386 14523 11389
rect 18873 11386 18939 11389
rect 14457 11384 18939 11386
rect 14457 11328 14462 11384
rect 14518 11328 18878 11384
rect 18934 11328 18939 11384
rect 14457 11326 18939 11328
rect 14457 11323 14523 11326
rect 18873 11323 18939 11326
rect 21541 11386 21607 11389
rect 25865 11386 25931 11389
rect 21541 11384 25931 11386
rect 21541 11328 21546 11384
rect 21602 11328 25870 11384
rect 25926 11328 25931 11384
rect 21541 11326 25931 11328
rect 21541 11323 21607 11326
rect 25865 11323 25931 11326
rect 38285 11386 38351 11389
rect 47117 11386 47183 11389
rect 38285 11384 47183 11386
rect 38285 11328 38290 11384
rect 38346 11328 47122 11384
rect 47178 11328 47183 11384
rect 38285 11326 47183 11328
rect 38285 11323 38351 11326
rect 47117 11323 47183 11326
rect 47301 11386 47367 11389
rect 53833 11386 53899 11389
rect 60774 11386 60780 11388
rect 47301 11384 53899 11386
rect 47301 11328 47306 11384
rect 47362 11328 53838 11384
rect 53894 11328 53899 11384
rect 47301 11326 53899 11328
rect 47301 11323 47367 11326
rect 53833 11323 53899 11326
rect 56366 11326 60780 11386
rect 24301 11250 24367 11253
rect 26233 11250 26299 11253
rect 24301 11248 26299 11250
rect 24301 11192 24306 11248
rect 24362 11192 26238 11248
rect 26294 11192 26299 11248
rect 24301 11190 26299 11192
rect 24301 11187 24367 11190
rect 26233 11187 26299 11190
rect 37089 11250 37155 11253
rect 38929 11250 38995 11253
rect 37089 11248 38995 11250
rect 37089 11192 37094 11248
rect 37150 11192 38934 11248
rect 38990 11192 38995 11248
rect 37089 11190 38995 11192
rect 37089 11187 37155 11190
rect 38929 11187 38995 11190
rect 41137 11250 41203 11253
rect 43713 11250 43779 11253
rect 41137 11248 43779 11250
rect 41137 11192 41142 11248
rect 41198 11192 43718 11248
rect 43774 11192 43779 11248
rect 41137 11190 43779 11192
rect 41137 11187 41203 11190
rect 43713 11187 43779 11190
rect 44357 11250 44423 11253
rect 56366 11250 56426 11326
rect 60774 11324 60780 11326
rect 60844 11324 60850 11388
rect 60958 11324 60964 11388
rect 61028 11386 61034 11388
rect 67590 11386 67650 11462
rect 68737 11459 68803 11462
rect 77764 11456 78080 11457
rect 77764 11392 77770 11456
rect 77834 11392 77850 11456
rect 77914 11392 77930 11456
rect 77994 11392 78010 11456
rect 78074 11392 78080 11456
rect 77764 11391 78080 11392
rect 61028 11326 67650 11386
rect 67817 11386 67883 11389
rect 69197 11386 69263 11389
rect 67817 11384 69263 11386
rect 67817 11328 67822 11384
rect 67878 11328 69202 11384
rect 69258 11328 69263 11384
rect 67817 11326 69263 11328
rect 61028 11324 61034 11326
rect 67817 11323 67883 11326
rect 69197 11323 69263 11326
rect 44357 11248 56426 11250
rect 44357 11192 44362 11248
rect 44418 11192 56426 11248
rect 44357 11190 56426 11192
rect 58065 11250 58131 11253
rect 58801 11250 58867 11253
rect 64321 11252 64387 11253
rect 58065 11248 58867 11250
rect 58065 11192 58070 11248
rect 58126 11192 58806 11248
rect 58862 11192 58867 11248
rect 58065 11190 58867 11192
rect 44357 11187 44423 11190
rect 58065 11187 58131 11190
rect 58801 11187 58867 11190
rect 64270 11188 64276 11252
rect 64340 11250 64387 11252
rect 66529 11250 66595 11253
rect 67541 11250 67607 11253
rect 64340 11248 64432 11250
rect 64382 11192 64432 11248
rect 64340 11190 64432 11192
rect 66529 11248 67607 11250
rect 66529 11192 66534 11248
rect 66590 11192 67546 11248
rect 67602 11192 67607 11248
rect 66529 11190 67607 11192
rect 64340 11188 64387 11190
rect 64321 11187 64387 11188
rect 66529 11187 66595 11190
rect 67541 11187 67607 11190
rect 67725 11250 67791 11253
rect 69381 11250 69447 11253
rect 67725 11248 69447 11250
rect 67725 11192 67730 11248
rect 67786 11192 69386 11248
rect 69442 11192 69447 11248
rect 67725 11190 69447 11192
rect 67725 11187 67791 11190
rect 69381 11187 69447 11190
rect 24301 11114 24367 11117
rect 28901 11114 28967 11117
rect 30741 11114 30807 11117
rect 38101 11114 38167 11117
rect 24301 11112 30807 11114
rect 24301 11056 24306 11112
rect 24362 11056 28906 11112
rect 28962 11056 30746 11112
rect 30802 11056 30807 11112
rect 24301 11054 30807 11056
rect 24301 11051 24367 11054
rect 28901 11051 28967 11054
rect 30741 11051 30807 11054
rect 37230 11112 38167 11114
rect 37230 11056 38106 11112
rect 38162 11056 38167 11112
rect 37230 11054 38167 11056
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 29729 10978 29795 10981
rect 37230 10978 37290 11054
rect 38101 11051 38167 11054
rect 44817 11114 44883 11117
rect 45829 11114 45895 11117
rect 44817 11112 45895 11114
rect 44817 11056 44822 11112
rect 44878 11056 45834 11112
rect 45890 11056 45895 11112
rect 44817 11054 45895 11056
rect 44817 11051 44883 11054
rect 45829 11051 45895 11054
rect 49601 11114 49667 11117
rect 52269 11114 52335 11117
rect 49601 11112 52335 11114
rect 49601 11056 49606 11112
rect 49662 11056 52274 11112
rect 52330 11056 52335 11112
rect 49601 11054 52335 11056
rect 49601 11051 49667 11054
rect 52269 11051 52335 11054
rect 55213 11114 55279 11117
rect 60774 11114 60780 11116
rect 55213 11112 60780 11114
rect 55213 11056 55218 11112
rect 55274 11056 60780 11112
rect 55213 11054 60780 11056
rect 55213 11051 55279 11054
rect 60774 11052 60780 11054
rect 60844 11052 60850 11116
rect 60958 11052 60964 11116
rect 61028 11114 61034 11116
rect 64505 11114 64571 11117
rect 61028 11112 64571 11114
rect 61028 11056 64510 11112
rect 64566 11056 64571 11112
rect 61028 11054 64571 11056
rect 61028 11052 61034 11054
rect 64505 11051 64571 11054
rect 64873 11114 64939 11117
rect 69289 11114 69355 11117
rect 64873 11112 69355 11114
rect 64873 11056 64878 11112
rect 64934 11056 69294 11112
rect 69350 11056 69355 11112
rect 64873 11054 69355 11056
rect 64873 11051 64939 11054
rect 69289 11051 69355 11054
rect 29729 10976 37290 10978
rect 29729 10920 29734 10976
rect 29790 10920 37290 10976
rect 29729 10918 37290 10920
rect 37733 10978 37799 10981
rect 41137 10978 41203 10981
rect 37733 10976 41203 10978
rect 37733 10920 37738 10976
rect 37794 10920 41142 10976
rect 41198 10920 41203 10976
rect 37733 10918 41203 10920
rect 29729 10915 29795 10918
rect 37733 10915 37799 10918
rect 41137 10915 41203 10918
rect 50889 10978 50955 10981
rect 51349 10978 51415 10981
rect 50889 10976 51415 10978
rect 50889 10920 50894 10976
rect 50950 10920 51354 10976
rect 51410 10920 51415 10976
rect 50889 10918 51415 10920
rect 50889 10915 50955 10918
rect 51349 10915 51415 10918
rect 53741 10978 53807 10981
rect 59353 10978 59419 10981
rect 53741 10976 59419 10978
rect 53741 10920 53746 10976
rect 53802 10920 59358 10976
rect 59414 10920 59419 10976
rect 53741 10918 59419 10920
rect 53741 10915 53807 10918
rect 59353 10915 59419 10918
rect 60641 10978 60707 10981
rect 62849 10978 62915 10981
rect 60641 10976 62915 10978
rect 60641 10920 60646 10976
rect 60702 10920 62854 10976
rect 62910 10920 62915 10976
rect 60641 10918 62915 10920
rect 60641 10915 60707 10918
rect 62849 10915 62915 10918
rect 87413 10978 87479 10981
rect 89200 10978 90000 11008
rect 87413 10976 90000 10978
rect 87413 10920 87418 10976
rect 87474 10920 90000 10976
rect 87413 10918 90000 10920
rect 87413 10915 87479 10918
rect 22894 10912 23210 10913
rect 22894 10848 22900 10912
rect 22964 10848 22980 10912
rect 23044 10848 23060 10912
rect 23124 10848 23140 10912
rect 23204 10848 23210 10912
rect 22894 10847 23210 10848
rect 44842 10912 45158 10913
rect 44842 10848 44848 10912
rect 44912 10848 44928 10912
rect 44992 10848 45008 10912
rect 45072 10848 45088 10912
rect 45152 10848 45158 10912
rect 44842 10847 45158 10848
rect 66790 10912 67106 10913
rect 66790 10848 66796 10912
rect 66860 10848 66876 10912
rect 66940 10848 66956 10912
rect 67020 10848 67036 10912
rect 67100 10848 67106 10912
rect 89200 10888 90000 10918
rect 66790 10847 67106 10848
rect 31477 10842 31543 10845
rect 37089 10842 37155 10845
rect 31477 10840 37155 10842
rect 31477 10784 31482 10840
rect 31538 10784 37094 10840
rect 37150 10784 37155 10840
rect 31477 10782 37155 10784
rect 31477 10779 31543 10782
rect 37089 10779 37155 10782
rect 38837 10842 38903 10845
rect 39481 10842 39547 10845
rect 38837 10840 39547 10842
rect 38837 10784 38842 10840
rect 38898 10784 39486 10840
rect 39542 10784 39547 10840
rect 38837 10782 39547 10784
rect 38837 10779 38903 10782
rect 39481 10779 39547 10782
rect 49509 10842 49575 10845
rect 53373 10842 53439 10845
rect 49509 10840 53439 10842
rect 49509 10784 49514 10840
rect 49570 10784 53378 10840
rect 53434 10784 53439 10840
rect 49509 10782 53439 10784
rect 49509 10779 49575 10782
rect 53373 10779 53439 10782
rect 53649 10842 53715 10845
rect 63401 10842 63467 10845
rect 53649 10840 63467 10842
rect 53649 10784 53654 10840
rect 53710 10784 63406 10840
rect 63462 10784 63467 10840
rect 53649 10782 63467 10784
rect 53649 10779 53715 10782
rect 63401 10779 63467 10782
rect 1577 10706 1643 10709
rect 56961 10706 57027 10709
rect 1577 10704 57027 10706
rect 1577 10648 1582 10704
rect 1638 10648 56966 10704
rect 57022 10648 57027 10704
rect 1577 10646 57027 10648
rect 1577 10643 1643 10646
rect 56961 10643 57027 10646
rect 63033 10706 63099 10709
rect 63401 10706 63467 10709
rect 63033 10704 63467 10706
rect 63033 10648 63038 10704
rect 63094 10648 63406 10704
rect 63462 10648 63467 10704
rect 63033 10646 63467 10648
rect 63033 10643 63099 10646
rect 63401 10643 63467 10646
rect 38561 10570 38627 10573
rect 41413 10570 41479 10573
rect 38561 10568 41479 10570
rect 38561 10512 38566 10568
rect 38622 10512 41418 10568
rect 41474 10512 41479 10568
rect 38561 10510 41479 10512
rect 38561 10507 38627 10510
rect 41413 10507 41479 10510
rect 45277 10570 45343 10573
rect 46749 10570 46815 10573
rect 45277 10568 46815 10570
rect 45277 10512 45282 10568
rect 45338 10512 46754 10568
rect 46810 10512 46815 10568
rect 45277 10510 46815 10512
rect 45277 10507 45343 10510
rect 46749 10507 46815 10510
rect 52637 10570 52703 10573
rect 53465 10570 53531 10573
rect 59629 10570 59695 10573
rect 52637 10568 59695 10570
rect 52637 10512 52642 10568
rect 52698 10512 53470 10568
rect 53526 10512 59634 10568
rect 59690 10512 59695 10568
rect 52637 10510 59695 10512
rect 52637 10507 52703 10510
rect 53465 10507 53531 10510
rect 59629 10507 59695 10510
rect 60774 10508 60780 10572
rect 60844 10570 60850 10572
rect 63769 10570 63835 10573
rect 60844 10568 63835 10570
rect 60844 10512 63774 10568
rect 63830 10512 63835 10568
rect 60844 10510 63835 10512
rect 60844 10508 60850 10510
rect 63769 10507 63835 10510
rect 45185 10434 45251 10437
rect 47209 10434 47275 10437
rect 45185 10432 47275 10434
rect 45185 10376 45190 10432
rect 45246 10376 47214 10432
rect 47270 10376 47275 10432
rect 45185 10374 47275 10376
rect 45185 10371 45251 10374
rect 47209 10371 47275 10374
rect 52545 10434 52611 10437
rect 55397 10434 55463 10437
rect 52545 10432 55463 10434
rect 52545 10376 52550 10432
rect 52606 10376 55402 10432
rect 55458 10376 55463 10432
rect 52545 10374 55463 10376
rect 52545 10371 52611 10374
rect 55397 10371 55463 10374
rect 61837 10434 61903 10437
rect 67449 10434 67515 10437
rect 61837 10432 67515 10434
rect 61837 10376 61842 10432
rect 61898 10376 67454 10432
rect 67510 10376 67515 10432
rect 61837 10374 67515 10376
rect 61837 10371 61903 10374
rect 67449 10371 67515 10374
rect 11920 10368 12236 10369
rect 0 10298 800 10328
rect 11920 10304 11926 10368
rect 11990 10304 12006 10368
rect 12070 10304 12086 10368
rect 12150 10304 12166 10368
rect 12230 10304 12236 10368
rect 11920 10303 12236 10304
rect 33868 10368 34184 10369
rect 33868 10304 33874 10368
rect 33938 10304 33954 10368
rect 34018 10304 34034 10368
rect 34098 10304 34114 10368
rect 34178 10304 34184 10368
rect 33868 10303 34184 10304
rect 55816 10368 56132 10369
rect 55816 10304 55822 10368
rect 55886 10304 55902 10368
rect 55966 10304 55982 10368
rect 56046 10304 56062 10368
rect 56126 10304 56132 10368
rect 55816 10303 56132 10304
rect 77764 10368 78080 10369
rect 77764 10304 77770 10368
rect 77834 10304 77850 10368
rect 77914 10304 77930 10368
rect 77994 10304 78010 10368
rect 78074 10304 78080 10368
rect 77764 10303 78080 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 42149 10298 42215 10301
rect 52085 10298 52151 10301
rect 42149 10296 52151 10298
rect 42149 10240 42154 10296
rect 42210 10240 52090 10296
rect 52146 10240 52151 10296
rect 42149 10238 52151 10240
rect 42149 10235 42215 10238
rect 52085 10235 52151 10238
rect 56910 10236 56916 10300
rect 56980 10298 56986 10300
rect 63493 10298 63559 10301
rect 56980 10296 63559 10298
rect 56980 10240 63498 10296
rect 63554 10240 63559 10296
rect 56980 10238 63559 10240
rect 56980 10236 56986 10238
rect 63493 10235 63559 10238
rect 88057 10298 88123 10301
rect 89200 10298 90000 10328
rect 88057 10296 90000 10298
rect 88057 10240 88062 10296
rect 88118 10240 90000 10296
rect 88057 10238 90000 10240
rect 88057 10235 88123 10238
rect 89200 10208 90000 10238
rect 43345 10162 43411 10165
rect 47853 10162 47919 10165
rect 43345 10160 47919 10162
rect 43345 10104 43350 10160
rect 43406 10104 47858 10160
rect 47914 10104 47919 10160
rect 43345 10102 47919 10104
rect 43345 10099 43411 10102
rect 47853 10099 47919 10102
rect 50797 10162 50863 10165
rect 57605 10162 57671 10165
rect 50797 10160 57671 10162
rect 50797 10104 50802 10160
rect 50858 10104 57610 10160
rect 57666 10104 57671 10160
rect 50797 10102 57671 10104
rect 50797 10099 50863 10102
rect 57605 10099 57671 10102
rect 38653 10026 38719 10029
rect 39113 10026 39179 10029
rect 38653 10024 39179 10026
rect 38653 9968 38658 10024
rect 38714 9968 39118 10024
rect 39174 9968 39179 10024
rect 38653 9966 39179 9968
rect 38653 9963 38719 9966
rect 39113 9963 39179 9966
rect 22894 9824 23210 9825
rect 22894 9760 22900 9824
rect 22964 9760 22980 9824
rect 23044 9760 23060 9824
rect 23124 9760 23140 9824
rect 23204 9760 23210 9824
rect 22894 9759 23210 9760
rect 44842 9824 45158 9825
rect 44842 9760 44848 9824
rect 44912 9760 44928 9824
rect 44992 9760 45008 9824
rect 45072 9760 45088 9824
rect 45152 9760 45158 9824
rect 44842 9759 45158 9760
rect 66790 9824 67106 9825
rect 66790 9760 66796 9824
rect 66860 9760 66876 9824
rect 66940 9760 66956 9824
rect 67020 9760 67036 9824
rect 67100 9760 67106 9824
rect 66790 9759 67106 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 11920 9280 12236 9281
rect 11920 9216 11926 9280
rect 11990 9216 12006 9280
rect 12070 9216 12086 9280
rect 12150 9216 12166 9280
rect 12230 9216 12236 9280
rect 11920 9215 12236 9216
rect 33868 9280 34184 9281
rect 33868 9216 33874 9280
rect 33938 9216 33954 9280
rect 34018 9216 34034 9280
rect 34098 9216 34114 9280
rect 34178 9216 34184 9280
rect 33868 9215 34184 9216
rect 55816 9280 56132 9281
rect 55816 9216 55822 9280
rect 55886 9216 55902 9280
rect 55966 9216 55982 9280
rect 56046 9216 56062 9280
rect 56126 9216 56132 9280
rect 55816 9215 56132 9216
rect 77764 9280 78080 9281
rect 77764 9216 77770 9280
rect 77834 9216 77850 9280
rect 77914 9216 77930 9280
rect 77994 9216 78010 9280
rect 78074 9216 78080 9280
rect 77764 9215 78080 9216
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 87413 8938 87479 8941
rect 89200 8938 90000 8968
rect 87413 8936 90000 8938
rect 87413 8880 87418 8936
rect 87474 8880 90000 8936
rect 87413 8878 90000 8880
rect 87413 8875 87479 8878
rect 89200 8848 90000 8878
rect 22894 8736 23210 8737
rect 22894 8672 22900 8736
rect 22964 8672 22980 8736
rect 23044 8672 23060 8736
rect 23124 8672 23140 8736
rect 23204 8672 23210 8736
rect 22894 8671 23210 8672
rect 44842 8736 45158 8737
rect 44842 8672 44848 8736
rect 44912 8672 44928 8736
rect 44992 8672 45008 8736
rect 45072 8672 45088 8736
rect 45152 8672 45158 8736
rect 44842 8671 45158 8672
rect 66790 8736 67106 8737
rect 66790 8672 66796 8736
rect 66860 8672 66876 8736
rect 66940 8672 66956 8736
rect 67020 8672 67036 8736
rect 67100 8672 67106 8736
rect 66790 8671 67106 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 88241 8258 88307 8261
rect 89200 8258 90000 8288
rect 88241 8256 90000 8258
rect 88241 8200 88246 8256
rect 88302 8200 90000 8256
rect 88241 8198 90000 8200
rect 88241 8195 88307 8198
rect 11920 8192 12236 8193
rect 11920 8128 11926 8192
rect 11990 8128 12006 8192
rect 12070 8128 12086 8192
rect 12150 8128 12166 8192
rect 12230 8128 12236 8192
rect 11920 8127 12236 8128
rect 33868 8192 34184 8193
rect 33868 8128 33874 8192
rect 33938 8128 33954 8192
rect 34018 8128 34034 8192
rect 34098 8128 34114 8192
rect 34178 8128 34184 8192
rect 33868 8127 34184 8128
rect 55816 8192 56132 8193
rect 55816 8128 55822 8192
rect 55886 8128 55902 8192
rect 55966 8128 55982 8192
rect 56046 8128 56062 8192
rect 56126 8128 56132 8192
rect 55816 8127 56132 8128
rect 77764 8192 78080 8193
rect 77764 8128 77770 8192
rect 77834 8128 77850 8192
rect 77914 8128 77930 8192
rect 77994 8128 78010 8192
rect 78074 8128 78080 8192
rect 89200 8168 90000 8198
rect 77764 8127 78080 8128
rect 22894 7648 23210 7649
rect 22894 7584 22900 7648
rect 22964 7584 22980 7648
rect 23044 7584 23060 7648
rect 23124 7584 23140 7648
rect 23204 7584 23210 7648
rect 22894 7583 23210 7584
rect 44842 7648 45158 7649
rect 44842 7584 44848 7648
rect 44912 7584 44928 7648
rect 44992 7584 45008 7648
rect 45072 7584 45088 7648
rect 45152 7584 45158 7648
rect 44842 7583 45158 7584
rect 66790 7648 67106 7649
rect 66790 7584 66796 7648
rect 66860 7584 66876 7648
rect 66940 7584 66956 7648
rect 67020 7584 67036 7648
rect 67100 7584 67106 7648
rect 66790 7583 67106 7584
rect 88057 7578 88123 7581
rect 89200 7578 90000 7608
rect 88057 7576 90000 7578
rect 88057 7520 88062 7576
rect 88118 7520 90000 7576
rect 88057 7518 90000 7520
rect 88057 7515 88123 7518
rect 89200 7488 90000 7518
rect 11920 7104 12236 7105
rect 11920 7040 11926 7104
rect 11990 7040 12006 7104
rect 12070 7040 12086 7104
rect 12150 7040 12166 7104
rect 12230 7040 12236 7104
rect 11920 7039 12236 7040
rect 33868 7104 34184 7105
rect 33868 7040 33874 7104
rect 33938 7040 33954 7104
rect 34018 7040 34034 7104
rect 34098 7040 34114 7104
rect 34178 7040 34184 7104
rect 33868 7039 34184 7040
rect 55816 7104 56132 7105
rect 55816 7040 55822 7104
rect 55886 7040 55902 7104
rect 55966 7040 55982 7104
rect 56046 7040 56062 7104
rect 56126 7040 56132 7104
rect 55816 7039 56132 7040
rect 77764 7104 78080 7105
rect 77764 7040 77770 7104
rect 77834 7040 77850 7104
rect 77914 7040 77930 7104
rect 77994 7040 78010 7104
rect 78074 7040 78080 7104
rect 77764 7039 78080 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 88057 6898 88123 6901
rect 89200 6898 90000 6928
rect 88057 6896 90000 6898
rect 88057 6840 88062 6896
rect 88118 6840 90000 6896
rect 88057 6838 90000 6840
rect 88057 6835 88123 6838
rect 89200 6808 90000 6838
rect 22894 6560 23210 6561
rect 22894 6496 22900 6560
rect 22964 6496 22980 6560
rect 23044 6496 23060 6560
rect 23124 6496 23140 6560
rect 23204 6496 23210 6560
rect 22894 6495 23210 6496
rect 44842 6560 45158 6561
rect 44842 6496 44848 6560
rect 44912 6496 44928 6560
rect 44992 6496 45008 6560
rect 45072 6496 45088 6560
rect 45152 6496 45158 6560
rect 44842 6495 45158 6496
rect 66790 6560 67106 6561
rect 66790 6496 66796 6560
rect 66860 6496 66876 6560
rect 66940 6496 66956 6560
rect 67020 6496 67036 6560
rect 67100 6496 67106 6560
rect 66790 6495 67106 6496
rect 0 6218 800 6248
rect 1761 6218 1827 6221
rect 0 6216 1827 6218
rect 0 6160 1766 6216
rect 1822 6160 1827 6216
rect 0 6158 1827 6160
rect 0 6128 800 6158
rect 1761 6155 1827 6158
rect 87413 6218 87479 6221
rect 89200 6218 90000 6248
rect 87413 6216 90000 6218
rect 87413 6160 87418 6216
rect 87474 6160 90000 6216
rect 87413 6158 90000 6160
rect 87413 6155 87479 6158
rect 89200 6128 90000 6158
rect 11920 6016 12236 6017
rect 11920 5952 11926 6016
rect 11990 5952 12006 6016
rect 12070 5952 12086 6016
rect 12150 5952 12166 6016
rect 12230 5952 12236 6016
rect 11920 5951 12236 5952
rect 33868 6016 34184 6017
rect 33868 5952 33874 6016
rect 33938 5952 33954 6016
rect 34018 5952 34034 6016
rect 34098 5952 34114 6016
rect 34178 5952 34184 6016
rect 33868 5951 34184 5952
rect 55816 6016 56132 6017
rect 55816 5952 55822 6016
rect 55886 5952 55902 6016
rect 55966 5952 55982 6016
rect 56046 5952 56062 6016
rect 56126 5952 56132 6016
rect 55816 5951 56132 5952
rect 77764 6016 78080 6017
rect 77764 5952 77770 6016
rect 77834 5952 77850 6016
rect 77914 5952 77930 6016
rect 77994 5952 78010 6016
rect 78074 5952 78080 6016
rect 77764 5951 78080 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 87965 5538 88031 5541
rect 89200 5538 90000 5568
rect 87965 5536 90000 5538
rect 87965 5480 87970 5536
rect 88026 5480 90000 5536
rect 87965 5478 90000 5480
rect 87965 5475 88031 5478
rect 22894 5472 23210 5473
rect 22894 5408 22900 5472
rect 22964 5408 22980 5472
rect 23044 5408 23060 5472
rect 23124 5408 23140 5472
rect 23204 5408 23210 5472
rect 22894 5407 23210 5408
rect 44842 5472 45158 5473
rect 44842 5408 44848 5472
rect 44912 5408 44928 5472
rect 44992 5408 45008 5472
rect 45072 5408 45088 5472
rect 45152 5408 45158 5472
rect 44842 5407 45158 5408
rect 66790 5472 67106 5473
rect 66790 5408 66796 5472
rect 66860 5408 66876 5472
rect 66940 5408 66956 5472
rect 67020 5408 67036 5472
rect 67100 5408 67106 5472
rect 89200 5448 90000 5478
rect 66790 5407 67106 5408
rect 11920 4928 12236 4929
rect 0 4768 800 4888
rect 11920 4864 11926 4928
rect 11990 4864 12006 4928
rect 12070 4864 12086 4928
rect 12150 4864 12166 4928
rect 12230 4864 12236 4928
rect 11920 4863 12236 4864
rect 33868 4928 34184 4929
rect 33868 4864 33874 4928
rect 33938 4864 33954 4928
rect 34018 4864 34034 4928
rect 34098 4864 34114 4928
rect 34178 4864 34184 4928
rect 33868 4863 34184 4864
rect 55816 4928 56132 4929
rect 55816 4864 55822 4928
rect 55886 4864 55902 4928
rect 55966 4864 55982 4928
rect 56046 4864 56062 4928
rect 56126 4864 56132 4928
rect 55816 4863 56132 4864
rect 77764 4928 78080 4929
rect 77764 4864 77770 4928
rect 77834 4864 77850 4928
rect 77914 4864 77930 4928
rect 77994 4864 78010 4928
rect 78074 4864 78080 4928
rect 77764 4863 78080 4864
rect 88057 4858 88123 4861
rect 89200 4858 90000 4888
rect 88057 4856 90000 4858
rect 88057 4800 88062 4856
rect 88118 4800 90000 4856
rect 88057 4798 90000 4800
rect 88057 4795 88123 4798
rect 89200 4768 90000 4798
rect 22894 4384 23210 4385
rect 22894 4320 22900 4384
rect 22964 4320 22980 4384
rect 23044 4320 23060 4384
rect 23124 4320 23140 4384
rect 23204 4320 23210 4384
rect 22894 4319 23210 4320
rect 44842 4384 45158 4385
rect 44842 4320 44848 4384
rect 44912 4320 44928 4384
rect 44992 4320 45008 4384
rect 45072 4320 45088 4384
rect 45152 4320 45158 4384
rect 44842 4319 45158 4320
rect 66790 4384 67106 4385
rect 66790 4320 66796 4384
rect 66860 4320 66876 4384
rect 66940 4320 66956 4384
rect 67020 4320 67036 4384
rect 67100 4320 67106 4384
rect 66790 4319 67106 4320
rect 0 4178 800 4208
rect 1577 4178 1643 4181
rect 0 4176 1643 4178
rect 0 4120 1582 4176
rect 1638 4120 1643 4176
rect 0 4118 1643 4120
rect 0 4088 800 4118
rect 1577 4115 1643 4118
rect 88057 4178 88123 4181
rect 89200 4178 90000 4208
rect 88057 4176 90000 4178
rect 88057 4120 88062 4176
rect 88118 4120 90000 4176
rect 88057 4118 90000 4120
rect 88057 4115 88123 4118
rect 89200 4088 90000 4118
rect 43437 4042 43503 4045
rect 46473 4042 46539 4045
rect 43437 4040 46539 4042
rect 43437 3984 43442 4040
rect 43498 3984 46478 4040
rect 46534 3984 46539 4040
rect 43437 3982 46539 3984
rect 43437 3979 43503 3982
rect 46473 3979 46539 3982
rect 51441 4042 51507 4045
rect 52545 4042 52611 4045
rect 51441 4040 52611 4042
rect 51441 3984 51446 4040
rect 51502 3984 52550 4040
rect 52606 3984 52611 4040
rect 51441 3982 52611 3984
rect 51441 3979 51507 3982
rect 52545 3979 52611 3982
rect 11920 3840 12236 3841
rect 11920 3776 11926 3840
rect 11990 3776 12006 3840
rect 12070 3776 12086 3840
rect 12150 3776 12166 3840
rect 12230 3776 12236 3840
rect 11920 3775 12236 3776
rect 33868 3840 34184 3841
rect 33868 3776 33874 3840
rect 33938 3776 33954 3840
rect 34018 3776 34034 3840
rect 34098 3776 34114 3840
rect 34178 3776 34184 3840
rect 33868 3775 34184 3776
rect 55816 3840 56132 3841
rect 55816 3776 55822 3840
rect 55886 3776 55902 3840
rect 55966 3776 55982 3840
rect 56046 3776 56062 3840
rect 56126 3776 56132 3840
rect 55816 3775 56132 3776
rect 77764 3840 78080 3841
rect 77764 3776 77770 3840
rect 77834 3776 77850 3840
rect 77914 3776 77930 3840
rect 77994 3776 78010 3840
rect 78074 3776 78080 3840
rect 77764 3775 78080 3776
rect 42609 3770 42675 3773
rect 48221 3770 48287 3773
rect 42609 3768 48287 3770
rect 42609 3712 42614 3768
rect 42670 3712 48226 3768
rect 48282 3712 48287 3768
rect 42609 3710 48287 3712
rect 42609 3707 42675 3710
rect 48221 3707 48287 3710
rect 0 3498 800 3528
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 800 3438
rect 1393 3435 1459 3438
rect 43437 3498 43503 3501
rect 48129 3498 48195 3501
rect 43437 3496 48195 3498
rect 43437 3440 43442 3496
rect 43498 3440 48134 3496
rect 48190 3440 48195 3496
rect 43437 3438 48195 3440
rect 43437 3435 43503 3438
rect 48129 3435 48195 3438
rect 48865 3498 48931 3501
rect 49509 3498 49575 3501
rect 48865 3496 49575 3498
rect 48865 3440 48870 3496
rect 48926 3440 49514 3496
rect 49570 3440 49575 3496
rect 48865 3438 49575 3440
rect 48865 3435 48931 3438
rect 49509 3435 49575 3438
rect 50521 3498 50587 3501
rect 51809 3498 51875 3501
rect 52913 3498 52979 3501
rect 50521 3496 52979 3498
rect 50521 3440 50526 3496
rect 50582 3440 51814 3496
rect 51870 3440 52918 3496
rect 52974 3440 52979 3496
rect 50521 3438 52979 3440
rect 50521 3435 50587 3438
rect 51809 3435 51875 3438
rect 52913 3435 52979 3438
rect 88333 3498 88399 3501
rect 89200 3498 90000 3528
rect 88333 3496 90000 3498
rect 88333 3440 88338 3496
rect 88394 3440 90000 3496
rect 88333 3438 90000 3440
rect 88333 3435 88399 3438
rect 89200 3408 90000 3438
rect 50245 3362 50311 3365
rect 52177 3362 52243 3365
rect 50245 3360 52243 3362
rect 50245 3304 50250 3360
rect 50306 3304 52182 3360
rect 52238 3304 52243 3360
rect 50245 3302 52243 3304
rect 50245 3299 50311 3302
rect 52177 3299 52243 3302
rect 22894 3296 23210 3297
rect 22894 3232 22900 3296
rect 22964 3232 22980 3296
rect 23044 3232 23060 3296
rect 23124 3232 23140 3296
rect 23204 3232 23210 3296
rect 22894 3231 23210 3232
rect 44842 3296 45158 3297
rect 44842 3232 44848 3296
rect 44912 3232 44928 3296
rect 44992 3232 45008 3296
rect 45072 3232 45088 3296
rect 45152 3232 45158 3296
rect 44842 3231 45158 3232
rect 66790 3296 67106 3297
rect 66790 3232 66796 3296
rect 66860 3232 66876 3296
rect 66940 3232 66956 3296
rect 67020 3232 67036 3296
rect 67100 3232 67106 3296
rect 66790 3231 67106 3232
rect 49233 3226 49299 3229
rect 51993 3226 52059 3229
rect 49233 3224 52059 3226
rect 49233 3168 49238 3224
rect 49294 3168 51998 3224
rect 52054 3168 52059 3224
rect 49233 3166 52059 3168
rect 49233 3163 49299 3166
rect 51993 3163 52059 3166
rect 25957 3090 26023 3093
rect 28533 3090 28599 3093
rect 25957 3088 28599 3090
rect 25957 3032 25962 3088
rect 26018 3032 28538 3088
rect 28594 3032 28599 3088
rect 25957 3030 28599 3032
rect 25957 3027 26023 3030
rect 28533 3027 28599 3030
rect 39941 2954 40007 2957
rect 45277 2954 45343 2957
rect 39941 2952 45343 2954
rect 39941 2896 39946 2952
rect 40002 2896 45282 2952
rect 45338 2896 45343 2952
rect 39941 2894 45343 2896
rect 39941 2891 40007 2894
rect 45277 2891 45343 2894
rect 45461 2954 45527 2957
rect 49785 2954 49851 2957
rect 45461 2952 49851 2954
rect 45461 2896 45466 2952
rect 45522 2896 49790 2952
rect 49846 2896 49851 2952
rect 45461 2894 49851 2896
rect 45461 2891 45527 2894
rect 49785 2891 49851 2894
rect 0 2818 800 2848
rect 1485 2818 1551 2821
rect 0 2816 1551 2818
rect 0 2760 1490 2816
rect 1546 2760 1551 2816
rect 0 2758 1551 2760
rect 0 2728 800 2758
rect 1485 2755 1551 2758
rect 40953 2818 41019 2821
rect 45553 2818 45619 2821
rect 40953 2816 45619 2818
rect 40953 2760 40958 2816
rect 41014 2760 45558 2816
rect 45614 2760 45619 2816
rect 40953 2758 45619 2760
rect 40953 2755 41019 2758
rect 45553 2755 45619 2758
rect 46565 2818 46631 2821
rect 50613 2818 50679 2821
rect 46565 2816 50679 2818
rect 46565 2760 46570 2816
rect 46626 2760 50618 2816
rect 50674 2760 50679 2816
rect 46565 2758 50679 2760
rect 46565 2755 46631 2758
rect 50613 2755 50679 2758
rect 88057 2818 88123 2821
rect 89200 2818 90000 2848
rect 88057 2816 90000 2818
rect 88057 2760 88062 2816
rect 88118 2760 90000 2816
rect 88057 2758 90000 2760
rect 88057 2755 88123 2758
rect 11920 2752 12236 2753
rect 11920 2688 11926 2752
rect 11990 2688 12006 2752
rect 12070 2688 12086 2752
rect 12150 2688 12166 2752
rect 12230 2688 12236 2752
rect 11920 2687 12236 2688
rect 33868 2752 34184 2753
rect 33868 2688 33874 2752
rect 33938 2688 33954 2752
rect 34018 2688 34034 2752
rect 34098 2688 34114 2752
rect 34178 2688 34184 2752
rect 33868 2687 34184 2688
rect 55816 2752 56132 2753
rect 55816 2688 55822 2752
rect 55886 2688 55902 2752
rect 55966 2688 55982 2752
rect 56046 2688 56062 2752
rect 56126 2688 56132 2752
rect 55816 2687 56132 2688
rect 77764 2752 78080 2753
rect 77764 2688 77770 2752
rect 77834 2688 77850 2752
rect 77914 2688 77930 2752
rect 77994 2688 78010 2752
rect 78074 2688 78080 2752
rect 89200 2728 90000 2758
rect 77764 2687 78080 2688
rect 26325 2546 26391 2549
rect 80789 2546 80855 2549
rect 26325 2544 80855 2546
rect 26325 2488 26330 2544
rect 26386 2488 80794 2544
rect 80850 2488 80855 2544
rect 26325 2486 80855 2488
rect 26325 2483 26391 2486
rect 80789 2483 80855 2486
rect 2681 2410 2747 2413
rect 56501 2410 56567 2413
rect 2681 2408 56567 2410
rect 2681 2352 2686 2408
rect 2742 2352 56506 2408
rect 56562 2352 56567 2408
rect 2681 2350 56567 2352
rect 2681 2347 2747 2350
rect 56501 2347 56567 2350
rect 24209 2274 24275 2277
rect 28257 2274 28323 2277
rect 24209 2272 28323 2274
rect 24209 2216 24214 2272
rect 24270 2216 28262 2272
rect 28318 2216 28323 2272
rect 24209 2214 28323 2216
rect 24209 2211 24275 2214
rect 28257 2211 28323 2214
rect 22894 2208 23210 2209
rect 0 2138 800 2168
rect 22894 2144 22900 2208
rect 22964 2144 22980 2208
rect 23044 2144 23060 2208
rect 23124 2144 23140 2208
rect 23204 2144 23210 2208
rect 22894 2143 23210 2144
rect 44842 2208 45158 2209
rect 44842 2144 44848 2208
rect 44912 2144 44928 2208
rect 44992 2144 45008 2208
rect 45072 2144 45088 2208
rect 45152 2144 45158 2208
rect 44842 2143 45158 2144
rect 66790 2208 67106 2209
rect 66790 2144 66796 2208
rect 66860 2144 66876 2208
rect 66940 2144 66956 2208
rect 67020 2144 67036 2208
rect 67100 2144 67106 2208
rect 66790 2143 67106 2144
rect 2957 2138 3023 2141
rect 0 2136 3023 2138
rect 0 2080 2962 2136
rect 3018 2080 3023 2136
rect 0 2078 3023 2080
rect 0 2048 800 2078
rect 2957 2075 3023 2078
rect 34053 2138 34119 2141
rect 40309 2138 40375 2141
rect 34053 2136 40375 2138
rect 34053 2080 34058 2136
rect 34114 2080 40314 2136
rect 40370 2080 40375 2136
rect 34053 2078 40375 2080
rect 34053 2075 34119 2078
rect 40309 2075 40375 2078
rect 88149 2138 88215 2141
rect 89200 2138 90000 2168
rect 88149 2136 90000 2138
rect 88149 2080 88154 2136
rect 88210 2080 90000 2136
rect 88149 2078 90000 2080
rect 88149 2075 88215 2078
rect 89200 2048 90000 2078
rect 30281 2002 30347 2005
rect 31845 2002 31911 2005
rect 30281 2000 31911 2002
rect 30281 1944 30286 2000
rect 30342 1944 31850 2000
rect 31906 1944 31911 2000
rect 30281 1942 31911 1944
rect 30281 1939 30347 1942
rect 31845 1939 31911 1942
rect 45553 2002 45619 2005
rect 48865 2002 48931 2005
rect 45553 2000 48931 2002
rect 45553 1944 45558 2000
rect 45614 1944 48870 2000
rect 48926 1944 48931 2000
rect 45553 1942 48931 1944
rect 45553 1939 45619 1942
rect 48865 1939 48931 1942
rect 26325 1866 26391 1869
rect 31661 1866 31727 1869
rect 26325 1864 31727 1866
rect 26325 1808 26330 1864
rect 26386 1808 31666 1864
rect 31722 1808 31727 1864
rect 26325 1806 31727 1808
rect 26325 1803 26391 1806
rect 31661 1803 31727 1806
rect 38653 1866 38719 1869
rect 45829 1866 45895 1869
rect 38653 1864 45895 1866
rect 38653 1808 38658 1864
rect 38714 1808 45834 1864
rect 45890 1808 45895 1864
rect 38653 1806 45895 1808
rect 38653 1803 38719 1806
rect 45829 1803 45895 1806
rect 31753 1730 31819 1733
rect 35709 1730 35775 1733
rect 31753 1728 35775 1730
rect 31753 1672 31758 1728
rect 31814 1672 35714 1728
rect 35770 1672 35775 1728
rect 31753 1670 35775 1672
rect 31753 1667 31819 1670
rect 35709 1667 35775 1670
rect 45553 1730 45619 1733
rect 48497 1730 48563 1733
rect 45553 1728 48563 1730
rect 45553 1672 45558 1728
rect 45614 1672 48502 1728
rect 48558 1672 48563 1728
rect 45553 1670 48563 1672
rect 45553 1667 45619 1670
rect 48497 1667 48563 1670
rect 27245 1594 27311 1597
rect 31845 1594 31911 1597
rect 27245 1592 31911 1594
rect 27245 1536 27250 1592
rect 27306 1536 31850 1592
rect 31906 1536 31911 1592
rect 27245 1534 31911 1536
rect 27245 1531 27311 1534
rect 31845 1531 31911 1534
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 4061 914 4127 917
rect 2454 912 4127 914
rect 2454 856 4066 912
rect 4122 856 4127 912
rect 2454 854 4127 856
rect 0 778 800 808
rect 2454 778 2514 854
rect 4061 851 4127 854
rect 86861 914 86927 917
rect 86861 912 86970 914
rect 86861 856 86866 912
rect 86922 856 86970 912
rect 86861 851 86970 856
rect 0 718 2514 778
rect 86910 778 86970 851
rect 89200 778 90000 808
rect 86910 718 90000 778
rect 0 688 800 718
rect 89200 688 90000 718
rect 86677 98 86743 101
rect 89200 98 90000 128
rect 86677 96 90000 98
rect 86677 40 86682 96
rect 86738 40 90000 96
rect 86677 38 90000 40
rect 86677 35 86743 38
rect 89200 8 90000 38
<< via3 >>
rect 11926 27772 11990 27776
rect 11926 27716 11930 27772
rect 11930 27716 11986 27772
rect 11986 27716 11990 27772
rect 11926 27712 11990 27716
rect 12006 27772 12070 27776
rect 12006 27716 12010 27772
rect 12010 27716 12066 27772
rect 12066 27716 12070 27772
rect 12006 27712 12070 27716
rect 12086 27772 12150 27776
rect 12086 27716 12090 27772
rect 12090 27716 12146 27772
rect 12146 27716 12150 27772
rect 12086 27712 12150 27716
rect 12166 27772 12230 27776
rect 12166 27716 12170 27772
rect 12170 27716 12226 27772
rect 12226 27716 12230 27772
rect 12166 27712 12230 27716
rect 33874 27772 33938 27776
rect 33874 27716 33878 27772
rect 33878 27716 33934 27772
rect 33934 27716 33938 27772
rect 33874 27712 33938 27716
rect 33954 27772 34018 27776
rect 33954 27716 33958 27772
rect 33958 27716 34014 27772
rect 34014 27716 34018 27772
rect 33954 27712 34018 27716
rect 34034 27772 34098 27776
rect 34034 27716 34038 27772
rect 34038 27716 34094 27772
rect 34094 27716 34098 27772
rect 34034 27712 34098 27716
rect 34114 27772 34178 27776
rect 34114 27716 34118 27772
rect 34118 27716 34174 27772
rect 34174 27716 34178 27772
rect 34114 27712 34178 27716
rect 55822 27772 55886 27776
rect 55822 27716 55826 27772
rect 55826 27716 55882 27772
rect 55882 27716 55886 27772
rect 55822 27712 55886 27716
rect 55902 27772 55966 27776
rect 55902 27716 55906 27772
rect 55906 27716 55962 27772
rect 55962 27716 55966 27772
rect 55902 27712 55966 27716
rect 55982 27772 56046 27776
rect 55982 27716 55986 27772
rect 55986 27716 56042 27772
rect 56042 27716 56046 27772
rect 55982 27712 56046 27716
rect 56062 27772 56126 27776
rect 56062 27716 56066 27772
rect 56066 27716 56122 27772
rect 56122 27716 56126 27772
rect 56062 27712 56126 27716
rect 77770 27772 77834 27776
rect 77770 27716 77774 27772
rect 77774 27716 77830 27772
rect 77830 27716 77834 27772
rect 77770 27712 77834 27716
rect 77850 27772 77914 27776
rect 77850 27716 77854 27772
rect 77854 27716 77910 27772
rect 77910 27716 77914 27772
rect 77850 27712 77914 27716
rect 77930 27772 77994 27776
rect 77930 27716 77934 27772
rect 77934 27716 77990 27772
rect 77990 27716 77994 27772
rect 77930 27712 77994 27716
rect 78010 27772 78074 27776
rect 78010 27716 78014 27772
rect 78014 27716 78070 27772
rect 78070 27716 78074 27772
rect 78010 27712 78074 27716
rect 22900 27228 22964 27232
rect 22900 27172 22904 27228
rect 22904 27172 22960 27228
rect 22960 27172 22964 27228
rect 22900 27168 22964 27172
rect 22980 27228 23044 27232
rect 22980 27172 22984 27228
rect 22984 27172 23040 27228
rect 23040 27172 23044 27228
rect 22980 27168 23044 27172
rect 23060 27228 23124 27232
rect 23060 27172 23064 27228
rect 23064 27172 23120 27228
rect 23120 27172 23124 27228
rect 23060 27168 23124 27172
rect 23140 27228 23204 27232
rect 23140 27172 23144 27228
rect 23144 27172 23200 27228
rect 23200 27172 23204 27228
rect 23140 27168 23204 27172
rect 44848 27228 44912 27232
rect 44848 27172 44852 27228
rect 44852 27172 44908 27228
rect 44908 27172 44912 27228
rect 44848 27168 44912 27172
rect 44928 27228 44992 27232
rect 44928 27172 44932 27228
rect 44932 27172 44988 27228
rect 44988 27172 44992 27228
rect 44928 27168 44992 27172
rect 45008 27228 45072 27232
rect 45008 27172 45012 27228
rect 45012 27172 45068 27228
rect 45068 27172 45072 27228
rect 45008 27168 45072 27172
rect 45088 27228 45152 27232
rect 45088 27172 45092 27228
rect 45092 27172 45148 27228
rect 45148 27172 45152 27228
rect 45088 27168 45152 27172
rect 66796 27228 66860 27232
rect 66796 27172 66800 27228
rect 66800 27172 66856 27228
rect 66856 27172 66860 27228
rect 66796 27168 66860 27172
rect 66876 27228 66940 27232
rect 66876 27172 66880 27228
rect 66880 27172 66936 27228
rect 66936 27172 66940 27228
rect 66876 27168 66940 27172
rect 66956 27228 67020 27232
rect 66956 27172 66960 27228
rect 66960 27172 67016 27228
rect 67016 27172 67020 27228
rect 66956 27168 67020 27172
rect 67036 27228 67100 27232
rect 67036 27172 67040 27228
rect 67040 27172 67096 27228
rect 67096 27172 67100 27228
rect 67036 27168 67100 27172
rect 11926 26684 11990 26688
rect 11926 26628 11930 26684
rect 11930 26628 11986 26684
rect 11986 26628 11990 26684
rect 11926 26624 11990 26628
rect 12006 26684 12070 26688
rect 12006 26628 12010 26684
rect 12010 26628 12066 26684
rect 12066 26628 12070 26684
rect 12006 26624 12070 26628
rect 12086 26684 12150 26688
rect 12086 26628 12090 26684
rect 12090 26628 12146 26684
rect 12146 26628 12150 26684
rect 12086 26624 12150 26628
rect 12166 26684 12230 26688
rect 12166 26628 12170 26684
rect 12170 26628 12226 26684
rect 12226 26628 12230 26684
rect 12166 26624 12230 26628
rect 33874 26684 33938 26688
rect 33874 26628 33878 26684
rect 33878 26628 33934 26684
rect 33934 26628 33938 26684
rect 33874 26624 33938 26628
rect 33954 26684 34018 26688
rect 33954 26628 33958 26684
rect 33958 26628 34014 26684
rect 34014 26628 34018 26684
rect 33954 26624 34018 26628
rect 34034 26684 34098 26688
rect 34034 26628 34038 26684
rect 34038 26628 34094 26684
rect 34094 26628 34098 26684
rect 34034 26624 34098 26628
rect 34114 26684 34178 26688
rect 34114 26628 34118 26684
rect 34118 26628 34174 26684
rect 34174 26628 34178 26684
rect 34114 26624 34178 26628
rect 55822 26684 55886 26688
rect 55822 26628 55826 26684
rect 55826 26628 55882 26684
rect 55882 26628 55886 26684
rect 55822 26624 55886 26628
rect 55902 26684 55966 26688
rect 55902 26628 55906 26684
rect 55906 26628 55962 26684
rect 55962 26628 55966 26684
rect 55902 26624 55966 26628
rect 55982 26684 56046 26688
rect 55982 26628 55986 26684
rect 55986 26628 56042 26684
rect 56042 26628 56046 26684
rect 55982 26624 56046 26628
rect 56062 26684 56126 26688
rect 56062 26628 56066 26684
rect 56066 26628 56122 26684
rect 56122 26628 56126 26684
rect 56062 26624 56126 26628
rect 77770 26684 77834 26688
rect 77770 26628 77774 26684
rect 77774 26628 77830 26684
rect 77830 26628 77834 26684
rect 77770 26624 77834 26628
rect 77850 26684 77914 26688
rect 77850 26628 77854 26684
rect 77854 26628 77910 26684
rect 77910 26628 77914 26684
rect 77850 26624 77914 26628
rect 77930 26684 77994 26688
rect 77930 26628 77934 26684
rect 77934 26628 77990 26684
rect 77990 26628 77994 26684
rect 77930 26624 77994 26628
rect 78010 26684 78074 26688
rect 78010 26628 78014 26684
rect 78014 26628 78070 26684
rect 78070 26628 78074 26684
rect 78010 26624 78074 26628
rect 22900 26140 22964 26144
rect 22900 26084 22904 26140
rect 22904 26084 22960 26140
rect 22960 26084 22964 26140
rect 22900 26080 22964 26084
rect 22980 26140 23044 26144
rect 22980 26084 22984 26140
rect 22984 26084 23040 26140
rect 23040 26084 23044 26140
rect 22980 26080 23044 26084
rect 23060 26140 23124 26144
rect 23060 26084 23064 26140
rect 23064 26084 23120 26140
rect 23120 26084 23124 26140
rect 23060 26080 23124 26084
rect 23140 26140 23204 26144
rect 23140 26084 23144 26140
rect 23144 26084 23200 26140
rect 23200 26084 23204 26140
rect 23140 26080 23204 26084
rect 44848 26140 44912 26144
rect 44848 26084 44852 26140
rect 44852 26084 44908 26140
rect 44908 26084 44912 26140
rect 44848 26080 44912 26084
rect 44928 26140 44992 26144
rect 44928 26084 44932 26140
rect 44932 26084 44988 26140
rect 44988 26084 44992 26140
rect 44928 26080 44992 26084
rect 45008 26140 45072 26144
rect 45008 26084 45012 26140
rect 45012 26084 45068 26140
rect 45068 26084 45072 26140
rect 45008 26080 45072 26084
rect 45088 26140 45152 26144
rect 45088 26084 45092 26140
rect 45092 26084 45148 26140
rect 45148 26084 45152 26140
rect 45088 26080 45152 26084
rect 66796 26140 66860 26144
rect 66796 26084 66800 26140
rect 66800 26084 66856 26140
rect 66856 26084 66860 26140
rect 66796 26080 66860 26084
rect 66876 26140 66940 26144
rect 66876 26084 66880 26140
rect 66880 26084 66936 26140
rect 66936 26084 66940 26140
rect 66876 26080 66940 26084
rect 66956 26140 67020 26144
rect 66956 26084 66960 26140
rect 66960 26084 67016 26140
rect 67016 26084 67020 26140
rect 66956 26080 67020 26084
rect 67036 26140 67100 26144
rect 67036 26084 67040 26140
rect 67040 26084 67096 26140
rect 67096 26084 67100 26140
rect 67036 26080 67100 26084
rect 28028 25740 28092 25804
rect 11926 25596 11990 25600
rect 11926 25540 11930 25596
rect 11930 25540 11986 25596
rect 11986 25540 11990 25596
rect 11926 25536 11990 25540
rect 12006 25596 12070 25600
rect 12006 25540 12010 25596
rect 12010 25540 12066 25596
rect 12066 25540 12070 25596
rect 12006 25536 12070 25540
rect 12086 25596 12150 25600
rect 12086 25540 12090 25596
rect 12090 25540 12146 25596
rect 12146 25540 12150 25596
rect 12086 25536 12150 25540
rect 12166 25596 12230 25600
rect 12166 25540 12170 25596
rect 12170 25540 12226 25596
rect 12226 25540 12230 25596
rect 12166 25536 12230 25540
rect 33874 25596 33938 25600
rect 33874 25540 33878 25596
rect 33878 25540 33934 25596
rect 33934 25540 33938 25596
rect 33874 25536 33938 25540
rect 33954 25596 34018 25600
rect 33954 25540 33958 25596
rect 33958 25540 34014 25596
rect 34014 25540 34018 25596
rect 33954 25536 34018 25540
rect 34034 25596 34098 25600
rect 34034 25540 34038 25596
rect 34038 25540 34094 25596
rect 34094 25540 34098 25596
rect 34034 25536 34098 25540
rect 34114 25596 34178 25600
rect 34114 25540 34118 25596
rect 34118 25540 34174 25596
rect 34174 25540 34178 25596
rect 34114 25536 34178 25540
rect 55822 25596 55886 25600
rect 55822 25540 55826 25596
rect 55826 25540 55882 25596
rect 55882 25540 55886 25596
rect 55822 25536 55886 25540
rect 55902 25596 55966 25600
rect 55902 25540 55906 25596
rect 55906 25540 55962 25596
rect 55962 25540 55966 25596
rect 55902 25536 55966 25540
rect 55982 25596 56046 25600
rect 55982 25540 55986 25596
rect 55986 25540 56042 25596
rect 56042 25540 56046 25596
rect 55982 25536 56046 25540
rect 56062 25596 56126 25600
rect 56062 25540 56066 25596
rect 56066 25540 56122 25596
rect 56122 25540 56126 25596
rect 56062 25536 56126 25540
rect 77770 25596 77834 25600
rect 77770 25540 77774 25596
rect 77774 25540 77830 25596
rect 77830 25540 77834 25596
rect 77770 25536 77834 25540
rect 77850 25596 77914 25600
rect 77850 25540 77854 25596
rect 77854 25540 77910 25596
rect 77910 25540 77914 25596
rect 77850 25536 77914 25540
rect 77930 25596 77994 25600
rect 77930 25540 77934 25596
rect 77934 25540 77990 25596
rect 77990 25540 77994 25596
rect 77930 25536 77994 25540
rect 78010 25596 78074 25600
rect 78010 25540 78014 25596
rect 78014 25540 78070 25596
rect 78070 25540 78074 25596
rect 78010 25536 78074 25540
rect 22900 25052 22964 25056
rect 22900 24996 22904 25052
rect 22904 24996 22960 25052
rect 22960 24996 22964 25052
rect 22900 24992 22964 24996
rect 22980 25052 23044 25056
rect 22980 24996 22984 25052
rect 22984 24996 23040 25052
rect 23040 24996 23044 25052
rect 22980 24992 23044 24996
rect 23060 25052 23124 25056
rect 23060 24996 23064 25052
rect 23064 24996 23120 25052
rect 23120 24996 23124 25052
rect 23060 24992 23124 24996
rect 23140 25052 23204 25056
rect 23140 24996 23144 25052
rect 23144 24996 23200 25052
rect 23200 24996 23204 25052
rect 23140 24992 23204 24996
rect 44848 25052 44912 25056
rect 44848 24996 44852 25052
rect 44852 24996 44908 25052
rect 44908 24996 44912 25052
rect 44848 24992 44912 24996
rect 44928 25052 44992 25056
rect 44928 24996 44932 25052
rect 44932 24996 44988 25052
rect 44988 24996 44992 25052
rect 44928 24992 44992 24996
rect 45008 25052 45072 25056
rect 45008 24996 45012 25052
rect 45012 24996 45068 25052
rect 45068 24996 45072 25052
rect 45008 24992 45072 24996
rect 45088 25052 45152 25056
rect 45088 24996 45092 25052
rect 45092 24996 45148 25052
rect 45148 24996 45152 25052
rect 45088 24992 45152 24996
rect 66796 25052 66860 25056
rect 66796 24996 66800 25052
rect 66800 24996 66856 25052
rect 66856 24996 66860 25052
rect 66796 24992 66860 24996
rect 66876 25052 66940 25056
rect 66876 24996 66880 25052
rect 66880 24996 66936 25052
rect 66936 24996 66940 25052
rect 66876 24992 66940 24996
rect 66956 25052 67020 25056
rect 66956 24996 66960 25052
rect 66960 24996 67016 25052
rect 67016 24996 67020 25052
rect 66956 24992 67020 24996
rect 67036 25052 67100 25056
rect 67036 24996 67040 25052
rect 67040 24996 67096 25052
rect 67096 24996 67100 25052
rect 67036 24992 67100 24996
rect 11926 24508 11990 24512
rect 11926 24452 11930 24508
rect 11930 24452 11986 24508
rect 11986 24452 11990 24508
rect 11926 24448 11990 24452
rect 12006 24508 12070 24512
rect 12006 24452 12010 24508
rect 12010 24452 12066 24508
rect 12066 24452 12070 24508
rect 12006 24448 12070 24452
rect 12086 24508 12150 24512
rect 12086 24452 12090 24508
rect 12090 24452 12146 24508
rect 12146 24452 12150 24508
rect 12086 24448 12150 24452
rect 12166 24508 12230 24512
rect 12166 24452 12170 24508
rect 12170 24452 12226 24508
rect 12226 24452 12230 24508
rect 12166 24448 12230 24452
rect 33874 24508 33938 24512
rect 33874 24452 33878 24508
rect 33878 24452 33934 24508
rect 33934 24452 33938 24508
rect 33874 24448 33938 24452
rect 33954 24508 34018 24512
rect 33954 24452 33958 24508
rect 33958 24452 34014 24508
rect 34014 24452 34018 24508
rect 33954 24448 34018 24452
rect 34034 24508 34098 24512
rect 34034 24452 34038 24508
rect 34038 24452 34094 24508
rect 34094 24452 34098 24508
rect 34034 24448 34098 24452
rect 34114 24508 34178 24512
rect 34114 24452 34118 24508
rect 34118 24452 34174 24508
rect 34174 24452 34178 24508
rect 34114 24448 34178 24452
rect 55822 24508 55886 24512
rect 55822 24452 55826 24508
rect 55826 24452 55882 24508
rect 55882 24452 55886 24508
rect 55822 24448 55886 24452
rect 55902 24508 55966 24512
rect 55902 24452 55906 24508
rect 55906 24452 55962 24508
rect 55962 24452 55966 24508
rect 55902 24448 55966 24452
rect 55982 24508 56046 24512
rect 55982 24452 55986 24508
rect 55986 24452 56042 24508
rect 56042 24452 56046 24508
rect 55982 24448 56046 24452
rect 56062 24508 56126 24512
rect 56062 24452 56066 24508
rect 56066 24452 56122 24508
rect 56122 24452 56126 24508
rect 56062 24448 56126 24452
rect 77770 24508 77834 24512
rect 77770 24452 77774 24508
rect 77774 24452 77830 24508
rect 77830 24452 77834 24508
rect 77770 24448 77834 24452
rect 77850 24508 77914 24512
rect 77850 24452 77854 24508
rect 77854 24452 77910 24508
rect 77910 24452 77914 24508
rect 77850 24448 77914 24452
rect 77930 24508 77994 24512
rect 77930 24452 77934 24508
rect 77934 24452 77990 24508
rect 77990 24452 77994 24508
rect 77930 24448 77994 24452
rect 78010 24508 78074 24512
rect 78010 24452 78014 24508
rect 78014 24452 78070 24508
rect 78070 24452 78074 24508
rect 78010 24448 78074 24452
rect 27476 24108 27540 24172
rect 22900 23964 22964 23968
rect 22900 23908 22904 23964
rect 22904 23908 22960 23964
rect 22960 23908 22964 23964
rect 22900 23904 22964 23908
rect 22980 23964 23044 23968
rect 22980 23908 22984 23964
rect 22984 23908 23040 23964
rect 23040 23908 23044 23964
rect 22980 23904 23044 23908
rect 23060 23964 23124 23968
rect 23060 23908 23064 23964
rect 23064 23908 23120 23964
rect 23120 23908 23124 23964
rect 23060 23904 23124 23908
rect 23140 23964 23204 23968
rect 23140 23908 23144 23964
rect 23144 23908 23200 23964
rect 23200 23908 23204 23964
rect 23140 23904 23204 23908
rect 44848 23964 44912 23968
rect 44848 23908 44852 23964
rect 44852 23908 44908 23964
rect 44908 23908 44912 23964
rect 44848 23904 44912 23908
rect 44928 23964 44992 23968
rect 44928 23908 44932 23964
rect 44932 23908 44988 23964
rect 44988 23908 44992 23964
rect 44928 23904 44992 23908
rect 45008 23964 45072 23968
rect 45008 23908 45012 23964
rect 45012 23908 45068 23964
rect 45068 23908 45072 23964
rect 45008 23904 45072 23908
rect 45088 23964 45152 23968
rect 45088 23908 45092 23964
rect 45092 23908 45148 23964
rect 45148 23908 45152 23964
rect 45088 23904 45152 23908
rect 66796 23964 66860 23968
rect 66796 23908 66800 23964
rect 66800 23908 66856 23964
rect 66856 23908 66860 23964
rect 66796 23904 66860 23908
rect 66876 23964 66940 23968
rect 66876 23908 66880 23964
rect 66880 23908 66936 23964
rect 66936 23908 66940 23964
rect 66876 23904 66940 23908
rect 66956 23964 67020 23968
rect 66956 23908 66960 23964
rect 66960 23908 67016 23964
rect 67016 23908 67020 23964
rect 66956 23904 67020 23908
rect 67036 23964 67100 23968
rect 67036 23908 67040 23964
rect 67040 23908 67096 23964
rect 67096 23908 67100 23964
rect 67036 23904 67100 23908
rect 11926 23420 11990 23424
rect 11926 23364 11930 23420
rect 11930 23364 11986 23420
rect 11986 23364 11990 23420
rect 11926 23360 11990 23364
rect 12006 23420 12070 23424
rect 12006 23364 12010 23420
rect 12010 23364 12066 23420
rect 12066 23364 12070 23420
rect 12006 23360 12070 23364
rect 12086 23420 12150 23424
rect 12086 23364 12090 23420
rect 12090 23364 12146 23420
rect 12146 23364 12150 23420
rect 12086 23360 12150 23364
rect 12166 23420 12230 23424
rect 12166 23364 12170 23420
rect 12170 23364 12226 23420
rect 12226 23364 12230 23420
rect 12166 23360 12230 23364
rect 33874 23420 33938 23424
rect 33874 23364 33878 23420
rect 33878 23364 33934 23420
rect 33934 23364 33938 23420
rect 33874 23360 33938 23364
rect 33954 23420 34018 23424
rect 33954 23364 33958 23420
rect 33958 23364 34014 23420
rect 34014 23364 34018 23420
rect 33954 23360 34018 23364
rect 34034 23420 34098 23424
rect 34034 23364 34038 23420
rect 34038 23364 34094 23420
rect 34094 23364 34098 23420
rect 34034 23360 34098 23364
rect 34114 23420 34178 23424
rect 34114 23364 34118 23420
rect 34118 23364 34174 23420
rect 34174 23364 34178 23420
rect 34114 23360 34178 23364
rect 55822 23420 55886 23424
rect 55822 23364 55826 23420
rect 55826 23364 55882 23420
rect 55882 23364 55886 23420
rect 55822 23360 55886 23364
rect 55902 23420 55966 23424
rect 55902 23364 55906 23420
rect 55906 23364 55962 23420
rect 55962 23364 55966 23420
rect 55902 23360 55966 23364
rect 55982 23420 56046 23424
rect 55982 23364 55986 23420
rect 55986 23364 56042 23420
rect 56042 23364 56046 23420
rect 55982 23360 56046 23364
rect 56062 23420 56126 23424
rect 56062 23364 56066 23420
rect 56066 23364 56122 23420
rect 56122 23364 56126 23420
rect 56062 23360 56126 23364
rect 77770 23420 77834 23424
rect 77770 23364 77774 23420
rect 77774 23364 77830 23420
rect 77830 23364 77834 23420
rect 77770 23360 77834 23364
rect 77850 23420 77914 23424
rect 77850 23364 77854 23420
rect 77854 23364 77910 23420
rect 77910 23364 77914 23420
rect 77850 23360 77914 23364
rect 77930 23420 77994 23424
rect 77930 23364 77934 23420
rect 77934 23364 77990 23420
rect 77990 23364 77994 23420
rect 77930 23360 77994 23364
rect 78010 23420 78074 23424
rect 78010 23364 78014 23420
rect 78014 23364 78070 23420
rect 78070 23364 78074 23420
rect 78010 23360 78074 23364
rect 22900 22876 22964 22880
rect 22900 22820 22904 22876
rect 22904 22820 22960 22876
rect 22960 22820 22964 22876
rect 22900 22816 22964 22820
rect 22980 22876 23044 22880
rect 22980 22820 22984 22876
rect 22984 22820 23040 22876
rect 23040 22820 23044 22876
rect 22980 22816 23044 22820
rect 23060 22876 23124 22880
rect 23060 22820 23064 22876
rect 23064 22820 23120 22876
rect 23120 22820 23124 22876
rect 23060 22816 23124 22820
rect 23140 22876 23204 22880
rect 23140 22820 23144 22876
rect 23144 22820 23200 22876
rect 23200 22820 23204 22876
rect 23140 22816 23204 22820
rect 44848 22876 44912 22880
rect 44848 22820 44852 22876
rect 44852 22820 44908 22876
rect 44908 22820 44912 22876
rect 44848 22816 44912 22820
rect 44928 22876 44992 22880
rect 44928 22820 44932 22876
rect 44932 22820 44988 22876
rect 44988 22820 44992 22876
rect 44928 22816 44992 22820
rect 45008 22876 45072 22880
rect 45008 22820 45012 22876
rect 45012 22820 45068 22876
rect 45068 22820 45072 22876
rect 45008 22816 45072 22820
rect 45088 22876 45152 22880
rect 45088 22820 45092 22876
rect 45092 22820 45148 22876
rect 45148 22820 45152 22876
rect 45088 22816 45152 22820
rect 66796 22876 66860 22880
rect 66796 22820 66800 22876
rect 66800 22820 66856 22876
rect 66856 22820 66860 22876
rect 66796 22816 66860 22820
rect 66876 22876 66940 22880
rect 66876 22820 66880 22876
rect 66880 22820 66936 22876
rect 66936 22820 66940 22876
rect 66876 22816 66940 22820
rect 66956 22876 67020 22880
rect 66956 22820 66960 22876
rect 66960 22820 67016 22876
rect 67016 22820 67020 22876
rect 66956 22816 67020 22820
rect 67036 22876 67100 22880
rect 67036 22820 67040 22876
rect 67040 22820 67096 22876
rect 67096 22820 67100 22876
rect 67036 22816 67100 22820
rect 11926 22332 11990 22336
rect 11926 22276 11930 22332
rect 11930 22276 11986 22332
rect 11986 22276 11990 22332
rect 11926 22272 11990 22276
rect 12006 22332 12070 22336
rect 12006 22276 12010 22332
rect 12010 22276 12066 22332
rect 12066 22276 12070 22332
rect 12006 22272 12070 22276
rect 12086 22332 12150 22336
rect 12086 22276 12090 22332
rect 12090 22276 12146 22332
rect 12146 22276 12150 22332
rect 12086 22272 12150 22276
rect 12166 22332 12230 22336
rect 12166 22276 12170 22332
rect 12170 22276 12226 22332
rect 12226 22276 12230 22332
rect 12166 22272 12230 22276
rect 33874 22332 33938 22336
rect 33874 22276 33878 22332
rect 33878 22276 33934 22332
rect 33934 22276 33938 22332
rect 33874 22272 33938 22276
rect 33954 22332 34018 22336
rect 33954 22276 33958 22332
rect 33958 22276 34014 22332
rect 34014 22276 34018 22332
rect 33954 22272 34018 22276
rect 34034 22332 34098 22336
rect 34034 22276 34038 22332
rect 34038 22276 34094 22332
rect 34094 22276 34098 22332
rect 34034 22272 34098 22276
rect 34114 22332 34178 22336
rect 34114 22276 34118 22332
rect 34118 22276 34174 22332
rect 34174 22276 34178 22332
rect 34114 22272 34178 22276
rect 55822 22332 55886 22336
rect 55822 22276 55826 22332
rect 55826 22276 55882 22332
rect 55882 22276 55886 22332
rect 55822 22272 55886 22276
rect 55902 22332 55966 22336
rect 55902 22276 55906 22332
rect 55906 22276 55962 22332
rect 55962 22276 55966 22332
rect 55902 22272 55966 22276
rect 55982 22332 56046 22336
rect 55982 22276 55986 22332
rect 55986 22276 56042 22332
rect 56042 22276 56046 22332
rect 55982 22272 56046 22276
rect 56062 22332 56126 22336
rect 56062 22276 56066 22332
rect 56066 22276 56122 22332
rect 56122 22276 56126 22332
rect 56062 22272 56126 22276
rect 77770 22332 77834 22336
rect 77770 22276 77774 22332
rect 77774 22276 77830 22332
rect 77830 22276 77834 22332
rect 77770 22272 77834 22276
rect 77850 22332 77914 22336
rect 77850 22276 77854 22332
rect 77854 22276 77910 22332
rect 77910 22276 77914 22332
rect 77850 22272 77914 22276
rect 77930 22332 77994 22336
rect 77930 22276 77934 22332
rect 77934 22276 77990 22332
rect 77990 22276 77994 22332
rect 77930 22272 77994 22276
rect 78010 22332 78074 22336
rect 78010 22276 78014 22332
rect 78014 22276 78070 22332
rect 78070 22276 78074 22332
rect 78010 22272 78074 22276
rect 22900 21788 22964 21792
rect 22900 21732 22904 21788
rect 22904 21732 22960 21788
rect 22960 21732 22964 21788
rect 22900 21728 22964 21732
rect 22980 21788 23044 21792
rect 22980 21732 22984 21788
rect 22984 21732 23040 21788
rect 23040 21732 23044 21788
rect 22980 21728 23044 21732
rect 23060 21788 23124 21792
rect 23060 21732 23064 21788
rect 23064 21732 23120 21788
rect 23120 21732 23124 21788
rect 23060 21728 23124 21732
rect 23140 21788 23204 21792
rect 23140 21732 23144 21788
rect 23144 21732 23200 21788
rect 23200 21732 23204 21788
rect 23140 21728 23204 21732
rect 44848 21788 44912 21792
rect 44848 21732 44852 21788
rect 44852 21732 44908 21788
rect 44908 21732 44912 21788
rect 44848 21728 44912 21732
rect 44928 21788 44992 21792
rect 44928 21732 44932 21788
rect 44932 21732 44988 21788
rect 44988 21732 44992 21788
rect 44928 21728 44992 21732
rect 45008 21788 45072 21792
rect 45008 21732 45012 21788
rect 45012 21732 45068 21788
rect 45068 21732 45072 21788
rect 45008 21728 45072 21732
rect 45088 21788 45152 21792
rect 45088 21732 45092 21788
rect 45092 21732 45148 21788
rect 45148 21732 45152 21788
rect 45088 21728 45152 21732
rect 66796 21788 66860 21792
rect 66796 21732 66800 21788
rect 66800 21732 66856 21788
rect 66856 21732 66860 21788
rect 66796 21728 66860 21732
rect 66876 21788 66940 21792
rect 66876 21732 66880 21788
rect 66880 21732 66936 21788
rect 66936 21732 66940 21788
rect 66876 21728 66940 21732
rect 66956 21788 67020 21792
rect 66956 21732 66960 21788
rect 66960 21732 67016 21788
rect 67016 21732 67020 21788
rect 66956 21728 67020 21732
rect 67036 21788 67100 21792
rect 67036 21732 67040 21788
rect 67040 21732 67096 21788
rect 67096 21732 67100 21788
rect 67036 21728 67100 21732
rect 26556 21388 26620 21452
rect 11926 21244 11990 21248
rect 11926 21188 11930 21244
rect 11930 21188 11986 21244
rect 11986 21188 11990 21244
rect 11926 21184 11990 21188
rect 12006 21244 12070 21248
rect 12006 21188 12010 21244
rect 12010 21188 12066 21244
rect 12066 21188 12070 21244
rect 12006 21184 12070 21188
rect 12086 21244 12150 21248
rect 12086 21188 12090 21244
rect 12090 21188 12146 21244
rect 12146 21188 12150 21244
rect 12086 21184 12150 21188
rect 12166 21244 12230 21248
rect 12166 21188 12170 21244
rect 12170 21188 12226 21244
rect 12226 21188 12230 21244
rect 12166 21184 12230 21188
rect 33874 21244 33938 21248
rect 33874 21188 33878 21244
rect 33878 21188 33934 21244
rect 33934 21188 33938 21244
rect 33874 21184 33938 21188
rect 33954 21244 34018 21248
rect 33954 21188 33958 21244
rect 33958 21188 34014 21244
rect 34014 21188 34018 21244
rect 33954 21184 34018 21188
rect 34034 21244 34098 21248
rect 34034 21188 34038 21244
rect 34038 21188 34094 21244
rect 34094 21188 34098 21244
rect 34034 21184 34098 21188
rect 34114 21244 34178 21248
rect 34114 21188 34118 21244
rect 34118 21188 34174 21244
rect 34174 21188 34178 21244
rect 34114 21184 34178 21188
rect 55822 21244 55886 21248
rect 55822 21188 55826 21244
rect 55826 21188 55882 21244
rect 55882 21188 55886 21244
rect 55822 21184 55886 21188
rect 55902 21244 55966 21248
rect 55902 21188 55906 21244
rect 55906 21188 55962 21244
rect 55962 21188 55966 21244
rect 55902 21184 55966 21188
rect 55982 21244 56046 21248
rect 55982 21188 55986 21244
rect 55986 21188 56042 21244
rect 56042 21188 56046 21244
rect 55982 21184 56046 21188
rect 56062 21244 56126 21248
rect 56062 21188 56066 21244
rect 56066 21188 56122 21244
rect 56122 21188 56126 21244
rect 56062 21184 56126 21188
rect 77770 21244 77834 21248
rect 77770 21188 77774 21244
rect 77774 21188 77830 21244
rect 77830 21188 77834 21244
rect 77770 21184 77834 21188
rect 77850 21244 77914 21248
rect 77850 21188 77854 21244
rect 77854 21188 77910 21244
rect 77910 21188 77914 21244
rect 77850 21184 77914 21188
rect 77930 21244 77994 21248
rect 77930 21188 77934 21244
rect 77934 21188 77990 21244
rect 77990 21188 77994 21244
rect 77930 21184 77994 21188
rect 78010 21244 78074 21248
rect 78010 21188 78014 21244
rect 78014 21188 78070 21244
rect 78070 21188 78074 21244
rect 78010 21184 78074 21188
rect 22900 20700 22964 20704
rect 22900 20644 22904 20700
rect 22904 20644 22960 20700
rect 22960 20644 22964 20700
rect 22900 20640 22964 20644
rect 22980 20700 23044 20704
rect 22980 20644 22984 20700
rect 22984 20644 23040 20700
rect 23040 20644 23044 20700
rect 22980 20640 23044 20644
rect 23060 20700 23124 20704
rect 23060 20644 23064 20700
rect 23064 20644 23120 20700
rect 23120 20644 23124 20700
rect 23060 20640 23124 20644
rect 23140 20700 23204 20704
rect 23140 20644 23144 20700
rect 23144 20644 23200 20700
rect 23200 20644 23204 20700
rect 23140 20640 23204 20644
rect 44848 20700 44912 20704
rect 44848 20644 44852 20700
rect 44852 20644 44908 20700
rect 44908 20644 44912 20700
rect 44848 20640 44912 20644
rect 44928 20700 44992 20704
rect 44928 20644 44932 20700
rect 44932 20644 44988 20700
rect 44988 20644 44992 20700
rect 44928 20640 44992 20644
rect 45008 20700 45072 20704
rect 45008 20644 45012 20700
rect 45012 20644 45068 20700
rect 45068 20644 45072 20700
rect 45008 20640 45072 20644
rect 45088 20700 45152 20704
rect 45088 20644 45092 20700
rect 45092 20644 45148 20700
rect 45148 20644 45152 20700
rect 45088 20640 45152 20644
rect 66796 20700 66860 20704
rect 66796 20644 66800 20700
rect 66800 20644 66856 20700
rect 66856 20644 66860 20700
rect 66796 20640 66860 20644
rect 66876 20700 66940 20704
rect 66876 20644 66880 20700
rect 66880 20644 66936 20700
rect 66936 20644 66940 20700
rect 66876 20640 66940 20644
rect 66956 20700 67020 20704
rect 66956 20644 66960 20700
rect 66960 20644 67016 20700
rect 67016 20644 67020 20700
rect 66956 20640 67020 20644
rect 67036 20700 67100 20704
rect 67036 20644 67040 20700
rect 67040 20644 67096 20700
rect 67096 20644 67100 20700
rect 67036 20640 67100 20644
rect 11926 20156 11990 20160
rect 11926 20100 11930 20156
rect 11930 20100 11986 20156
rect 11986 20100 11990 20156
rect 11926 20096 11990 20100
rect 12006 20156 12070 20160
rect 12006 20100 12010 20156
rect 12010 20100 12066 20156
rect 12066 20100 12070 20156
rect 12006 20096 12070 20100
rect 12086 20156 12150 20160
rect 12086 20100 12090 20156
rect 12090 20100 12146 20156
rect 12146 20100 12150 20156
rect 12086 20096 12150 20100
rect 12166 20156 12230 20160
rect 12166 20100 12170 20156
rect 12170 20100 12226 20156
rect 12226 20100 12230 20156
rect 12166 20096 12230 20100
rect 33874 20156 33938 20160
rect 33874 20100 33878 20156
rect 33878 20100 33934 20156
rect 33934 20100 33938 20156
rect 33874 20096 33938 20100
rect 33954 20156 34018 20160
rect 33954 20100 33958 20156
rect 33958 20100 34014 20156
rect 34014 20100 34018 20156
rect 33954 20096 34018 20100
rect 34034 20156 34098 20160
rect 34034 20100 34038 20156
rect 34038 20100 34094 20156
rect 34094 20100 34098 20156
rect 34034 20096 34098 20100
rect 34114 20156 34178 20160
rect 34114 20100 34118 20156
rect 34118 20100 34174 20156
rect 34174 20100 34178 20156
rect 34114 20096 34178 20100
rect 55822 20156 55886 20160
rect 55822 20100 55826 20156
rect 55826 20100 55882 20156
rect 55882 20100 55886 20156
rect 55822 20096 55886 20100
rect 55902 20156 55966 20160
rect 55902 20100 55906 20156
rect 55906 20100 55962 20156
rect 55962 20100 55966 20156
rect 55902 20096 55966 20100
rect 55982 20156 56046 20160
rect 55982 20100 55986 20156
rect 55986 20100 56042 20156
rect 56042 20100 56046 20156
rect 55982 20096 56046 20100
rect 56062 20156 56126 20160
rect 56062 20100 56066 20156
rect 56066 20100 56122 20156
rect 56122 20100 56126 20156
rect 56062 20096 56126 20100
rect 77770 20156 77834 20160
rect 77770 20100 77774 20156
rect 77774 20100 77830 20156
rect 77830 20100 77834 20156
rect 77770 20096 77834 20100
rect 77850 20156 77914 20160
rect 77850 20100 77854 20156
rect 77854 20100 77910 20156
rect 77910 20100 77914 20156
rect 77850 20096 77914 20100
rect 77930 20156 77994 20160
rect 77930 20100 77934 20156
rect 77934 20100 77990 20156
rect 77990 20100 77994 20156
rect 77930 20096 77994 20100
rect 78010 20156 78074 20160
rect 78010 20100 78014 20156
rect 78014 20100 78070 20156
rect 78070 20100 78074 20156
rect 78010 20096 78074 20100
rect 22900 19612 22964 19616
rect 22900 19556 22904 19612
rect 22904 19556 22960 19612
rect 22960 19556 22964 19612
rect 22900 19552 22964 19556
rect 22980 19612 23044 19616
rect 22980 19556 22984 19612
rect 22984 19556 23040 19612
rect 23040 19556 23044 19612
rect 22980 19552 23044 19556
rect 23060 19612 23124 19616
rect 23060 19556 23064 19612
rect 23064 19556 23120 19612
rect 23120 19556 23124 19612
rect 23060 19552 23124 19556
rect 23140 19612 23204 19616
rect 23140 19556 23144 19612
rect 23144 19556 23200 19612
rect 23200 19556 23204 19612
rect 23140 19552 23204 19556
rect 44848 19612 44912 19616
rect 44848 19556 44852 19612
rect 44852 19556 44908 19612
rect 44908 19556 44912 19612
rect 44848 19552 44912 19556
rect 44928 19612 44992 19616
rect 44928 19556 44932 19612
rect 44932 19556 44988 19612
rect 44988 19556 44992 19612
rect 44928 19552 44992 19556
rect 45008 19612 45072 19616
rect 45008 19556 45012 19612
rect 45012 19556 45068 19612
rect 45068 19556 45072 19612
rect 45008 19552 45072 19556
rect 45088 19612 45152 19616
rect 45088 19556 45092 19612
rect 45092 19556 45148 19612
rect 45148 19556 45152 19612
rect 45088 19552 45152 19556
rect 66796 19612 66860 19616
rect 66796 19556 66800 19612
rect 66800 19556 66856 19612
rect 66856 19556 66860 19612
rect 66796 19552 66860 19556
rect 66876 19612 66940 19616
rect 66876 19556 66880 19612
rect 66880 19556 66936 19612
rect 66936 19556 66940 19612
rect 66876 19552 66940 19556
rect 66956 19612 67020 19616
rect 66956 19556 66960 19612
rect 66960 19556 67016 19612
rect 67016 19556 67020 19612
rect 66956 19552 67020 19556
rect 67036 19612 67100 19616
rect 67036 19556 67040 19612
rect 67040 19556 67096 19612
rect 67096 19556 67100 19612
rect 67036 19552 67100 19556
rect 11926 19068 11990 19072
rect 11926 19012 11930 19068
rect 11930 19012 11986 19068
rect 11986 19012 11990 19068
rect 11926 19008 11990 19012
rect 12006 19068 12070 19072
rect 12006 19012 12010 19068
rect 12010 19012 12066 19068
rect 12066 19012 12070 19068
rect 12006 19008 12070 19012
rect 12086 19068 12150 19072
rect 12086 19012 12090 19068
rect 12090 19012 12146 19068
rect 12146 19012 12150 19068
rect 12086 19008 12150 19012
rect 12166 19068 12230 19072
rect 12166 19012 12170 19068
rect 12170 19012 12226 19068
rect 12226 19012 12230 19068
rect 12166 19008 12230 19012
rect 33874 19068 33938 19072
rect 33874 19012 33878 19068
rect 33878 19012 33934 19068
rect 33934 19012 33938 19068
rect 33874 19008 33938 19012
rect 33954 19068 34018 19072
rect 33954 19012 33958 19068
rect 33958 19012 34014 19068
rect 34014 19012 34018 19068
rect 33954 19008 34018 19012
rect 34034 19068 34098 19072
rect 34034 19012 34038 19068
rect 34038 19012 34094 19068
rect 34094 19012 34098 19068
rect 34034 19008 34098 19012
rect 34114 19068 34178 19072
rect 34114 19012 34118 19068
rect 34118 19012 34174 19068
rect 34174 19012 34178 19068
rect 34114 19008 34178 19012
rect 55822 19068 55886 19072
rect 55822 19012 55826 19068
rect 55826 19012 55882 19068
rect 55882 19012 55886 19068
rect 55822 19008 55886 19012
rect 55902 19068 55966 19072
rect 55902 19012 55906 19068
rect 55906 19012 55962 19068
rect 55962 19012 55966 19068
rect 55902 19008 55966 19012
rect 55982 19068 56046 19072
rect 55982 19012 55986 19068
rect 55986 19012 56042 19068
rect 56042 19012 56046 19068
rect 55982 19008 56046 19012
rect 56062 19068 56126 19072
rect 56062 19012 56066 19068
rect 56066 19012 56122 19068
rect 56122 19012 56126 19068
rect 56062 19008 56126 19012
rect 77770 19068 77834 19072
rect 77770 19012 77774 19068
rect 77774 19012 77830 19068
rect 77830 19012 77834 19068
rect 77770 19008 77834 19012
rect 77850 19068 77914 19072
rect 77850 19012 77854 19068
rect 77854 19012 77910 19068
rect 77910 19012 77914 19068
rect 77850 19008 77914 19012
rect 77930 19068 77994 19072
rect 77930 19012 77934 19068
rect 77934 19012 77990 19068
rect 77990 19012 77994 19068
rect 77930 19008 77994 19012
rect 78010 19068 78074 19072
rect 78010 19012 78014 19068
rect 78014 19012 78070 19068
rect 78070 19012 78074 19068
rect 78010 19008 78074 19012
rect 22900 18524 22964 18528
rect 22900 18468 22904 18524
rect 22904 18468 22960 18524
rect 22960 18468 22964 18524
rect 22900 18464 22964 18468
rect 22980 18524 23044 18528
rect 22980 18468 22984 18524
rect 22984 18468 23040 18524
rect 23040 18468 23044 18524
rect 22980 18464 23044 18468
rect 23060 18524 23124 18528
rect 23060 18468 23064 18524
rect 23064 18468 23120 18524
rect 23120 18468 23124 18524
rect 23060 18464 23124 18468
rect 23140 18524 23204 18528
rect 23140 18468 23144 18524
rect 23144 18468 23200 18524
rect 23200 18468 23204 18524
rect 23140 18464 23204 18468
rect 44848 18524 44912 18528
rect 44848 18468 44852 18524
rect 44852 18468 44908 18524
rect 44908 18468 44912 18524
rect 44848 18464 44912 18468
rect 44928 18524 44992 18528
rect 44928 18468 44932 18524
rect 44932 18468 44988 18524
rect 44988 18468 44992 18524
rect 44928 18464 44992 18468
rect 45008 18524 45072 18528
rect 45008 18468 45012 18524
rect 45012 18468 45068 18524
rect 45068 18468 45072 18524
rect 45008 18464 45072 18468
rect 45088 18524 45152 18528
rect 45088 18468 45092 18524
rect 45092 18468 45148 18524
rect 45148 18468 45152 18524
rect 45088 18464 45152 18468
rect 66796 18524 66860 18528
rect 66796 18468 66800 18524
rect 66800 18468 66856 18524
rect 66856 18468 66860 18524
rect 66796 18464 66860 18468
rect 66876 18524 66940 18528
rect 66876 18468 66880 18524
rect 66880 18468 66936 18524
rect 66936 18468 66940 18524
rect 66876 18464 66940 18468
rect 66956 18524 67020 18528
rect 66956 18468 66960 18524
rect 66960 18468 67016 18524
rect 67016 18468 67020 18524
rect 66956 18464 67020 18468
rect 67036 18524 67100 18528
rect 67036 18468 67040 18524
rect 67040 18468 67096 18524
rect 67096 18468 67100 18524
rect 67036 18464 67100 18468
rect 56364 18320 56428 18324
rect 56364 18264 56378 18320
rect 56378 18264 56428 18320
rect 56364 18260 56428 18264
rect 11926 17980 11990 17984
rect 11926 17924 11930 17980
rect 11930 17924 11986 17980
rect 11986 17924 11990 17980
rect 11926 17920 11990 17924
rect 12006 17980 12070 17984
rect 12006 17924 12010 17980
rect 12010 17924 12066 17980
rect 12066 17924 12070 17980
rect 12006 17920 12070 17924
rect 12086 17980 12150 17984
rect 12086 17924 12090 17980
rect 12090 17924 12146 17980
rect 12146 17924 12150 17980
rect 12086 17920 12150 17924
rect 12166 17980 12230 17984
rect 12166 17924 12170 17980
rect 12170 17924 12226 17980
rect 12226 17924 12230 17980
rect 12166 17920 12230 17924
rect 33874 17980 33938 17984
rect 33874 17924 33878 17980
rect 33878 17924 33934 17980
rect 33934 17924 33938 17980
rect 33874 17920 33938 17924
rect 33954 17980 34018 17984
rect 33954 17924 33958 17980
rect 33958 17924 34014 17980
rect 34014 17924 34018 17980
rect 33954 17920 34018 17924
rect 34034 17980 34098 17984
rect 34034 17924 34038 17980
rect 34038 17924 34094 17980
rect 34094 17924 34098 17980
rect 34034 17920 34098 17924
rect 34114 17980 34178 17984
rect 34114 17924 34118 17980
rect 34118 17924 34174 17980
rect 34174 17924 34178 17980
rect 34114 17920 34178 17924
rect 55822 17980 55886 17984
rect 55822 17924 55826 17980
rect 55826 17924 55882 17980
rect 55882 17924 55886 17980
rect 55822 17920 55886 17924
rect 55902 17980 55966 17984
rect 55902 17924 55906 17980
rect 55906 17924 55962 17980
rect 55962 17924 55966 17980
rect 55902 17920 55966 17924
rect 55982 17980 56046 17984
rect 55982 17924 55986 17980
rect 55986 17924 56042 17980
rect 56042 17924 56046 17980
rect 55982 17920 56046 17924
rect 56062 17980 56126 17984
rect 56062 17924 56066 17980
rect 56066 17924 56122 17980
rect 56122 17924 56126 17980
rect 56062 17920 56126 17924
rect 77770 17980 77834 17984
rect 77770 17924 77774 17980
rect 77774 17924 77830 17980
rect 77830 17924 77834 17980
rect 77770 17920 77834 17924
rect 77850 17980 77914 17984
rect 77850 17924 77854 17980
rect 77854 17924 77910 17980
rect 77910 17924 77914 17980
rect 77850 17920 77914 17924
rect 77930 17980 77994 17984
rect 77930 17924 77934 17980
rect 77934 17924 77990 17980
rect 77990 17924 77994 17980
rect 77930 17920 77994 17924
rect 78010 17980 78074 17984
rect 78010 17924 78014 17980
rect 78014 17924 78070 17980
rect 78070 17924 78074 17980
rect 78010 17920 78074 17924
rect 22900 17436 22964 17440
rect 22900 17380 22904 17436
rect 22904 17380 22960 17436
rect 22960 17380 22964 17436
rect 22900 17376 22964 17380
rect 22980 17436 23044 17440
rect 22980 17380 22984 17436
rect 22984 17380 23040 17436
rect 23040 17380 23044 17436
rect 22980 17376 23044 17380
rect 23060 17436 23124 17440
rect 23060 17380 23064 17436
rect 23064 17380 23120 17436
rect 23120 17380 23124 17436
rect 23060 17376 23124 17380
rect 23140 17436 23204 17440
rect 23140 17380 23144 17436
rect 23144 17380 23200 17436
rect 23200 17380 23204 17436
rect 23140 17376 23204 17380
rect 44848 17436 44912 17440
rect 44848 17380 44852 17436
rect 44852 17380 44908 17436
rect 44908 17380 44912 17436
rect 44848 17376 44912 17380
rect 44928 17436 44992 17440
rect 44928 17380 44932 17436
rect 44932 17380 44988 17436
rect 44988 17380 44992 17436
rect 44928 17376 44992 17380
rect 45008 17436 45072 17440
rect 45008 17380 45012 17436
rect 45012 17380 45068 17436
rect 45068 17380 45072 17436
rect 45008 17376 45072 17380
rect 45088 17436 45152 17440
rect 45088 17380 45092 17436
rect 45092 17380 45148 17436
rect 45148 17380 45152 17436
rect 45088 17376 45152 17380
rect 66796 17436 66860 17440
rect 66796 17380 66800 17436
rect 66800 17380 66856 17436
rect 66856 17380 66860 17436
rect 66796 17376 66860 17380
rect 66876 17436 66940 17440
rect 66876 17380 66880 17436
rect 66880 17380 66936 17436
rect 66936 17380 66940 17436
rect 66876 17376 66940 17380
rect 66956 17436 67020 17440
rect 66956 17380 66960 17436
rect 66960 17380 67016 17436
rect 67016 17380 67020 17436
rect 66956 17376 67020 17380
rect 67036 17436 67100 17440
rect 67036 17380 67040 17436
rect 67040 17380 67096 17436
rect 67096 17380 67100 17436
rect 67036 17376 67100 17380
rect 11926 16892 11990 16896
rect 11926 16836 11930 16892
rect 11930 16836 11986 16892
rect 11986 16836 11990 16892
rect 11926 16832 11990 16836
rect 12006 16892 12070 16896
rect 12006 16836 12010 16892
rect 12010 16836 12066 16892
rect 12066 16836 12070 16892
rect 12006 16832 12070 16836
rect 12086 16892 12150 16896
rect 12086 16836 12090 16892
rect 12090 16836 12146 16892
rect 12146 16836 12150 16892
rect 12086 16832 12150 16836
rect 12166 16892 12230 16896
rect 12166 16836 12170 16892
rect 12170 16836 12226 16892
rect 12226 16836 12230 16892
rect 12166 16832 12230 16836
rect 33874 16892 33938 16896
rect 33874 16836 33878 16892
rect 33878 16836 33934 16892
rect 33934 16836 33938 16892
rect 33874 16832 33938 16836
rect 33954 16892 34018 16896
rect 33954 16836 33958 16892
rect 33958 16836 34014 16892
rect 34014 16836 34018 16892
rect 33954 16832 34018 16836
rect 34034 16892 34098 16896
rect 34034 16836 34038 16892
rect 34038 16836 34094 16892
rect 34094 16836 34098 16892
rect 34034 16832 34098 16836
rect 34114 16892 34178 16896
rect 34114 16836 34118 16892
rect 34118 16836 34174 16892
rect 34174 16836 34178 16892
rect 34114 16832 34178 16836
rect 55822 16892 55886 16896
rect 55822 16836 55826 16892
rect 55826 16836 55882 16892
rect 55882 16836 55886 16892
rect 55822 16832 55886 16836
rect 55902 16892 55966 16896
rect 55902 16836 55906 16892
rect 55906 16836 55962 16892
rect 55962 16836 55966 16892
rect 55902 16832 55966 16836
rect 55982 16892 56046 16896
rect 55982 16836 55986 16892
rect 55986 16836 56042 16892
rect 56042 16836 56046 16892
rect 55982 16832 56046 16836
rect 56062 16892 56126 16896
rect 56062 16836 56066 16892
rect 56066 16836 56122 16892
rect 56122 16836 56126 16892
rect 56062 16832 56126 16836
rect 77770 16892 77834 16896
rect 77770 16836 77774 16892
rect 77774 16836 77830 16892
rect 77830 16836 77834 16892
rect 77770 16832 77834 16836
rect 77850 16892 77914 16896
rect 77850 16836 77854 16892
rect 77854 16836 77910 16892
rect 77910 16836 77914 16892
rect 77850 16832 77914 16836
rect 77930 16892 77994 16896
rect 77930 16836 77934 16892
rect 77934 16836 77990 16892
rect 77990 16836 77994 16892
rect 77930 16832 77994 16836
rect 78010 16892 78074 16896
rect 78010 16836 78014 16892
rect 78014 16836 78070 16892
rect 78070 16836 78074 16892
rect 78010 16832 78074 16836
rect 22900 16348 22964 16352
rect 22900 16292 22904 16348
rect 22904 16292 22960 16348
rect 22960 16292 22964 16348
rect 22900 16288 22964 16292
rect 22980 16348 23044 16352
rect 22980 16292 22984 16348
rect 22984 16292 23040 16348
rect 23040 16292 23044 16348
rect 22980 16288 23044 16292
rect 23060 16348 23124 16352
rect 23060 16292 23064 16348
rect 23064 16292 23120 16348
rect 23120 16292 23124 16348
rect 23060 16288 23124 16292
rect 23140 16348 23204 16352
rect 23140 16292 23144 16348
rect 23144 16292 23200 16348
rect 23200 16292 23204 16348
rect 23140 16288 23204 16292
rect 44848 16348 44912 16352
rect 44848 16292 44852 16348
rect 44852 16292 44908 16348
rect 44908 16292 44912 16348
rect 44848 16288 44912 16292
rect 44928 16348 44992 16352
rect 44928 16292 44932 16348
rect 44932 16292 44988 16348
rect 44988 16292 44992 16348
rect 44928 16288 44992 16292
rect 45008 16348 45072 16352
rect 45008 16292 45012 16348
rect 45012 16292 45068 16348
rect 45068 16292 45072 16348
rect 45008 16288 45072 16292
rect 45088 16348 45152 16352
rect 45088 16292 45092 16348
rect 45092 16292 45148 16348
rect 45148 16292 45152 16348
rect 45088 16288 45152 16292
rect 66796 16348 66860 16352
rect 66796 16292 66800 16348
rect 66800 16292 66856 16348
rect 66856 16292 66860 16348
rect 66796 16288 66860 16292
rect 66876 16348 66940 16352
rect 66876 16292 66880 16348
rect 66880 16292 66936 16348
rect 66936 16292 66940 16348
rect 66876 16288 66940 16292
rect 66956 16348 67020 16352
rect 66956 16292 66960 16348
rect 66960 16292 67016 16348
rect 67016 16292 67020 16348
rect 66956 16288 67020 16292
rect 67036 16348 67100 16352
rect 67036 16292 67040 16348
rect 67040 16292 67096 16348
rect 67096 16292 67100 16348
rect 67036 16288 67100 16292
rect 55628 16084 55692 16148
rect 11926 15804 11990 15808
rect 11926 15748 11930 15804
rect 11930 15748 11986 15804
rect 11986 15748 11990 15804
rect 11926 15744 11990 15748
rect 12006 15804 12070 15808
rect 12006 15748 12010 15804
rect 12010 15748 12066 15804
rect 12066 15748 12070 15804
rect 12006 15744 12070 15748
rect 12086 15804 12150 15808
rect 12086 15748 12090 15804
rect 12090 15748 12146 15804
rect 12146 15748 12150 15804
rect 12086 15744 12150 15748
rect 12166 15804 12230 15808
rect 12166 15748 12170 15804
rect 12170 15748 12226 15804
rect 12226 15748 12230 15804
rect 12166 15744 12230 15748
rect 33874 15804 33938 15808
rect 33874 15748 33878 15804
rect 33878 15748 33934 15804
rect 33934 15748 33938 15804
rect 33874 15744 33938 15748
rect 33954 15804 34018 15808
rect 33954 15748 33958 15804
rect 33958 15748 34014 15804
rect 34014 15748 34018 15804
rect 33954 15744 34018 15748
rect 34034 15804 34098 15808
rect 34034 15748 34038 15804
rect 34038 15748 34094 15804
rect 34094 15748 34098 15804
rect 34034 15744 34098 15748
rect 34114 15804 34178 15808
rect 34114 15748 34118 15804
rect 34118 15748 34174 15804
rect 34174 15748 34178 15804
rect 34114 15744 34178 15748
rect 55822 15804 55886 15808
rect 55822 15748 55826 15804
rect 55826 15748 55882 15804
rect 55882 15748 55886 15804
rect 55822 15744 55886 15748
rect 55902 15804 55966 15808
rect 55902 15748 55906 15804
rect 55906 15748 55962 15804
rect 55962 15748 55966 15804
rect 55902 15744 55966 15748
rect 55982 15804 56046 15808
rect 55982 15748 55986 15804
rect 55986 15748 56042 15804
rect 56042 15748 56046 15804
rect 55982 15744 56046 15748
rect 56062 15804 56126 15808
rect 56062 15748 56066 15804
rect 56066 15748 56122 15804
rect 56122 15748 56126 15804
rect 56062 15744 56126 15748
rect 77770 15804 77834 15808
rect 77770 15748 77774 15804
rect 77774 15748 77830 15804
rect 77830 15748 77834 15804
rect 77770 15744 77834 15748
rect 77850 15804 77914 15808
rect 77850 15748 77854 15804
rect 77854 15748 77910 15804
rect 77910 15748 77914 15804
rect 77850 15744 77914 15748
rect 77930 15804 77994 15808
rect 77930 15748 77934 15804
rect 77934 15748 77990 15804
rect 77990 15748 77994 15804
rect 77930 15744 77994 15748
rect 78010 15804 78074 15808
rect 78010 15748 78014 15804
rect 78014 15748 78070 15804
rect 78070 15748 78074 15804
rect 78010 15744 78074 15748
rect 28028 15540 28092 15604
rect 22900 15260 22964 15264
rect 22900 15204 22904 15260
rect 22904 15204 22960 15260
rect 22960 15204 22964 15260
rect 22900 15200 22964 15204
rect 22980 15260 23044 15264
rect 22980 15204 22984 15260
rect 22984 15204 23040 15260
rect 23040 15204 23044 15260
rect 22980 15200 23044 15204
rect 23060 15260 23124 15264
rect 23060 15204 23064 15260
rect 23064 15204 23120 15260
rect 23120 15204 23124 15260
rect 23060 15200 23124 15204
rect 23140 15260 23204 15264
rect 23140 15204 23144 15260
rect 23144 15204 23200 15260
rect 23200 15204 23204 15260
rect 23140 15200 23204 15204
rect 44848 15260 44912 15264
rect 44848 15204 44852 15260
rect 44852 15204 44908 15260
rect 44908 15204 44912 15260
rect 44848 15200 44912 15204
rect 44928 15260 44992 15264
rect 44928 15204 44932 15260
rect 44932 15204 44988 15260
rect 44988 15204 44992 15260
rect 44928 15200 44992 15204
rect 45008 15260 45072 15264
rect 45008 15204 45012 15260
rect 45012 15204 45068 15260
rect 45068 15204 45072 15260
rect 45008 15200 45072 15204
rect 45088 15260 45152 15264
rect 45088 15204 45092 15260
rect 45092 15204 45148 15260
rect 45148 15204 45152 15260
rect 45088 15200 45152 15204
rect 66796 15260 66860 15264
rect 66796 15204 66800 15260
rect 66800 15204 66856 15260
rect 66856 15204 66860 15260
rect 66796 15200 66860 15204
rect 66876 15260 66940 15264
rect 66876 15204 66880 15260
rect 66880 15204 66936 15260
rect 66936 15204 66940 15260
rect 66876 15200 66940 15204
rect 66956 15260 67020 15264
rect 66956 15204 66960 15260
rect 66960 15204 67016 15260
rect 67016 15204 67020 15260
rect 66956 15200 67020 15204
rect 67036 15260 67100 15264
rect 67036 15204 67040 15260
rect 67040 15204 67096 15260
rect 67096 15204 67100 15260
rect 67036 15200 67100 15204
rect 27476 15132 27540 15196
rect 11926 14716 11990 14720
rect 11926 14660 11930 14716
rect 11930 14660 11986 14716
rect 11986 14660 11990 14716
rect 11926 14656 11990 14660
rect 12006 14716 12070 14720
rect 12006 14660 12010 14716
rect 12010 14660 12066 14716
rect 12066 14660 12070 14716
rect 12006 14656 12070 14660
rect 12086 14716 12150 14720
rect 12086 14660 12090 14716
rect 12090 14660 12146 14716
rect 12146 14660 12150 14716
rect 12086 14656 12150 14660
rect 12166 14716 12230 14720
rect 12166 14660 12170 14716
rect 12170 14660 12226 14716
rect 12226 14660 12230 14716
rect 12166 14656 12230 14660
rect 33874 14716 33938 14720
rect 33874 14660 33878 14716
rect 33878 14660 33934 14716
rect 33934 14660 33938 14716
rect 33874 14656 33938 14660
rect 33954 14716 34018 14720
rect 33954 14660 33958 14716
rect 33958 14660 34014 14716
rect 34014 14660 34018 14716
rect 33954 14656 34018 14660
rect 34034 14716 34098 14720
rect 34034 14660 34038 14716
rect 34038 14660 34094 14716
rect 34094 14660 34098 14716
rect 34034 14656 34098 14660
rect 34114 14716 34178 14720
rect 34114 14660 34118 14716
rect 34118 14660 34174 14716
rect 34174 14660 34178 14716
rect 34114 14656 34178 14660
rect 56916 14784 56980 14788
rect 56916 14728 56930 14784
rect 56930 14728 56980 14784
rect 56916 14724 56980 14728
rect 55822 14716 55886 14720
rect 55822 14660 55826 14716
rect 55826 14660 55882 14716
rect 55882 14660 55886 14716
rect 55822 14656 55886 14660
rect 55902 14716 55966 14720
rect 55902 14660 55906 14716
rect 55906 14660 55962 14716
rect 55962 14660 55966 14716
rect 55902 14656 55966 14660
rect 55982 14716 56046 14720
rect 55982 14660 55986 14716
rect 55986 14660 56042 14716
rect 56042 14660 56046 14716
rect 55982 14656 56046 14660
rect 56062 14716 56126 14720
rect 56062 14660 56066 14716
rect 56066 14660 56122 14716
rect 56122 14660 56126 14716
rect 56062 14656 56126 14660
rect 77770 14716 77834 14720
rect 77770 14660 77774 14716
rect 77774 14660 77830 14716
rect 77830 14660 77834 14716
rect 77770 14656 77834 14660
rect 77850 14716 77914 14720
rect 77850 14660 77854 14716
rect 77854 14660 77910 14716
rect 77910 14660 77914 14716
rect 77850 14656 77914 14660
rect 77930 14716 77994 14720
rect 77930 14660 77934 14716
rect 77934 14660 77990 14716
rect 77990 14660 77994 14716
rect 77930 14656 77994 14660
rect 78010 14716 78074 14720
rect 78010 14660 78014 14716
rect 78014 14660 78070 14716
rect 78070 14660 78074 14716
rect 78010 14656 78074 14660
rect 63908 14316 63972 14380
rect 22900 14172 22964 14176
rect 22900 14116 22904 14172
rect 22904 14116 22960 14172
rect 22960 14116 22964 14172
rect 22900 14112 22964 14116
rect 22980 14172 23044 14176
rect 22980 14116 22984 14172
rect 22984 14116 23040 14172
rect 23040 14116 23044 14172
rect 22980 14112 23044 14116
rect 23060 14172 23124 14176
rect 23060 14116 23064 14172
rect 23064 14116 23120 14172
rect 23120 14116 23124 14172
rect 23060 14112 23124 14116
rect 23140 14172 23204 14176
rect 23140 14116 23144 14172
rect 23144 14116 23200 14172
rect 23200 14116 23204 14172
rect 23140 14112 23204 14116
rect 44848 14172 44912 14176
rect 44848 14116 44852 14172
rect 44852 14116 44908 14172
rect 44908 14116 44912 14172
rect 44848 14112 44912 14116
rect 44928 14172 44992 14176
rect 44928 14116 44932 14172
rect 44932 14116 44988 14172
rect 44988 14116 44992 14172
rect 44928 14112 44992 14116
rect 45008 14172 45072 14176
rect 45008 14116 45012 14172
rect 45012 14116 45068 14172
rect 45068 14116 45072 14172
rect 45008 14112 45072 14116
rect 45088 14172 45152 14176
rect 45088 14116 45092 14172
rect 45092 14116 45148 14172
rect 45148 14116 45152 14172
rect 45088 14112 45152 14116
rect 66796 14172 66860 14176
rect 66796 14116 66800 14172
rect 66800 14116 66856 14172
rect 66856 14116 66860 14172
rect 66796 14112 66860 14116
rect 66876 14172 66940 14176
rect 66876 14116 66880 14172
rect 66880 14116 66936 14172
rect 66936 14116 66940 14172
rect 66876 14112 66940 14116
rect 66956 14172 67020 14176
rect 66956 14116 66960 14172
rect 66960 14116 67016 14172
rect 67016 14116 67020 14172
rect 66956 14112 67020 14116
rect 67036 14172 67100 14176
rect 67036 14116 67040 14172
rect 67040 14116 67096 14172
rect 67096 14116 67100 14172
rect 67036 14112 67100 14116
rect 11926 13628 11990 13632
rect 11926 13572 11930 13628
rect 11930 13572 11986 13628
rect 11986 13572 11990 13628
rect 11926 13568 11990 13572
rect 12006 13628 12070 13632
rect 12006 13572 12010 13628
rect 12010 13572 12066 13628
rect 12066 13572 12070 13628
rect 12006 13568 12070 13572
rect 12086 13628 12150 13632
rect 12086 13572 12090 13628
rect 12090 13572 12146 13628
rect 12146 13572 12150 13628
rect 12086 13568 12150 13572
rect 12166 13628 12230 13632
rect 12166 13572 12170 13628
rect 12170 13572 12226 13628
rect 12226 13572 12230 13628
rect 12166 13568 12230 13572
rect 33874 13628 33938 13632
rect 33874 13572 33878 13628
rect 33878 13572 33934 13628
rect 33934 13572 33938 13628
rect 33874 13568 33938 13572
rect 33954 13628 34018 13632
rect 33954 13572 33958 13628
rect 33958 13572 34014 13628
rect 34014 13572 34018 13628
rect 33954 13568 34018 13572
rect 34034 13628 34098 13632
rect 34034 13572 34038 13628
rect 34038 13572 34094 13628
rect 34094 13572 34098 13628
rect 34034 13568 34098 13572
rect 34114 13628 34178 13632
rect 34114 13572 34118 13628
rect 34118 13572 34174 13628
rect 34174 13572 34178 13628
rect 34114 13568 34178 13572
rect 55822 13628 55886 13632
rect 55822 13572 55826 13628
rect 55826 13572 55882 13628
rect 55882 13572 55886 13628
rect 55822 13568 55886 13572
rect 55902 13628 55966 13632
rect 55902 13572 55906 13628
rect 55906 13572 55962 13628
rect 55962 13572 55966 13628
rect 55902 13568 55966 13572
rect 55982 13628 56046 13632
rect 55982 13572 55986 13628
rect 55986 13572 56042 13628
rect 56042 13572 56046 13628
rect 55982 13568 56046 13572
rect 56062 13628 56126 13632
rect 56062 13572 56066 13628
rect 56066 13572 56122 13628
rect 56122 13572 56126 13628
rect 56062 13568 56126 13572
rect 77770 13628 77834 13632
rect 77770 13572 77774 13628
rect 77774 13572 77830 13628
rect 77830 13572 77834 13628
rect 77770 13568 77834 13572
rect 77850 13628 77914 13632
rect 77850 13572 77854 13628
rect 77854 13572 77910 13628
rect 77910 13572 77914 13628
rect 77850 13568 77914 13572
rect 77930 13628 77994 13632
rect 77930 13572 77934 13628
rect 77934 13572 77990 13628
rect 77990 13572 77994 13628
rect 77930 13568 77994 13572
rect 78010 13628 78074 13632
rect 78010 13572 78014 13628
rect 78014 13572 78070 13628
rect 78070 13572 78074 13628
rect 78010 13568 78074 13572
rect 55628 13500 55692 13564
rect 22900 13084 22964 13088
rect 22900 13028 22904 13084
rect 22904 13028 22960 13084
rect 22960 13028 22964 13084
rect 22900 13024 22964 13028
rect 22980 13084 23044 13088
rect 22980 13028 22984 13084
rect 22984 13028 23040 13084
rect 23040 13028 23044 13084
rect 22980 13024 23044 13028
rect 23060 13084 23124 13088
rect 23060 13028 23064 13084
rect 23064 13028 23120 13084
rect 23120 13028 23124 13084
rect 23060 13024 23124 13028
rect 23140 13084 23204 13088
rect 23140 13028 23144 13084
rect 23144 13028 23200 13084
rect 23200 13028 23204 13084
rect 23140 13024 23204 13028
rect 44848 13084 44912 13088
rect 44848 13028 44852 13084
rect 44852 13028 44908 13084
rect 44908 13028 44912 13084
rect 44848 13024 44912 13028
rect 44928 13084 44992 13088
rect 44928 13028 44932 13084
rect 44932 13028 44988 13084
rect 44988 13028 44992 13084
rect 44928 13024 44992 13028
rect 45008 13084 45072 13088
rect 45008 13028 45012 13084
rect 45012 13028 45068 13084
rect 45068 13028 45072 13084
rect 45008 13024 45072 13028
rect 45088 13084 45152 13088
rect 45088 13028 45092 13084
rect 45092 13028 45148 13084
rect 45148 13028 45152 13084
rect 45088 13024 45152 13028
rect 26556 12880 26620 12884
rect 26556 12824 26570 12880
rect 26570 12824 26620 12880
rect 26556 12820 26620 12824
rect 66796 13084 66860 13088
rect 66796 13028 66800 13084
rect 66800 13028 66856 13084
rect 66856 13028 66860 13084
rect 66796 13024 66860 13028
rect 66876 13084 66940 13088
rect 66876 13028 66880 13084
rect 66880 13028 66936 13084
rect 66936 13028 66940 13084
rect 66876 13024 66940 13028
rect 66956 13084 67020 13088
rect 66956 13028 66960 13084
rect 66960 13028 67016 13084
rect 67016 13028 67020 13084
rect 66956 13024 67020 13028
rect 67036 13084 67100 13088
rect 67036 13028 67040 13084
rect 67040 13028 67096 13084
rect 67096 13028 67100 13084
rect 67036 13024 67100 13028
rect 64276 12548 64340 12612
rect 11926 12540 11990 12544
rect 11926 12484 11930 12540
rect 11930 12484 11986 12540
rect 11986 12484 11990 12540
rect 11926 12480 11990 12484
rect 12006 12540 12070 12544
rect 12006 12484 12010 12540
rect 12010 12484 12066 12540
rect 12066 12484 12070 12540
rect 12006 12480 12070 12484
rect 12086 12540 12150 12544
rect 12086 12484 12090 12540
rect 12090 12484 12146 12540
rect 12146 12484 12150 12540
rect 12086 12480 12150 12484
rect 12166 12540 12230 12544
rect 12166 12484 12170 12540
rect 12170 12484 12226 12540
rect 12226 12484 12230 12540
rect 12166 12480 12230 12484
rect 33874 12540 33938 12544
rect 33874 12484 33878 12540
rect 33878 12484 33934 12540
rect 33934 12484 33938 12540
rect 33874 12480 33938 12484
rect 33954 12540 34018 12544
rect 33954 12484 33958 12540
rect 33958 12484 34014 12540
rect 34014 12484 34018 12540
rect 33954 12480 34018 12484
rect 34034 12540 34098 12544
rect 34034 12484 34038 12540
rect 34038 12484 34094 12540
rect 34094 12484 34098 12540
rect 34034 12480 34098 12484
rect 34114 12540 34178 12544
rect 34114 12484 34118 12540
rect 34118 12484 34174 12540
rect 34174 12484 34178 12540
rect 34114 12480 34178 12484
rect 55822 12540 55886 12544
rect 55822 12484 55826 12540
rect 55826 12484 55882 12540
rect 55882 12484 55886 12540
rect 55822 12480 55886 12484
rect 55902 12540 55966 12544
rect 55902 12484 55906 12540
rect 55906 12484 55962 12540
rect 55962 12484 55966 12540
rect 55902 12480 55966 12484
rect 55982 12540 56046 12544
rect 55982 12484 55986 12540
rect 55986 12484 56042 12540
rect 56042 12484 56046 12540
rect 55982 12480 56046 12484
rect 56062 12540 56126 12544
rect 56062 12484 56066 12540
rect 56066 12484 56122 12540
rect 56122 12484 56126 12540
rect 56062 12480 56126 12484
rect 77770 12540 77834 12544
rect 77770 12484 77774 12540
rect 77774 12484 77830 12540
rect 77830 12484 77834 12540
rect 77770 12480 77834 12484
rect 77850 12540 77914 12544
rect 77850 12484 77854 12540
rect 77854 12484 77910 12540
rect 77910 12484 77914 12540
rect 77850 12480 77914 12484
rect 77930 12540 77994 12544
rect 77930 12484 77934 12540
rect 77934 12484 77990 12540
rect 77990 12484 77994 12540
rect 77930 12480 77994 12484
rect 78010 12540 78074 12544
rect 78010 12484 78014 12540
rect 78014 12484 78070 12540
rect 78070 12484 78074 12540
rect 78010 12480 78074 12484
rect 63724 12472 63788 12476
rect 63724 12416 63738 12472
rect 63738 12416 63788 12472
rect 63724 12412 63788 12416
rect 22900 11996 22964 12000
rect 22900 11940 22904 11996
rect 22904 11940 22960 11996
rect 22960 11940 22964 11996
rect 22900 11936 22964 11940
rect 22980 11996 23044 12000
rect 22980 11940 22984 11996
rect 22984 11940 23040 11996
rect 23040 11940 23044 11996
rect 22980 11936 23044 11940
rect 23060 11996 23124 12000
rect 23060 11940 23064 11996
rect 23064 11940 23120 11996
rect 23120 11940 23124 11996
rect 23060 11936 23124 11940
rect 23140 11996 23204 12000
rect 23140 11940 23144 11996
rect 23144 11940 23200 11996
rect 23200 11940 23204 11996
rect 23140 11936 23204 11940
rect 44848 11996 44912 12000
rect 44848 11940 44852 11996
rect 44852 11940 44908 11996
rect 44908 11940 44912 11996
rect 44848 11936 44912 11940
rect 44928 11996 44992 12000
rect 44928 11940 44932 11996
rect 44932 11940 44988 11996
rect 44988 11940 44992 11996
rect 44928 11936 44992 11940
rect 45008 11996 45072 12000
rect 45008 11940 45012 11996
rect 45012 11940 45068 11996
rect 45068 11940 45072 11996
rect 45008 11936 45072 11940
rect 45088 11996 45152 12000
rect 45088 11940 45092 11996
rect 45092 11940 45148 11996
rect 45148 11940 45152 11996
rect 45088 11936 45152 11940
rect 66796 11996 66860 12000
rect 66796 11940 66800 11996
rect 66800 11940 66856 11996
rect 66856 11940 66860 11996
rect 66796 11936 66860 11940
rect 66876 11996 66940 12000
rect 66876 11940 66880 11996
rect 66880 11940 66936 11996
rect 66936 11940 66940 11996
rect 66876 11936 66940 11940
rect 66956 11996 67020 12000
rect 66956 11940 66960 11996
rect 66960 11940 67016 11996
rect 67016 11940 67020 11996
rect 66956 11936 67020 11940
rect 67036 11996 67100 12000
rect 67036 11940 67040 11996
rect 67040 11940 67096 11996
rect 67096 11940 67100 11996
rect 67036 11936 67100 11940
rect 63724 11928 63788 11932
rect 63724 11872 63774 11928
rect 63774 11872 63788 11928
rect 63724 11868 63788 11872
rect 60964 11732 61028 11796
rect 56364 11520 56428 11524
rect 56364 11464 56414 11520
rect 56414 11464 56428 11520
rect 56364 11460 56428 11464
rect 63908 11460 63972 11524
rect 11926 11452 11990 11456
rect 11926 11396 11930 11452
rect 11930 11396 11986 11452
rect 11986 11396 11990 11452
rect 11926 11392 11990 11396
rect 12006 11452 12070 11456
rect 12006 11396 12010 11452
rect 12010 11396 12066 11452
rect 12066 11396 12070 11452
rect 12006 11392 12070 11396
rect 12086 11452 12150 11456
rect 12086 11396 12090 11452
rect 12090 11396 12146 11452
rect 12146 11396 12150 11452
rect 12086 11392 12150 11396
rect 12166 11452 12230 11456
rect 12166 11396 12170 11452
rect 12170 11396 12226 11452
rect 12226 11396 12230 11452
rect 12166 11392 12230 11396
rect 33874 11452 33938 11456
rect 33874 11396 33878 11452
rect 33878 11396 33934 11452
rect 33934 11396 33938 11452
rect 33874 11392 33938 11396
rect 33954 11452 34018 11456
rect 33954 11396 33958 11452
rect 33958 11396 34014 11452
rect 34014 11396 34018 11452
rect 33954 11392 34018 11396
rect 34034 11452 34098 11456
rect 34034 11396 34038 11452
rect 34038 11396 34094 11452
rect 34094 11396 34098 11452
rect 34034 11392 34098 11396
rect 34114 11452 34178 11456
rect 34114 11396 34118 11452
rect 34118 11396 34174 11452
rect 34174 11396 34178 11452
rect 34114 11392 34178 11396
rect 55822 11452 55886 11456
rect 55822 11396 55826 11452
rect 55826 11396 55882 11452
rect 55882 11396 55886 11452
rect 55822 11392 55886 11396
rect 55902 11452 55966 11456
rect 55902 11396 55906 11452
rect 55906 11396 55962 11452
rect 55962 11396 55966 11452
rect 55902 11392 55966 11396
rect 55982 11452 56046 11456
rect 55982 11396 55986 11452
rect 55986 11396 56042 11452
rect 56042 11396 56046 11452
rect 55982 11392 56046 11396
rect 56062 11452 56126 11456
rect 56062 11396 56066 11452
rect 56066 11396 56122 11452
rect 56122 11396 56126 11452
rect 56062 11392 56126 11396
rect 60780 11324 60844 11388
rect 60964 11324 61028 11388
rect 77770 11452 77834 11456
rect 77770 11396 77774 11452
rect 77774 11396 77830 11452
rect 77830 11396 77834 11452
rect 77770 11392 77834 11396
rect 77850 11452 77914 11456
rect 77850 11396 77854 11452
rect 77854 11396 77910 11452
rect 77910 11396 77914 11452
rect 77850 11392 77914 11396
rect 77930 11452 77994 11456
rect 77930 11396 77934 11452
rect 77934 11396 77990 11452
rect 77990 11396 77994 11452
rect 77930 11392 77994 11396
rect 78010 11452 78074 11456
rect 78010 11396 78014 11452
rect 78014 11396 78070 11452
rect 78070 11396 78074 11452
rect 78010 11392 78074 11396
rect 64276 11248 64340 11252
rect 64276 11192 64326 11248
rect 64326 11192 64340 11248
rect 64276 11188 64340 11192
rect 60780 11052 60844 11116
rect 60964 11052 61028 11116
rect 22900 10908 22964 10912
rect 22900 10852 22904 10908
rect 22904 10852 22960 10908
rect 22960 10852 22964 10908
rect 22900 10848 22964 10852
rect 22980 10908 23044 10912
rect 22980 10852 22984 10908
rect 22984 10852 23040 10908
rect 23040 10852 23044 10908
rect 22980 10848 23044 10852
rect 23060 10908 23124 10912
rect 23060 10852 23064 10908
rect 23064 10852 23120 10908
rect 23120 10852 23124 10908
rect 23060 10848 23124 10852
rect 23140 10908 23204 10912
rect 23140 10852 23144 10908
rect 23144 10852 23200 10908
rect 23200 10852 23204 10908
rect 23140 10848 23204 10852
rect 44848 10908 44912 10912
rect 44848 10852 44852 10908
rect 44852 10852 44908 10908
rect 44908 10852 44912 10908
rect 44848 10848 44912 10852
rect 44928 10908 44992 10912
rect 44928 10852 44932 10908
rect 44932 10852 44988 10908
rect 44988 10852 44992 10908
rect 44928 10848 44992 10852
rect 45008 10908 45072 10912
rect 45008 10852 45012 10908
rect 45012 10852 45068 10908
rect 45068 10852 45072 10908
rect 45008 10848 45072 10852
rect 45088 10908 45152 10912
rect 45088 10852 45092 10908
rect 45092 10852 45148 10908
rect 45148 10852 45152 10908
rect 45088 10848 45152 10852
rect 66796 10908 66860 10912
rect 66796 10852 66800 10908
rect 66800 10852 66856 10908
rect 66856 10852 66860 10908
rect 66796 10848 66860 10852
rect 66876 10908 66940 10912
rect 66876 10852 66880 10908
rect 66880 10852 66936 10908
rect 66936 10852 66940 10908
rect 66876 10848 66940 10852
rect 66956 10908 67020 10912
rect 66956 10852 66960 10908
rect 66960 10852 67016 10908
rect 67016 10852 67020 10908
rect 66956 10848 67020 10852
rect 67036 10908 67100 10912
rect 67036 10852 67040 10908
rect 67040 10852 67096 10908
rect 67096 10852 67100 10908
rect 67036 10848 67100 10852
rect 60780 10508 60844 10572
rect 11926 10364 11990 10368
rect 11926 10308 11930 10364
rect 11930 10308 11986 10364
rect 11986 10308 11990 10364
rect 11926 10304 11990 10308
rect 12006 10364 12070 10368
rect 12006 10308 12010 10364
rect 12010 10308 12066 10364
rect 12066 10308 12070 10364
rect 12006 10304 12070 10308
rect 12086 10364 12150 10368
rect 12086 10308 12090 10364
rect 12090 10308 12146 10364
rect 12146 10308 12150 10364
rect 12086 10304 12150 10308
rect 12166 10364 12230 10368
rect 12166 10308 12170 10364
rect 12170 10308 12226 10364
rect 12226 10308 12230 10364
rect 12166 10304 12230 10308
rect 33874 10364 33938 10368
rect 33874 10308 33878 10364
rect 33878 10308 33934 10364
rect 33934 10308 33938 10364
rect 33874 10304 33938 10308
rect 33954 10364 34018 10368
rect 33954 10308 33958 10364
rect 33958 10308 34014 10364
rect 34014 10308 34018 10364
rect 33954 10304 34018 10308
rect 34034 10364 34098 10368
rect 34034 10308 34038 10364
rect 34038 10308 34094 10364
rect 34094 10308 34098 10364
rect 34034 10304 34098 10308
rect 34114 10364 34178 10368
rect 34114 10308 34118 10364
rect 34118 10308 34174 10364
rect 34174 10308 34178 10364
rect 34114 10304 34178 10308
rect 55822 10364 55886 10368
rect 55822 10308 55826 10364
rect 55826 10308 55882 10364
rect 55882 10308 55886 10364
rect 55822 10304 55886 10308
rect 55902 10364 55966 10368
rect 55902 10308 55906 10364
rect 55906 10308 55962 10364
rect 55962 10308 55966 10364
rect 55902 10304 55966 10308
rect 55982 10364 56046 10368
rect 55982 10308 55986 10364
rect 55986 10308 56042 10364
rect 56042 10308 56046 10364
rect 55982 10304 56046 10308
rect 56062 10364 56126 10368
rect 56062 10308 56066 10364
rect 56066 10308 56122 10364
rect 56122 10308 56126 10364
rect 56062 10304 56126 10308
rect 77770 10364 77834 10368
rect 77770 10308 77774 10364
rect 77774 10308 77830 10364
rect 77830 10308 77834 10364
rect 77770 10304 77834 10308
rect 77850 10364 77914 10368
rect 77850 10308 77854 10364
rect 77854 10308 77910 10364
rect 77910 10308 77914 10364
rect 77850 10304 77914 10308
rect 77930 10364 77994 10368
rect 77930 10308 77934 10364
rect 77934 10308 77990 10364
rect 77990 10308 77994 10364
rect 77930 10304 77994 10308
rect 78010 10364 78074 10368
rect 78010 10308 78014 10364
rect 78014 10308 78070 10364
rect 78070 10308 78074 10364
rect 78010 10304 78074 10308
rect 56916 10236 56980 10300
rect 22900 9820 22964 9824
rect 22900 9764 22904 9820
rect 22904 9764 22960 9820
rect 22960 9764 22964 9820
rect 22900 9760 22964 9764
rect 22980 9820 23044 9824
rect 22980 9764 22984 9820
rect 22984 9764 23040 9820
rect 23040 9764 23044 9820
rect 22980 9760 23044 9764
rect 23060 9820 23124 9824
rect 23060 9764 23064 9820
rect 23064 9764 23120 9820
rect 23120 9764 23124 9820
rect 23060 9760 23124 9764
rect 23140 9820 23204 9824
rect 23140 9764 23144 9820
rect 23144 9764 23200 9820
rect 23200 9764 23204 9820
rect 23140 9760 23204 9764
rect 44848 9820 44912 9824
rect 44848 9764 44852 9820
rect 44852 9764 44908 9820
rect 44908 9764 44912 9820
rect 44848 9760 44912 9764
rect 44928 9820 44992 9824
rect 44928 9764 44932 9820
rect 44932 9764 44988 9820
rect 44988 9764 44992 9820
rect 44928 9760 44992 9764
rect 45008 9820 45072 9824
rect 45008 9764 45012 9820
rect 45012 9764 45068 9820
rect 45068 9764 45072 9820
rect 45008 9760 45072 9764
rect 45088 9820 45152 9824
rect 45088 9764 45092 9820
rect 45092 9764 45148 9820
rect 45148 9764 45152 9820
rect 45088 9760 45152 9764
rect 66796 9820 66860 9824
rect 66796 9764 66800 9820
rect 66800 9764 66856 9820
rect 66856 9764 66860 9820
rect 66796 9760 66860 9764
rect 66876 9820 66940 9824
rect 66876 9764 66880 9820
rect 66880 9764 66936 9820
rect 66936 9764 66940 9820
rect 66876 9760 66940 9764
rect 66956 9820 67020 9824
rect 66956 9764 66960 9820
rect 66960 9764 67016 9820
rect 67016 9764 67020 9820
rect 66956 9760 67020 9764
rect 67036 9820 67100 9824
rect 67036 9764 67040 9820
rect 67040 9764 67096 9820
rect 67096 9764 67100 9820
rect 67036 9760 67100 9764
rect 11926 9276 11990 9280
rect 11926 9220 11930 9276
rect 11930 9220 11986 9276
rect 11986 9220 11990 9276
rect 11926 9216 11990 9220
rect 12006 9276 12070 9280
rect 12006 9220 12010 9276
rect 12010 9220 12066 9276
rect 12066 9220 12070 9276
rect 12006 9216 12070 9220
rect 12086 9276 12150 9280
rect 12086 9220 12090 9276
rect 12090 9220 12146 9276
rect 12146 9220 12150 9276
rect 12086 9216 12150 9220
rect 12166 9276 12230 9280
rect 12166 9220 12170 9276
rect 12170 9220 12226 9276
rect 12226 9220 12230 9276
rect 12166 9216 12230 9220
rect 33874 9276 33938 9280
rect 33874 9220 33878 9276
rect 33878 9220 33934 9276
rect 33934 9220 33938 9276
rect 33874 9216 33938 9220
rect 33954 9276 34018 9280
rect 33954 9220 33958 9276
rect 33958 9220 34014 9276
rect 34014 9220 34018 9276
rect 33954 9216 34018 9220
rect 34034 9276 34098 9280
rect 34034 9220 34038 9276
rect 34038 9220 34094 9276
rect 34094 9220 34098 9276
rect 34034 9216 34098 9220
rect 34114 9276 34178 9280
rect 34114 9220 34118 9276
rect 34118 9220 34174 9276
rect 34174 9220 34178 9276
rect 34114 9216 34178 9220
rect 55822 9276 55886 9280
rect 55822 9220 55826 9276
rect 55826 9220 55882 9276
rect 55882 9220 55886 9276
rect 55822 9216 55886 9220
rect 55902 9276 55966 9280
rect 55902 9220 55906 9276
rect 55906 9220 55962 9276
rect 55962 9220 55966 9276
rect 55902 9216 55966 9220
rect 55982 9276 56046 9280
rect 55982 9220 55986 9276
rect 55986 9220 56042 9276
rect 56042 9220 56046 9276
rect 55982 9216 56046 9220
rect 56062 9276 56126 9280
rect 56062 9220 56066 9276
rect 56066 9220 56122 9276
rect 56122 9220 56126 9276
rect 56062 9216 56126 9220
rect 77770 9276 77834 9280
rect 77770 9220 77774 9276
rect 77774 9220 77830 9276
rect 77830 9220 77834 9276
rect 77770 9216 77834 9220
rect 77850 9276 77914 9280
rect 77850 9220 77854 9276
rect 77854 9220 77910 9276
rect 77910 9220 77914 9276
rect 77850 9216 77914 9220
rect 77930 9276 77994 9280
rect 77930 9220 77934 9276
rect 77934 9220 77990 9276
rect 77990 9220 77994 9276
rect 77930 9216 77994 9220
rect 78010 9276 78074 9280
rect 78010 9220 78014 9276
rect 78014 9220 78070 9276
rect 78070 9220 78074 9276
rect 78010 9216 78074 9220
rect 22900 8732 22964 8736
rect 22900 8676 22904 8732
rect 22904 8676 22960 8732
rect 22960 8676 22964 8732
rect 22900 8672 22964 8676
rect 22980 8732 23044 8736
rect 22980 8676 22984 8732
rect 22984 8676 23040 8732
rect 23040 8676 23044 8732
rect 22980 8672 23044 8676
rect 23060 8732 23124 8736
rect 23060 8676 23064 8732
rect 23064 8676 23120 8732
rect 23120 8676 23124 8732
rect 23060 8672 23124 8676
rect 23140 8732 23204 8736
rect 23140 8676 23144 8732
rect 23144 8676 23200 8732
rect 23200 8676 23204 8732
rect 23140 8672 23204 8676
rect 44848 8732 44912 8736
rect 44848 8676 44852 8732
rect 44852 8676 44908 8732
rect 44908 8676 44912 8732
rect 44848 8672 44912 8676
rect 44928 8732 44992 8736
rect 44928 8676 44932 8732
rect 44932 8676 44988 8732
rect 44988 8676 44992 8732
rect 44928 8672 44992 8676
rect 45008 8732 45072 8736
rect 45008 8676 45012 8732
rect 45012 8676 45068 8732
rect 45068 8676 45072 8732
rect 45008 8672 45072 8676
rect 45088 8732 45152 8736
rect 45088 8676 45092 8732
rect 45092 8676 45148 8732
rect 45148 8676 45152 8732
rect 45088 8672 45152 8676
rect 66796 8732 66860 8736
rect 66796 8676 66800 8732
rect 66800 8676 66856 8732
rect 66856 8676 66860 8732
rect 66796 8672 66860 8676
rect 66876 8732 66940 8736
rect 66876 8676 66880 8732
rect 66880 8676 66936 8732
rect 66936 8676 66940 8732
rect 66876 8672 66940 8676
rect 66956 8732 67020 8736
rect 66956 8676 66960 8732
rect 66960 8676 67016 8732
rect 67016 8676 67020 8732
rect 66956 8672 67020 8676
rect 67036 8732 67100 8736
rect 67036 8676 67040 8732
rect 67040 8676 67096 8732
rect 67096 8676 67100 8732
rect 67036 8672 67100 8676
rect 11926 8188 11990 8192
rect 11926 8132 11930 8188
rect 11930 8132 11986 8188
rect 11986 8132 11990 8188
rect 11926 8128 11990 8132
rect 12006 8188 12070 8192
rect 12006 8132 12010 8188
rect 12010 8132 12066 8188
rect 12066 8132 12070 8188
rect 12006 8128 12070 8132
rect 12086 8188 12150 8192
rect 12086 8132 12090 8188
rect 12090 8132 12146 8188
rect 12146 8132 12150 8188
rect 12086 8128 12150 8132
rect 12166 8188 12230 8192
rect 12166 8132 12170 8188
rect 12170 8132 12226 8188
rect 12226 8132 12230 8188
rect 12166 8128 12230 8132
rect 33874 8188 33938 8192
rect 33874 8132 33878 8188
rect 33878 8132 33934 8188
rect 33934 8132 33938 8188
rect 33874 8128 33938 8132
rect 33954 8188 34018 8192
rect 33954 8132 33958 8188
rect 33958 8132 34014 8188
rect 34014 8132 34018 8188
rect 33954 8128 34018 8132
rect 34034 8188 34098 8192
rect 34034 8132 34038 8188
rect 34038 8132 34094 8188
rect 34094 8132 34098 8188
rect 34034 8128 34098 8132
rect 34114 8188 34178 8192
rect 34114 8132 34118 8188
rect 34118 8132 34174 8188
rect 34174 8132 34178 8188
rect 34114 8128 34178 8132
rect 55822 8188 55886 8192
rect 55822 8132 55826 8188
rect 55826 8132 55882 8188
rect 55882 8132 55886 8188
rect 55822 8128 55886 8132
rect 55902 8188 55966 8192
rect 55902 8132 55906 8188
rect 55906 8132 55962 8188
rect 55962 8132 55966 8188
rect 55902 8128 55966 8132
rect 55982 8188 56046 8192
rect 55982 8132 55986 8188
rect 55986 8132 56042 8188
rect 56042 8132 56046 8188
rect 55982 8128 56046 8132
rect 56062 8188 56126 8192
rect 56062 8132 56066 8188
rect 56066 8132 56122 8188
rect 56122 8132 56126 8188
rect 56062 8128 56126 8132
rect 77770 8188 77834 8192
rect 77770 8132 77774 8188
rect 77774 8132 77830 8188
rect 77830 8132 77834 8188
rect 77770 8128 77834 8132
rect 77850 8188 77914 8192
rect 77850 8132 77854 8188
rect 77854 8132 77910 8188
rect 77910 8132 77914 8188
rect 77850 8128 77914 8132
rect 77930 8188 77994 8192
rect 77930 8132 77934 8188
rect 77934 8132 77990 8188
rect 77990 8132 77994 8188
rect 77930 8128 77994 8132
rect 78010 8188 78074 8192
rect 78010 8132 78014 8188
rect 78014 8132 78070 8188
rect 78070 8132 78074 8188
rect 78010 8128 78074 8132
rect 22900 7644 22964 7648
rect 22900 7588 22904 7644
rect 22904 7588 22960 7644
rect 22960 7588 22964 7644
rect 22900 7584 22964 7588
rect 22980 7644 23044 7648
rect 22980 7588 22984 7644
rect 22984 7588 23040 7644
rect 23040 7588 23044 7644
rect 22980 7584 23044 7588
rect 23060 7644 23124 7648
rect 23060 7588 23064 7644
rect 23064 7588 23120 7644
rect 23120 7588 23124 7644
rect 23060 7584 23124 7588
rect 23140 7644 23204 7648
rect 23140 7588 23144 7644
rect 23144 7588 23200 7644
rect 23200 7588 23204 7644
rect 23140 7584 23204 7588
rect 44848 7644 44912 7648
rect 44848 7588 44852 7644
rect 44852 7588 44908 7644
rect 44908 7588 44912 7644
rect 44848 7584 44912 7588
rect 44928 7644 44992 7648
rect 44928 7588 44932 7644
rect 44932 7588 44988 7644
rect 44988 7588 44992 7644
rect 44928 7584 44992 7588
rect 45008 7644 45072 7648
rect 45008 7588 45012 7644
rect 45012 7588 45068 7644
rect 45068 7588 45072 7644
rect 45008 7584 45072 7588
rect 45088 7644 45152 7648
rect 45088 7588 45092 7644
rect 45092 7588 45148 7644
rect 45148 7588 45152 7644
rect 45088 7584 45152 7588
rect 66796 7644 66860 7648
rect 66796 7588 66800 7644
rect 66800 7588 66856 7644
rect 66856 7588 66860 7644
rect 66796 7584 66860 7588
rect 66876 7644 66940 7648
rect 66876 7588 66880 7644
rect 66880 7588 66936 7644
rect 66936 7588 66940 7644
rect 66876 7584 66940 7588
rect 66956 7644 67020 7648
rect 66956 7588 66960 7644
rect 66960 7588 67016 7644
rect 67016 7588 67020 7644
rect 66956 7584 67020 7588
rect 67036 7644 67100 7648
rect 67036 7588 67040 7644
rect 67040 7588 67096 7644
rect 67096 7588 67100 7644
rect 67036 7584 67100 7588
rect 11926 7100 11990 7104
rect 11926 7044 11930 7100
rect 11930 7044 11986 7100
rect 11986 7044 11990 7100
rect 11926 7040 11990 7044
rect 12006 7100 12070 7104
rect 12006 7044 12010 7100
rect 12010 7044 12066 7100
rect 12066 7044 12070 7100
rect 12006 7040 12070 7044
rect 12086 7100 12150 7104
rect 12086 7044 12090 7100
rect 12090 7044 12146 7100
rect 12146 7044 12150 7100
rect 12086 7040 12150 7044
rect 12166 7100 12230 7104
rect 12166 7044 12170 7100
rect 12170 7044 12226 7100
rect 12226 7044 12230 7100
rect 12166 7040 12230 7044
rect 33874 7100 33938 7104
rect 33874 7044 33878 7100
rect 33878 7044 33934 7100
rect 33934 7044 33938 7100
rect 33874 7040 33938 7044
rect 33954 7100 34018 7104
rect 33954 7044 33958 7100
rect 33958 7044 34014 7100
rect 34014 7044 34018 7100
rect 33954 7040 34018 7044
rect 34034 7100 34098 7104
rect 34034 7044 34038 7100
rect 34038 7044 34094 7100
rect 34094 7044 34098 7100
rect 34034 7040 34098 7044
rect 34114 7100 34178 7104
rect 34114 7044 34118 7100
rect 34118 7044 34174 7100
rect 34174 7044 34178 7100
rect 34114 7040 34178 7044
rect 55822 7100 55886 7104
rect 55822 7044 55826 7100
rect 55826 7044 55882 7100
rect 55882 7044 55886 7100
rect 55822 7040 55886 7044
rect 55902 7100 55966 7104
rect 55902 7044 55906 7100
rect 55906 7044 55962 7100
rect 55962 7044 55966 7100
rect 55902 7040 55966 7044
rect 55982 7100 56046 7104
rect 55982 7044 55986 7100
rect 55986 7044 56042 7100
rect 56042 7044 56046 7100
rect 55982 7040 56046 7044
rect 56062 7100 56126 7104
rect 56062 7044 56066 7100
rect 56066 7044 56122 7100
rect 56122 7044 56126 7100
rect 56062 7040 56126 7044
rect 77770 7100 77834 7104
rect 77770 7044 77774 7100
rect 77774 7044 77830 7100
rect 77830 7044 77834 7100
rect 77770 7040 77834 7044
rect 77850 7100 77914 7104
rect 77850 7044 77854 7100
rect 77854 7044 77910 7100
rect 77910 7044 77914 7100
rect 77850 7040 77914 7044
rect 77930 7100 77994 7104
rect 77930 7044 77934 7100
rect 77934 7044 77990 7100
rect 77990 7044 77994 7100
rect 77930 7040 77994 7044
rect 78010 7100 78074 7104
rect 78010 7044 78014 7100
rect 78014 7044 78070 7100
rect 78070 7044 78074 7100
rect 78010 7040 78074 7044
rect 22900 6556 22964 6560
rect 22900 6500 22904 6556
rect 22904 6500 22960 6556
rect 22960 6500 22964 6556
rect 22900 6496 22964 6500
rect 22980 6556 23044 6560
rect 22980 6500 22984 6556
rect 22984 6500 23040 6556
rect 23040 6500 23044 6556
rect 22980 6496 23044 6500
rect 23060 6556 23124 6560
rect 23060 6500 23064 6556
rect 23064 6500 23120 6556
rect 23120 6500 23124 6556
rect 23060 6496 23124 6500
rect 23140 6556 23204 6560
rect 23140 6500 23144 6556
rect 23144 6500 23200 6556
rect 23200 6500 23204 6556
rect 23140 6496 23204 6500
rect 44848 6556 44912 6560
rect 44848 6500 44852 6556
rect 44852 6500 44908 6556
rect 44908 6500 44912 6556
rect 44848 6496 44912 6500
rect 44928 6556 44992 6560
rect 44928 6500 44932 6556
rect 44932 6500 44988 6556
rect 44988 6500 44992 6556
rect 44928 6496 44992 6500
rect 45008 6556 45072 6560
rect 45008 6500 45012 6556
rect 45012 6500 45068 6556
rect 45068 6500 45072 6556
rect 45008 6496 45072 6500
rect 45088 6556 45152 6560
rect 45088 6500 45092 6556
rect 45092 6500 45148 6556
rect 45148 6500 45152 6556
rect 45088 6496 45152 6500
rect 66796 6556 66860 6560
rect 66796 6500 66800 6556
rect 66800 6500 66856 6556
rect 66856 6500 66860 6556
rect 66796 6496 66860 6500
rect 66876 6556 66940 6560
rect 66876 6500 66880 6556
rect 66880 6500 66936 6556
rect 66936 6500 66940 6556
rect 66876 6496 66940 6500
rect 66956 6556 67020 6560
rect 66956 6500 66960 6556
rect 66960 6500 67016 6556
rect 67016 6500 67020 6556
rect 66956 6496 67020 6500
rect 67036 6556 67100 6560
rect 67036 6500 67040 6556
rect 67040 6500 67096 6556
rect 67096 6500 67100 6556
rect 67036 6496 67100 6500
rect 11926 6012 11990 6016
rect 11926 5956 11930 6012
rect 11930 5956 11986 6012
rect 11986 5956 11990 6012
rect 11926 5952 11990 5956
rect 12006 6012 12070 6016
rect 12006 5956 12010 6012
rect 12010 5956 12066 6012
rect 12066 5956 12070 6012
rect 12006 5952 12070 5956
rect 12086 6012 12150 6016
rect 12086 5956 12090 6012
rect 12090 5956 12146 6012
rect 12146 5956 12150 6012
rect 12086 5952 12150 5956
rect 12166 6012 12230 6016
rect 12166 5956 12170 6012
rect 12170 5956 12226 6012
rect 12226 5956 12230 6012
rect 12166 5952 12230 5956
rect 33874 6012 33938 6016
rect 33874 5956 33878 6012
rect 33878 5956 33934 6012
rect 33934 5956 33938 6012
rect 33874 5952 33938 5956
rect 33954 6012 34018 6016
rect 33954 5956 33958 6012
rect 33958 5956 34014 6012
rect 34014 5956 34018 6012
rect 33954 5952 34018 5956
rect 34034 6012 34098 6016
rect 34034 5956 34038 6012
rect 34038 5956 34094 6012
rect 34094 5956 34098 6012
rect 34034 5952 34098 5956
rect 34114 6012 34178 6016
rect 34114 5956 34118 6012
rect 34118 5956 34174 6012
rect 34174 5956 34178 6012
rect 34114 5952 34178 5956
rect 55822 6012 55886 6016
rect 55822 5956 55826 6012
rect 55826 5956 55882 6012
rect 55882 5956 55886 6012
rect 55822 5952 55886 5956
rect 55902 6012 55966 6016
rect 55902 5956 55906 6012
rect 55906 5956 55962 6012
rect 55962 5956 55966 6012
rect 55902 5952 55966 5956
rect 55982 6012 56046 6016
rect 55982 5956 55986 6012
rect 55986 5956 56042 6012
rect 56042 5956 56046 6012
rect 55982 5952 56046 5956
rect 56062 6012 56126 6016
rect 56062 5956 56066 6012
rect 56066 5956 56122 6012
rect 56122 5956 56126 6012
rect 56062 5952 56126 5956
rect 77770 6012 77834 6016
rect 77770 5956 77774 6012
rect 77774 5956 77830 6012
rect 77830 5956 77834 6012
rect 77770 5952 77834 5956
rect 77850 6012 77914 6016
rect 77850 5956 77854 6012
rect 77854 5956 77910 6012
rect 77910 5956 77914 6012
rect 77850 5952 77914 5956
rect 77930 6012 77994 6016
rect 77930 5956 77934 6012
rect 77934 5956 77990 6012
rect 77990 5956 77994 6012
rect 77930 5952 77994 5956
rect 78010 6012 78074 6016
rect 78010 5956 78014 6012
rect 78014 5956 78070 6012
rect 78070 5956 78074 6012
rect 78010 5952 78074 5956
rect 22900 5468 22964 5472
rect 22900 5412 22904 5468
rect 22904 5412 22960 5468
rect 22960 5412 22964 5468
rect 22900 5408 22964 5412
rect 22980 5468 23044 5472
rect 22980 5412 22984 5468
rect 22984 5412 23040 5468
rect 23040 5412 23044 5468
rect 22980 5408 23044 5412
rect 23060 5468 23124 5472
rect 23060 5412 23064 5468
rect 23064 5412 23120 5468
rect 23120 5412 23124 5468
rect 23060 5408 23124 5412
rect 23140 5468 23204 5472
rect 23140 5412 23144 5468
rect 23144 5412 23200 5468
rect 23200 5412 23204 5468
rect 23140 5408 23204 5412
rect 44848 5468 44912 5472
rect 44848 5412 44852 5468
rect 44852 5412 44908 5468
rect 44908 5412 44912 5468
rect 44848 5408 44912 5412
rect 44928 5468 44992 5472
rect 44928 5412 44932 5468
rect 44932 5412 44988 5468
rect 44988 5412 44992 5468
rect 44928 5408 44992 5412
rect 45008 5468 45072 5472
rect 45008 5412 45012 5468
rect 45012 5412 45068 5468
rect 45068 5412 45072 5468
rect 45008 5408 45072 5412
rect 45088 5468 45152 5472
rect 45088 5412 45092 5468
rect 45092 5412 45148 5468
rect 45148 5412 45152 5468
rect 45088 5408 45152 5412
rect 66796 5468 66860 5472
rect 66796 5412 66800 5468
rect 66800 5412 66856 5468
rect 66856 5412 66860 5468
rect 66796 5408 66860 5412
rect 66876 5468 66940 5472
rect 66876 5412 66880 5468
rect 66880 5412 66936 5468
rect 66936 5412 66940 5468
rect 66876 5408 66940 5412
rect 66956 5468 67020 5472
rect 66956 5412 66960 5468
rect 66960 5412 67016 5468
rect 67016 5412 67020 5468
rect 66956 5408 67020 5412
rect 67036 5468 67100 5472
rect 67036 5412 67040 5468
rect 67040 5412 67096 5468
rect 67096 5412 67100 5468
rect 67036 5408 67100 5412
rect 11926 4924 11990 4928
rect 11926 4868 11930 4924
rect 11930 4868 11986 4924
rect 11986 4868 11990 4924
rect 11926 4864 11990 4868
rect 12006 4924 12070 4928
rect 12006 4868 12010 4924
rect 12010 4868 12066 4924
rect 12066 4868 12070 4924
rect 12006 4864 12070 4868
rect 12086 4924 12150 4928
rect 12086 4868 12090 4924
rect 12090 4868 12146 4924
rect 12146 4868 12150 4924
rect 12086 4864 12150 4868
rect 12166 4924 12230 4928
rect 12166 4868 12170 4924
rect 12170 4868 12226 4924
rect 12226 4868 12230 4924
rect 12166 4864 12230 4868
rect 33874 4924 33938 4928
rect 33874 4868 33878 4924
rect 33878 4868 33934 4924
rect 33934 4868 33938 4924
rect 33874 4864 33938 4868
rect 33954 4924 34018 4928
rect 33954 4868 33958 4924
rect 33958 4868 34014 4924
rect 34014 4868 34018 4924
rect 33954 4864 34018 4868
rect 34034 4924 34098 4928
rect 34034 4868 34038 4924
rect 34038 4868 34094 4924
rect 34094 4868 34098 4924
rect 34034 4864 34098 4868
rect 34114 4924 34178 4928
rect 34114 4868 34118 4924
rect 34118 4868 34174 4924
rect 34174 4868 34178 4924
rect 34114 4864 34178 4868
rect 55822 4924 55886 4928
rect 55822 4868 55826 4924
rect 55826 4868 55882 4924
rect 55882 4868 55886 4924
rect 55822 4864 55886 4868
rect 55902 4924 55966 4928
rect 55902 4868 55906 4924
rect 55906 4868 55962 4924
rect 55962 4868 55966 4924
rect 55902 4864 55966 4868
rect 55982 4924 56046 4928
rect 55982 4868 55986 4924
rect 55986 4868 56042 4924
rect 56042 4868 56046 4924
rect 55982 4864 56046 4868
rect 56062 4924 56126 4928
rect 56062 4868 56066 4924
rect 56066 4868 56122 4924
rect 56122 4868 56126 4924
rect 56062 4864 56126 4868
rect 77770 4924 77834 4928
rect 77770 4868 77774 4924
rect 77774 4868 77830 4924
rect 77830 4868 77834 4924
rect 77770 4864 77834 4868
rect 77850 4924 77914 4928
rect 77850 4868 77854 4924
rect 77854 4868 77910 4924
rect 77910 4868 77914 4924
rect 77850 4864 77914 4868
rect 77930 4924 77994 4928
rect 77930 4868 77934 4924
rect 77934 4868 77990 4924
rect 77990 4868 77994 4924
rect 77930 4864 77994 4868
rect 78010 4924 78074 4928
rect 78010 4868 78014 4924
rect 78014 4868 78070 4924
rect 78070 4868 78074 4924
rect 78010 4864 78074 4868
rect 22900 4380 22964 4384
rect 22900 4324 22904 4380
rect 22904 4324 22960 4380
rect 22960 4324 22964 4380
rect 22900 4320 22964 4324
rect 22980 4380 23044 4384
rect 22980 4324 22984 4380
rect 22984 4324 23040 4380
rect 23040 4324 23044 4380
rect 22980 4320 23044 4324
rect 23060 4380 23124 4384
rect 23060 4324 23064 4380
rect 23064 4324 23120 4380
rect 23120 4324 23124 4380
rect 23060 4320 23124 4324
rect 23140 4380 23204 4384
rect 23140 4324 23144 4380
rect 23144 4324 23200 4380
rect 23200 4324 23204 4380
rect 23140 4320 23204 4324
rect 44848 4380 44912 4384
rect 44848 4324 44852 4380
rect 44852 4324 44908 4380
rect 44908 4324 44912 4380
rect 44848 4320 44912 4324
rect 44928 4380 44992 4384
rect 44928 4324 44932 4380
rect 44932 4324 44988 4380
rect 44988 4324 44992 4380
rect 44928 4320 44992 4324
rect 45008 4380 45072 4384
rect 45008 4324 45012 4380
rect 45012 4324 45068 4380
rect 45068 4324 45072 4380
rect 45008 4320 45072 4324
rect 45088 4380 45152 4384
rect 45088 4324 45092 4380
rect 45092 4324 45148 4380
rect 45148 4324 45152 4380
rect 45088 4320 45152 4324
rect 66796 4380 66860 4384
rect 66796 4324 66800 4380
rect 66800 4324 66856 4380
rect 66856 4324 66860 4380
rect 66796 4320 66860 4324
rect 66876 4380 66940 4384
rect 66876 4324 66880 4380
rect 66880 4324 66936 4380
rect 66936 4324 66940 4380
rect 66876 4320 66940 4324
rect 66956 4380 67020 4384
rect 66956 4324 66960 4380
rect 66960 4324 67016 4380
rect 67016 4324 67020 4380
rect 66956 4320 67020 4324
rect 67036 4380 67100 4384
rect 67036 4324 67040 4380
rect 67040 4324 67096 4380
rect 67096 4324 67100 4380
rect 67036 4320 67100 4324
rect 11926 3836 11990 3840
rect 11926 3780 11930 3836
rect 11930 3780 11986 3836
rect 11986 3780 11990 3836
rect 11926 3776 11990 3780
rect 12006 3836 12070 3840
rect 12006 3780 12010 3836
rect 12010 3780 12066 3836
rect 12066 3780 12070 3836
rect 12006 3776 12070 3780
rect 12086 3836 12150 3840
rect 12086 3780 12090 3836
rect 12090 3780 12146 3836
rect 12146 3780 12150 3836
rect 12086 3776 12150 3780
rect 12166 3836 12230 3840
rect 12166 3780 12170 3836
rect 12170 3780 12226 3836
rect 12226 3780 12230 3836
rect 12166 3776 12230 3780
rect 33874 3836 33938 3840
rect 33874 3780 33878 3836
rect 33878 3780 33934 3836
rect 33934 3780 33938 3836
rect 33874 3776 33938 3780
rect 33954 3836 34018 3840
rect 33954 3780 33958 3836
rect 33958 3780 34014 3836
rect 34014 3780 34018 3836
rect 33954 3776 34018 3780
rect 34034 3836 34098 3840
rect 34034 3780 34038 3836
rect 34038 3780 34094 3836
rect 34094 3780 34098 3836
rect 34034 3776 34098 3780
rect 34114 3836 34178 3840
rect 34114 3780 34118 3836
rect 34118 3780 34174 3836
rect 34174 3780 34178 3836
rect 34114 3776 34178 3780
rect 55822 3836 55886 3840
rect 55822 3780 55826 3836
rect 55826 3780 55882 3836
rect 55882 3780 55886 3836
rect 55822 3776 55886 3780
rect 55902 3836 55966 3840
rect 55902 3780 55906 3836
rect 55906 3780 55962 3836
rect 55962 3780 55966 3836
rect 55902 3776 55966 3780
rect 55982 3836 56046 3840
rect 55982 3780 55986 3836
rect 55986 3780 56042 3836
rect 56042 3780 56046 3836
rect 55982 3776 56046 3780
rect 56062 3836 56126 3840
rect 56062 3780 56066 3836
rect 56066 3780 56122 3836
rect 56122 3780 56126 3836
rect 56062 3776 56126 3780
rect 77770 3836 77834 3840
rect 77770 3780 77774 3836
rect 77774 3780 77830 3836
rect 77830 3780 77834 3836
rect 77770 3776 77834 3780
rect 77850 3836 77914 3840
rect 77850 3780 77854 3836
rect 77854 3780 77910 3836
rect 77910 3780 77914 3836
rect 77850 3776 77914 3780
rect 77930 3836 77994 3840
rect 77930 3780 77934 3836
rect 77934 3780 77990 3836
rect 77990 3780 77994 3836
rect 77930 3776 77994 3780
rect 78010 3836 78074 3840
rect 78010 3780 78014 3836
rect 78014 3780 78070 3836
rect 78070 3780 78074 3836
rect 78010 3776 78074 3780
rect 22900 3292 22964 3296
rect 22900 3236 22904 3292
rect 22904 3236 22960 3292
rect 22960 3236 22964 3292
rect 22900 3232 22964 3236
rect 22980 3292 23044 3296
rect 22980 3236 22984 3292
rect 22984 3236 23040 3292
rect 23040 3236 23044 3292
rect 22980 3232 23044 3236
rect 23060 3292 23124 3296
rect 23060 3236 23064 3292
rect 23064 3236 23120 3292
rect 23120 3236 23124 3292
rect 23060 3232 23124 3236
rect 23140 3292 23204 3296
rect 23140 3236 23144 3292
rect 23144 3236 23200 3292
rect 23200 3236 23204 3292
rect 23140 3232 23204 3236
rect 44848 3292 44912 3296
rect 44848 3236 44852 3292
rect 44852 3236 44908 3292
rect 44908 3236 44912 3292
rect 44848 3232 44912 3236
rect 44928 3292 44992 3296
rect 44928 3236 44932 3292
rect 44932 3236 44988 3292
rect 44988 3236 44992 3292
rect 44928 3232 44992 3236
rect 45008 3292 45072 3296
rect 45008 3236 45012 3292
rect 45012 3236 45068 3292
rect 45068 3236 45072 3292
rect 45008 3232 45072 3236
rect 45088 3292 45152 3296
rect 45088 3236 45092 3292
rect 45092 3236 45148 3292
rect 45148 3236 45152 3292
rect 45088 3232 45152 3236
rect 66796 3292 66860 3296
rect 66796 3236 66800 3292
rect 66800 3236 66856 3292
rect 66856 3236 66860 3292
rect 66796 3232 66860 3236
rect 66876 3292 66940 3296
rect 66876 3236 66880 3292
rect 66880 3236 66936 3292
rect 66936 3236 66940 3292
rect 66876 3232 66940 3236
rect 66956 3292 67020 3296
rect 66956 3236 66960 3292
rect 66960 3236 67016 3292
rect 67016 3236 67020 3292
rect 66956 3232 67020 3236
rect 67036 3292 67100 3296
rect 67036 3236 67040 3292
rect 67040 3236 67096 3292
rect 67096 3236 67100 3292
rect 67036 3232 67100 3236
rect 11926 2748 11990 2752
rect 11926 2692 11930 2748
rect 11930 2692 11986 2748
rect 11986 2692 11990 2748
rect 11926 2688 11990 2692
rect 12006 2748 12070 2752
rect 12006 2692 12010 2748
rect 12010 2692 12066 2748
rect 12066 2692 12070 2748
rect 12006 2688 12070 2692
rect 12086 2748 12150 2752
rect 12086 2692 12090 2748
rect 12090 2692 12146 2748
rect 12146 2692 12150 2748
rect 12086 2688 12150 2692
rect 12166 2748 12230 2752
rect 12166 2692 12170 2748
rect 12170 2692 12226 2748
rect 12226 2692 12230 2748
rect 12166 2688 12230 2692
rect 33874 2748 33938 2752
rect 33874 2692 33878 2748
rect 33878 2692 33934 2748
rect 33934 2692 33938 2748
rect 33874 2688 33938 2692
rect 33954 2748 34018 2752
rect 33954 2692 33958 2748
rect 33958 2692 34014 2748
rect 34014 2692 34018 2748
rect 33954 2688 34018 2692
rect 34034 2748 34098 2752
rect 34034 2692 34038 2748
rect 34038 2692 34094 2748
rect 34094 2692 34098 2748
rect 34034 2688 34098 2692
rect 34114 2748 34178 2752
rect 34114 2692 34118 2748
rect 34118 2692 34174 2748
rect 34174 2692 34178 2748
rect 34114 2688 34178 2692
rect 55822 2748 55886 2752
rect 55822 2692 55826 2748
rect 55826 2692 55882 2748
rect 55882 2692 55886 2748
rect 55822 2688 55886 2692
rect 55902 2748 55966 2752
rect 55902 2692 55906 2748
rect 55906 2692 55962 2748
rect 55962 2692 55966 2748
rect 55902 2688 55966 2692
rect 55982 2748 56046 2752
rect 55982 2692 55986 2748
rect 55986 2692 56042 2748
rect 56042 2692 56046 2748
rect 55982 2688 56046 2692
rect 56062 2748 56126 2752
rect 56062 2692 56066 2748
rect 56066 2692 56122 2748
rect 56122 2692 56126 2748
rect 56062 2688 56126 2692
rect 77770 2748 77834 2752
rect 77770 2692 77774 2748
rect 77774 2692 77830 2748
rect 77830 2692 77834 2748
rect 77770 2688 77834 2692
rect 77850 2748 77914 2752
rect 77850 2692 77854 2748
rect 77854 2692 77910 2748
rect 77910 2692 77914 2748
rect 77850 2688 77914 2692
rect 77930 2748 77994 2752
rect 77930 2692 77934 2748
rect 77934 2692 77990 2748
rect 77990 2692 77994 2748
rect 77930 2688 77994 2692
rect 78010 2748 78074 2752
rect 78010 2692 78014 2748
rect 78014 2692 78070 2748
rect 78070 2692 78074 2748
rect 78010 2688 78074 2692
rect 22900 2204 22964 2208
rect 22900 2148 22904 2204
rect 22904 2148 22960 2204
rect 22960 2148 22964 2204
rect 22900 2144 22964 2148
rect 22980 2204 23044 2208
rect 22980 2148 22984 2204
rect 22984 2148 23040 2204
rect 23040 2148 23044 2204
rect 22980 2144 23044 2148
rect 23060 2204 23124 2208
rect 23060 2148 23064 2204
rect 23064 2148 23120 2204
rect 23120 2148 23124 2204
rect 23060 2144 23124 2148
rect 23140 2204 23204 2208
rect 23140 2148 23144 2204
rect 23144 2148 23200 2204
rect 23200 2148 23204 2204
rect 23140 2144 23204 2148
rect 44848 2204 44912 2208
rect 44848 2148 44852 2204
rect 44852 2148 44908 2204
rect 44908 2148 44912 2204
rect 44848 2144 44912 2148
rect 44928 2204 44992 2208
rect 44928 2148 44932 2204
rect 44932 2148 44988 2204
rect 44988 2148 44992 2204
rect 44928 2144 44992 2148
rect 45008 2204 45072 2208
rect 45008 2148 45012 2204
rect 45012 2148 45068 2204
rect 45068 2148 45072 2204
rect 45008 2144 45072 2148
rect 45088 2204 45152 2208
rect 45088 2148 45092 2204
rect 45092 2148 45148 2204
rect 45148 2148 45152 2204
rect 45088 2144 45152 2148
rect 66796 2204 66860 2208
rect 66796 2148 66800 2204
rect 66800 2148 66856 2204
rect 66856 2148 66860 2204
rect 66796 2144 66860 2148
rect 66876 2204 66940 2208
rect 66876 2148 66880 2204
rect 66880 2148 66936 2204
rect 66936 2148 66940 2204
rect 66876 2144 66940 2148
rect 66956 2204 67020 2208
rect 66956 2148 66960 2204
rect 66960 2148 67016 2204
rect 67016 2148 67020 2204
rect 66956 2144 67020 2148
rect 67036 2204 67100 2208
rect 67036 2148 67040 2204
rect 67040 2148 67096 2204
rect 67096 2148 67100 2204
rect 67036 2144 67100 2148
<< metal4 >>
rect 11918 27776 12238 27792
rect 11918 27712 11926 27776
rect 11990 27712 12006 27776
rect 12070 27712 12086 27776
rect 12150 27712 12166 27776
rect 12230 27712 12238 27776
rect 11918 26688 12238 27712
rect 11918 26624 11926 26688
rect 11990 26624 12006 26688
rect 12070 26624 12086 26688
rect 12150 26624 12166 26688
rect 12230 26624 12238 26688
rect 11918 25600 12238 26624
rect 11918 25536 11926 25600
rect 11990 25536 12006 25600
rect 12070 25536 12086 25600
rect 12150 25536 12166 25600
rect 12230 25536 12238 25600
rect 11918 24512 12238 25536
rect 11918 24448 11926 24512
rect 11990 24448 12006 24512
rect 12070 24448 12086 24512
rect 12150 24448 12166 24512
rect 12230 24448 12238 24512
rect 11918 23424 12238 24448
rect 11918 23360 11926 23424
rect 11990 23360 12006 23424
rect 12070 23360 12086 23424
rect 12150 23360 12166 23424
rect 12230 23360 12238 23424
rect 11918 22336 12238 23360
rect 11918 22272 11926 22336
rect 11990 22272 12006 22336
rect 12070 22272 12086 22336
rect 12150 22272 12166 22336
rect 12230 22272 12238 22336
rect 11918 21248 12238 22272
rect 11918 21184 11926 21248
rect 11990 21184 12006 21248
rect 12070 21184 12086 21248
rect 12150 21184 12166 21248
rect 12230 21184 12238 21248
rect 11918 20160 12238 21184
rect 11918 20096 11926 20160
rect 11990 20096 12006 20160
rect 12070 20096 12086 20160
rect 12150 20096 12166 20160
rect 12230 20096 12238 20160
rect 11918 19072 12238 20096
rect 11918 19008 11926 19072
rect 11990 19008 12006 19072
rect 12070 19008 12086 19072
rect 12150 19008 12166 19072
rect 12230 19008 12238 19072
rect 11918 17984 12238 19008
rect 11918 17920 11926 17984
rect 11990 17920 12006 17984
rect 12070 17920 12086 17984
rect 12150 17920 12166 17984
rect 12230 17920 12238 17984
rect 11918 16896 12238 17920
rect 11918 16832 11926 16896
rect 11990 16832 12006 16896
rect 12070 16832 12086 16896
rect 12150 16832 12166 16896
rect 12230 16832 12238 16896
rect 11918 15808 12238 16832
rect 11918 15744 11926 15808
rect 11990 15744 12006 15808
rect 12070 15744 12086 15808
rect 12150 15744 12166 15808
rect 12230 15744 12238 15808
rect 11918 14720 12238 15744
rect 11918 14656 11926 14720
rect 11990 14656 12006 14720
rect 12070 14656 12086 14720
rect 12150 14656 12166 14720
rect 12230 14656 12238 14720
rect 11918 13632 12238 14656
rect 11918 13568 11926 13632
rect 11990 13568 12006 13632
rect 12070 13568 12086 13632
rect 12150 13568 12166 13632
rect 12230 13568 12238 13632
rect 11918 12544 12238 13568
rect 11918 12480 11926 12544
rect 11990 12480 12006 12544
rect 12070 12480 12086 12544
rect 12150 12480 12166 12544
rect 12230 12480 12238 12544
rect 11918 11456 12238 12480
rect 11918 11392 11926 11456
rect 11990 11392 12006 11456
rect 12070 11392 12086 11456
rect 12150 11392 12166 11456
rect 12230 11392 12238 11456
rect 11918 10368 12238 11392
rect 11918 10304 11926 10368
rect 11990 10304 12006 10368
rect 12070 10304 12086 10368
rect 12150 10304 12166 10368
rect 12230 10304 12238 10368
rect 11918 9280 12238 10304
rect 11918 9216 11926 9280
rect 11990 9216 12006 9280
rect 12070 9216 12086 9280
rect 12150 9216 12166 9280
rect 12230 9216 12238 9280
rect 11918 8192 12238 9216
rect 11918 8128 11926 8192
rect 11990 8128 12006 8192
rect 12070 8128 12086 8192
rect 12150 8128 12166 8192
rect 12230 8128 12238 8192
rect 11918 7104 12238 8128
rect 11918 7040 11926 7104
rect 11990 7040 12006 7104
rect 12070 7040 12086 7104
rect 12150 7040 12166 7104
rect 12230 7040 12238 7104
rect 11918 6016 12238 7040
rect 11918 5952 11926 6016
rect 11990 5952 12006 6016
rect 12070 5952 12086 6016
rect 12150 5952 12166 6016
rect 12230 5952 12238 6016
rect 11918 4928 12238 5952
rect 11918 4864 11926 4928
rect 11990 4864 12006 4928
rect 12070 4864 12086 4928
rect 12150 4864 12166 4928
rect 12230 4864 12238 4928
rect 11918 3840 12238 4864
rect 11918 3776 11926 3840
rect 11990 3776 12006 3840
rect 12070 3776 12086 3840
rect 12150 3776 12166 3840
rect 12230 3776 12238 3840
rect 11918 2752 12238 3776
rect 11918 2688 11926 2752
rect 11990 2688 12006 2752
rect 12070 2688 12086 2752
rect 12150 2688 12166 2752
rect 12230 2688 12238 2752
rect 11918 2128 12238 2688
rect 22892 27232 23212 27792
rect 22892 27168 22900 27232
rect 22964 27168 22980 27232
rect 23044 27168 23060 27232
rect 23124 27168 23140 27232
rect 23204 27168 23212 27232
rect 22892 26144 23212 27168
rect 22892 26080 22900 26144
rect 22964 26080 22980 26144
rect 23044 26080 23060 26144
rect 23124 26080 23140 26144
rect 23204 26080 23212 26144
rect 22892 25056 23212 26080
rect 33866 27776 34186 27792
rect 33866 27712 33874 27776
rect 33938 27712 33954 27776
rect 34018 27712 34034 27776
rect 34098 27712 34114 27776
rect 34178 27712 34186 27776
rect 33866 26688 34186 27712
rect 33866 26624 33874 26688
rect 33938 26624 33954 26688
rect 34018 26624 34034 26688
rect 34098 26624 34114 26688
rect 34178 26624 34186 26688
rect 28027 25804 28093 25805
rect 28027 25740 28028 25804
rect 28092 25740 28093 25804
rect 28027 25739 28093 25740
rect 22892 24992 22900 25056
rect 22964 24992 22980 25056
rect 23044 24992 23060 25056
rect 23124 24992 23140 25056
rect 23204 24992 23212 25056
rect 22892 23968 23212 24992
rect 27475 24172 27541 24173
rect 27475 24108 27476 24172
rect 27540 24108 27541 24172
rect 27475 24107 27541 24108
rect 22892 23904 22900 23968
rect 22964 23904 22980 23968
rect 23044 23904 23060 23968
rect 23124 23904 23140 23968
rect 23204 23904 23212 23968
rect 22892 22880 23212 23904
rect 22892 22816 22900 22880
rect 22964 22816 22980 22880
rect 23044 22816 23060 22880
rect 23124 22816 23140 22880
rect 23204 22816 23212 22880
rect 22892 21792 23212 22816
rect 22892 21728 22900 21792
rect 22964 21728 22980 21792
rect 23044 21728 23060 21792
rect 23124 21728 23140 21792
rect 23204 21728 23212 21792
rect 22892 20704 23212 21728
rect 26555 21452 26621 21453
rect 26555 21388 26556 21452
rect 26620 21388 26621 21452
rect 26555 21387 26621 21388
rect 22892 20640 22900 20704
rect 22964 20640 22980 20704
rect 23044 20640 23060 20704
rect 23124 20640 23140 20704
rect 23204 20640 23212 20704
rect 22892 19616 23212 20640
rect 22892 19552 22900 19616
rect 22964 19552 22980 19616
rect 23044 19552 23060 19616
rect 23124 19552 23140 19616
rect 23204 19552 23212 19616
rect 22892 18528 23212 19552
rect 22892 18464 22900 18528
rect 22964 18464 22980 18528
rect 23044 18464 23060 18528
rect 23124 18464 23140 18528
rect 23204 18464 23212 18528
rect 22892 17440 23212 18464
rect 22892 17376 22900 17440
rect 22964 17376 22980 17440
rect 23044 17376 23060 17440
rect 23124 17376 23140 17440
rect 23204 17376 23212 17440
rect 22892 16352 23212 17376
rect 22892 16288 22900 16352
rect 22964 16288 22980 16352
rect 23044 16288 23060 16352
rect 23124 16288 23140 16352
rect 23204 16288 23212 16352
rect 22892 15264 23212 16288
rect 22892 15200 22900 15264
rect 22964 15200 22980 15264
rect 23044 15200 23060 15264
rect 23124 15200 23140 15264
rect 23204 15200 23212 15264
rect 22892 14176 23212 15200
rect 22892 14112 22900 14176
rect 22964 14112 22980 14176
rect 23044 14112 23060 14176
rect 23124 14112 23140 14176
rect 23204 14112 23212 14176
rect 22892 13088 23212 14112
rect 22892 13024 22900 13088
rect 22964 13024 22980 13088
rect 23044 13024 23060 13088
rect 23124 13024 23140 13088
rect 23204 13024 23212 13088
rect 22892 12000 23212 13024
rect 26558 12885 26618 21387
rect 27478 15197 27538 24107
rect 28030 15605 28090 25739
rect 33866 25600 34186 26624
rect 33866 25536 33874 25600
rect 33938 25536 33954 25600
rect 34018 25536 34034 25600
rect 34098 25536 34114 25600
rect 34178 25536 34186 25600
rect 33866 24512 34186 25536
rect 33866 24448 33874 24512
rect 33938 24448 33954 24512
rect 34018 24448 34034 24512
rect 34098 24448 34114 24512
rect 34178 24448 34186 24512
rect 33866 23424 34186 24448
rect 33866 23360 33874 23424
rect 33938 23360 33954 23424
rect 34018 23360 34034 23424
rect 34098 23360 34114 23424
rect 34178 23360 34186 23424
rect 33866 22336 34186 23360
rect 33866 22272 33874 22336
rect 33938 22272 33954 22336
rect 34018 22272 34034 22336
rect 34098 22272 34114 22336
rect 34178 22272 34186 22336
rect 33866 21248 34186 22272
rect 33866 21184 33874 21248
rect 33938 21184 33954 21248
rect 34018 21184 34034 21248
rect 34098 21184 34114 21248
rect 34178 21184 34186 21248
rect 33866 20160 34186 21184
rect 33866 20096 33874 20160
rect 33938 20096 33954 20160
rect 34018 20096 34034 20160
rect 34098 20096 34114 20160
rect 34178 20096 34186 20160
rect 33866 19072 34186 20096
rect 33866 19008 33874 19072
rect 33938 19008 33954 19072
rect 34018 19008 34034 19072
rect 34098 19008 34114 19072
rect 34178 19008 34186 19072
rect 33866 17984 34186 19008
rect 33866 17920 33874 17984
rect 33938 17920 33954 17984
rect 34018 17920 34034 17984
rect 34098 17920 34114 17984
rect 34178 17920 34186 17984
rect 33866 16896 34186 17920
rect 33866 16832 33874 16896
rect 33938 16832 33954 16896
rect 34018 16832 34034 16896
rect 34098 16832 34114 16896
rect 34178 16832 34186 16896
rect 33866 15808 34186 16832
rect 33866 15744 33874 15808
rect 33938 15744 33954 15808
rect 34018 15744 34034 15808
rect 34098 15744 34114 15808
rect 34178 15744 34186 15808
rect 28027 15604 28093 15605
rect 28027 15540 28028 15604
rect 28092 15540 28093 15604
rect 28027 15539 28093 15540
rect 27475 15196 27541 15197
rect 27475 15132 27476 15196
rect 27540 15132 27541 15196
rect 27475 15131 27541 15132
rect 33866 14720 34186 15744
rect 33866 14656 33874 14720
rect 33938 14656 33954 14720
rect 34018 14656 34034 14720
rect 34098 14656 34114 14720
rect 34178 14656 34186 14720
rect 33866 13632 34186 14656
rect 33866 13568 33874 13632
rect 33938 13568 33954 13632
rect 34018 13568 34034 13632
rect 34098 13568 34114 13632
rect 34178 13568 34186 13632
rect 26555 12884 26621 12885
rect 26555 12820 26556 12884
rect 26620 12820 26621 12884
rect 26555 12819 26621 12820
rect 22892 11936 22900 12000
rect 22964 11936 22980 12000
rect 23044 11936 23060 12000
rect 23124 11936 23140 12000
rect 23204 11936 23212 12000
rect 22892 10912 23212 11936
rect 22892 10848 22900 10912
rect 22964 10848 22980 10912
rect 23044 10848 23060 10912
rect 23124 10848 23140 10912
rect 23204 10848 23212 10912
rect 22892 9824 23212 10848
rect 22892 9760 22900 9824
rect 22964 9760 22980 9824
rect 23044 9760 23060 9824
rect 23124 9760 23140 9824
rect 23204 9760 23212 9824
rect 22892 8736 23212 9760
rect 22892 8672 22900 8736
rect 22964 8672 22980 8736
rect 23044 8672 23060 8736
rect 23124 8672 23140 8736
rect 23204 8672 23212 8736
rect 22892 7648 23212 8672
rect 22892 7584 22900 7648
rect 22964 7584 22980 7648
rect 23044 7584 23060 7648
rect 23124 7584 23140 7648
rect 23204 7584 23212 7648
rect 22892 6560 23212 7584
rect 22892 6496 22900 6560
rect 22964 6496 22980 6560
rect 23044 6496 23060 6560
rect 23124 6496 23140 6560
rect 23204 6496 23212 6560
rect 22892 5472 23212 6496
rect 22892 5408 22900 5472
rect 22964 5408 22980 5472
rect 23044 5408 23060 5472
rect 23124 5408 23140 5472
rect 23204 5408 23212 5472
rect 22892 4384 23212 5408
rect 22892 4320 22900 4384
rect 22964 4320 22980 4384
rect 23044 4320 23060 4384
rect 23124 4320 23140 4384
rect 23204 4320 23212 4384
rect 22892 3296 23212 4320
rect 22892 3232 22900 3296
rect 22964 3232 22980 3296
rect 23044 3232 23060 3296
rect 23124 3232 23140 3296
rect 23204 3232 23212 3296
rect 22892 2208 23212 3232
rect 22892 2144 22900 2208
rect 22964 2144 22980 2208
rect 23044 2144 23060 2208
rect 23124 2144 23140 2208
rect 23204 2144 23212 2208
rect 22892 2128 23212 2144
rect 33866 12544 34186 13568
rect 33866 12480 33874 12544
rect 33938 12480 33954 12544
rect 34018 12480 34034 12544
rect 34098 12480 34114 12544
rect 34178 12480 34186 12544
rect 33866 11456 34186 12480
rect 33866 11392 33874 11456
rect 33938 11392 33954 11456
rect 34018 11392 34034 11456
rect 34098 11392 34114 11456
rect 34178 11392 34186 11456
rect 33866 10368 34186 11392
rect 33866 10304 33874 10368
rect 33938 10304 33954 10368
rect 34018 10304 34034 10368
rect 34098 10304 34114 10368
rect 34178 10304 34186 10368
rect 33866 9280 34186 10304
rect 33866 9216 33874 9280
rect 33938 9216 33954 9280
rect 34018 9216 34034 9280
rect 34098 9216 34114 9280
rect 34178 9216 34186 9280
rect 33866 8192 34186 9216
rect 33866 8128 33874 8192
rect 33938 8128 33954 8192
rect 34018 8128 34034 8192
rect 34098 8128 34114 8192
rect 34178 8128 34186 8192
rect 33866 7104 34186 8128
rect 33866 7040 33874 7104
rect 33938 7040 33954 7104
rect 34018 7040 34034 7104
rect 34098 7040 34114 7104
rect 34178 7040 34186 7104
rect 33866 6016 34186 7040
rect 33866 5952 33874 6016
rect 33938 5952 33954 6016
rect 34018 5952 34034 6016
rect 34098 5952 34114 6016
rect 34178 5952 34186 6016
rect 33866 4928 34186 5952
rect 33866 4864 33874 4928
rect 33938 4864 33954 4928
rect 34018 4864 34034 4928
rect 34098 4864 34114 4928
rect 34178 4864 34186 4928
rect 33866 3840 34186 4864
rect 33866 3776 33874 3840
rect 33938 3776 33954 3840
rect 34018 3776 34034 3840
rect 34098 3776 34114 3840
rect 34178 3776 34186 3840
rect 33866 2752 34186 3776
rect 33866 2688 33874 2752
rect 33938 2688 33954 2752
rect 34018 2688 34034 2752
rect 34098 2688 34114 2752
rect 34178 2688 34186 2752
rect 33866 2128 34186 2688
rect 44840 27232 45160 27792
rect 44840 27168 44848 27232
rect 44912 27168 44928 27232
rect 44992 27168 45008 27232
rect 45072 27168 45088 27232
rect 45152 27168 45160 27232
rect 44840 26144 45160 27168
rect 44840 26080 44848 26144
rect 44912 26080 44928 26144
rect 44992 26080 45008 26144
rect 45072 26080 45088 26144
rect 45152 26080 45160 26144
rect 44840 25056 45160 26080
rect 44840 24992 44848 25056
rect 44912 24992 44928 25056
rect 44992 24992 45008 25056
rect 45072 24992 45088 25056
rect 45152 24992 45160 25056
rect 44840 23968 45160 24992
rect 44840 23904 44848 23968
rect 44912 23904 44928 23968
rect 44992 23904 45008 23968
rect 45072 23904 45088 23968
rect 45152 23904 45160 23968
rect 44840 22880 45160 23904
rect 44840 22816 44848 22880
rect 44912 22816 44928 22880
rect 44992 22816 45008 22880
rect 45072 22816 45088 22880
rect 45152 22816 45160 22880
rect 44840 21792 45160 22816
rect 44840 21728 44848 21792
rect 44912 21728 44928 21792
rect 44992 21728 45008 21792
rect 45072 21728 45088 21792
rect 45152 21728 45160 21792
rect 44840 20704 45160 21728
rect 44840 20640 44848 20704
rect 44912 20640 44928 20704
rect 44992 20640 45008 20704
rect 45072 20640 45088 20704
rect 45152 20640 45160 20704
rect 44840 19616 45160 20640
rect 44840 19552 44848 19616
rect 44912 19552 44928 19616
rect 44992 19552 45008 19616
rect 45072 19552 45088 19616
rect 45152 19552 45160 19616
rect 44840 18528 45160 19552
rect 44840 18464 44848 18528
rect 44912 18464 44928 18528
rect 44992 18464 45008 18528
rect 45072 18464 45088 18528
rect 45152 18464 45160 18528
rect 44840 17440 45160 18464
rect 44840 17376 44848 17440
rect 44912 17376 44928 17440
rect 44992 17376 45008 17440
rect 45072 17376 45088 17440
rect 45152 17376 45160 17440
rect 44840 16352 45160 17376
rect 44840 16288 44848 16352
rect 44912 16288 44928 16352
rect 44992 16288 45008 16352
rect 45072 16288 45088 16352
rect 45152 16288 45160 16352
rect 44840 15264 45160 16288
rect 55814 27776 56134 27792
rect 55814 27712 55822 27776
rect 55886 27712 55902 27776
rect 55966 27712 55982 27776
rect 56046 27712 56062 27776
rect 56126 27712 56134 27776
rect 55814 26688 56134 27712
rect 55814 26624 55822 26688
rect 55886 26624 55902 26688
rect 55966 26624 55982 26688
rect 56046 26624 56062 26688
rect 56126 26624 56134 26688
rect 55814 25600 56134 26624
rect 55814 25536 55822 25600
rect 55886 25536 55902 25600
rect 55966 25536 55982 25600
rect 56046 25536 56062 25600
rect 56126 25536 56134 25600
rect 55814 24512 56134 25536
rect 55814 24448 55822 24512
rect 55886 24448 55902 24512
rect 55966 24448 55982 24512
rect 56046 24448 56062 24512
rect 56126 24448 56134 24512
rect 55814 23424 56134 24448
rect 55814 23360 55822 23424
rect 55886 23360 55902 23424
rect 55966 23360 55982 23424
rect 56046 23360 56062 23424
rect 56126 23360 56134 23424
rect 55814 22336 56134 23360
rect 55814 22272 55822 22336
rect 55886 22272 55902 22336
rect 55966 22272 55982 22336
rect 56046 22272 56062 22336
rect 56126 22272 56134 22336
rect 55814 21248 56134 22272
rect 55814 21184 55822 21248
rect 55886 21184 55902 21248
rect 55966 21184 55982 21248
rect 56046 21184 56062 21248
rect 56126 21184 56134 21248
rect 55814 20160 56134 21184
rect 55814 20096 55822 20160
rect 55886 20096 55902 20160
rect 55966 20096 55982 20160
rect 56046 20096 56062 20160
rect 56126 20096 56134 20160
rect 55814 19072 56134 20096
rect 55814 19008 55822 19072
rect 55886 19008 55902 19072
rect 55966 19008 55982 19072
rect 56046 19008 56062 19072
rect 56126 19008 56134 19072
rect 55814 17984 56134 19008
rect 66788 27232 67108 27792
rect 66788 27168 66796 27232
rect 66860 27168 66876 27232
rect 66940 27168 66956 27232
rect 67020 27168 67036 27232
rect 67100 27168 67108 27232
rect 66788 26144 67108 27168
rect 66788 26080 66796 26144
rect 66860 26080 66876 26144
rect 66940 26080 66956 26144
rect 67020 26080 67036 26144
rect 67100 26080 67108 26144
rect 66788 25056 67108 26080
rect 66788 24992 66796 25056
rect 66860 24992 66876 25056
rect 66940 24992 66956 25056
rect 67020 24992 67036 25056
rect 67100 24992 67108 25056
rect 66788 23968 67108 24992
rect 66788 23904 66796 23968
rect 66860 23904 66876 23968
rect 66940 23904 66956 23968
rect 67020 23904 67036 23968
rect 67100 23904 67108 23968
rect 66788 22880 67108 23904
rect 66788 22816 66796 22880
rect 66860 22816 66876 22880
rect 66940 22816 66956 22880
rect 67020 22816 67036 22880
rect 67100 22816 67108 22880
rect 66788 21792 67108 22816
rect 66788 21728 66796 21792
rect 66860 21728 66876 21792
rect 66940 21728 66956 21792
rect 67020 21728 67036 21792
rect 67100 21728 67108 21792
rect 66788 20704 67108 21728
rect 66788 20640 66796 20704
rect 66860 20640 66876 20704
rect 66940 20640 66956 20704
rect 67020 20640 67036 20704
rect 67100 20640 67108 20704
rect 66788 19616 67108 20640
rect 66788 19552 66796 19616
rect 66860 19552 66876 19616
rect 66940 19552 66956 19616
rect 67020 19552 67036 19616
rect 67100 19552 67108 19616
rect 66788 18528 67108 19552
rect 66788 18464 66796 18528
rect 66860 18464 66876 18528
rect 66940 18464 66956 18528
rect 67020 18464 67036 18528
rect 67100 18464 67108 18528
rect 56363 18324 56429 18325
rect 56363 18260 56364 18324
rect 56428 18260 56429 18324
rect 56363 18259 56429 18260
rect 55814 17920 55822 17984
rect 55886 17920 55902 17984
rect 55966 17920 55982 17984
rect 56046 17920 56062 17984
rect 56126 17920 56134 17984
rect 55814 16896 56134 17920
rect 55814 16832 55822 16896
rect 55886 16832 55902 16896
rect 55966 16832 55982 16896
rect 56046 16832 56062 16896
rect 56126 16832 56134 16896
rect 55627 16148 55693 16149
rect 55627 16084 55628 16148
rect 55692 16084 55693 16148
rect 55627 16083 55693 16084
rect 44840 15200 44848 15264
rect 44912 15200 44928 15264
rect 44992 15200 45008 15264
rect 45072 15200 45088 15264
rect 45152 15200 45160 15264
rect 44840 14176 45160 15200
rect 44840 14112 44848 14176
rect 44912 14112 44928 14176
rect 44992 14112 45008 14176
rect 45072 14112 45088 14176
rect 45152 14112 45160 14176
rect 44840 13088 45160 14112
rect 55630 13565 55690 16083
rect 55814 15808 56134 16832
rect 55814 15744 55822 15808
rect 55886 15744 55902 15808
rect 55966 15744 55982 15808
rect 56046 15744 56062 15808
rect 56126 15744 56134 15808
rect 55814 14720 56134 15744
rect 55814 14656 55822 14720
rect 55886 14656 55902 14720
rect 55966 14656 55982 14720
rect 56046 14656 56062 14720
rect 56126 14656 56134 14720
rect 55814 13632 56134 14656
rect 55814 13568 55822 13632
rect 55886 13568 55902 13632
rect 55966 13568 55982 13632
rect 56046 13568 56062 13632
rect 56126 13568 56134 13632
rect 55627 13564 55693 13565
rect 55627 13500 55628 13564
rect 55692 13500 55693 13564
rect 55627 13499 55693 13500
rect 44840 13024 44848 13088
rect 44912 13024 44928 13088
rect 44992 13024 45008 13088
rect 45072 13024 45088 13088
rect 45152 13024 45160 13088
rect 44840 12000 45160 13024
rect 44840 11936 44848 12000
rect 44912 11936 44928 12000
rect 44992 11936 45008 12000
rect 45072 11936 45088 12000
rect 45152 11936 45160 12000
rect 44840 10912 45160 11936
rect 44840 10848 44848 10912
rect 44912 10848 44928 10912
rect 44992 10848 45008 10912
rect 45072 10848 45088 10912
rect 45152 10848 45160 10912
rect 44840 9824 45160 10848
rect 44840 9760 44848 9824
rect 44912 9760 44928 9824
rect 44992 9760 45008 9824
rect 45072 9760 45088 9824
rect 45152 9760 45160 9824
rect 44840 8736 45160 9760
rect 44840 8672 44848 8736
rect 44912 8672 44928 8736
rect 44992 8672 45008 8736
rect 45072 8672 45088 8736
rect 45152 8672 45160 8736
rect 44840 7648 45160 8672
rect 44840 7584 44848 7648
rect 44912 7584 44928 7648
rect 44992 7584 45008 7648
rect 45072 7584 45088 7648
rect 45152 7584 45160 7648
rect 44840 6560 45160 7584
rect 44840 6496 44848 6560
rect 44912 6496 44928 6560
rect 44992 6496 45008 6560
rect 45072 6496 45088 6560
rect 45152 6496 45160 6560
rect 44840 5472 45160 6496
rect 44840 5408 44848 5472
rect 44912 5408 44928 5472
rect 44992 5408 45008 5472
rect 45072 5408 45088 5472
rect 45152 5408 45160 5472
rect 44840 4384 45160 5408
rect 44840 4320 44848 4384
rect 44912 4320 44928 4384
rect 44992 4320 45008 4384
rect 45072 4320 45088 4384
rect 45152 4320 45160 4384
rect 44840 3296 45160 4320
rect 44840 3232 44848 3296
rect 44912 3232 44928 3296
rect 44992 3232 45008 3296
rect 45072 3232 45088 3296
rect 45152 3232 45160 3296
rect 44840 2208 45160 3232
rect 44840 2144 44848 2208
rect 44912 2144 44928 2208
rect 44992 2144 45008 2208
rect 45072 2144 45088 2208
rect 45152 2144 45160 2208
rect 44840 2128 45160 2144
rect 55814 12544 56134 13568
rect 55814 12480 55822 12544
rect 55886 12480 55902 12544
rect 55966 12480 55982 12544
rect 56046 12480 56062 12544
rect 56126 12480 56134 12544
rect 55814 11456 56134 12480
rect 56366 11525 56426 18259
rect 66788 17440 67108 18464
rect 66788 17376 66796 17440
rect 66860 17376 66876 17440
rect 66940 17376 66956 17440
rect 67020 17376 67036 17440
rect 67100 17376 67108 17440
rect 66788 16352 67108 17376
rect 66788 16288 66796 16352
rect 66860 16288 66876 16352
rect 66940 16288 66956 16352
rect 67020 16288 67036 16352
rect 67100 16288 67108 16352
rect 66788 15264 67108 16288
rect 66788 15200 66796 15264
rect 66860 15200 66876 15264
rect 66940 15200 66956 15264
rect 67020 15200 67036 15264
rect 67100 15200 67108 15264
rect 56915 14788 56981 14789
rect 56915 14724 56916 14788
rect 56980 14724 56981 14788
rect 56915 14723 56981 14724
rect 56363 11524 56429 11525
rect 56363 11460 56364 11524
rect 56428 11460 56429 11524
rect 56363 11459 56429 11460
rect 55814 11392 55822 11456
rect 55886 11392 55902 11456
rect 55966 11392 55982 11456
rect 56046 11392 56062 11456
rect 56126 11392 56134 11456
rect 55814 10368 56134 11392
rect 55814 10304 55822 10368
rect 55886 10304 55902 10368
rect 55966 10304 55982 10368
rect 56046 10304 56062 10368
rect 56126 10304 56134 10368
rect 55814 9280 56134 10304
rect 56918 10301 56978 14723
rect 63907 14380 63973 14381
rect 63907 14316 63908 14380
rect 63972 14316 63973 14380
rect 63907 14315 63973 14316
rect 63723 12476 63789 12477
rect 63723 12412 63724 12476
rect 63788 12412 63789 12476
rect 63723 12411 63789 12412
rect 63726 11933 63786 12411
rect 63723 11932 63789 11933
rect 63723 11868 63724 11932
rect 63788 11868 63789 11932
rect 63723 11867 63789 11868
rect 60963 11796 61029 11797
rect 60963 11732 60964 11796
rect 61028 11732 61029 11796
rect 60963 11731 61029 11732
rect 60966 11389 61026 11731
rect 63910 11525 63970 14315
rect 66788 14176 67108 15200
rect 66788 14112 66796 14176
rect 66860 14112 66876 14176
rect 66940 14112 66956 14176
rect 67020 14112 67036 14176
rect 67100 14112 67108 14176
rect 66788 13088 67108 14112
rect 66788 13024 66796 13088
rect 66860 13024 66876 13088
rect 66940 13024 66956 13088
rect 67020 13024 67036 13088
rect 67100 13024 67108 13088
rect 64275 12612 64341 12613
rect 64275 12548 64276 12612
rect 64340 12548 64341 12612
rect 64275 12547 64341 12548
rect 63907 11524 63973 11525
rect 63907 11460 63908 11524
rect 63972 11460 63973 11524
rect 63907 11459 63973 11460
rect 60779 11388 60845 11389
rect 60779 11324 60780 11388
rect 60844 11324 60845 11388
rect 60779 11323 60845 11324
rect 60963 11388 61029 11389
rect 60963 11324 60964 11388
rect 61028 11324 61029 11388
rect 60963 11323 61029 11324
rect 60782 11250 60842 11323
rect 64278 11253 64338 12547
rect 66788 12000 67108 13024
rect 66788 11936 66796 12000
rect 66860 11936 66876 12000
rect 66940 11936 66956 12000
rect 67020 11936 67036 12000
rect 67100 11936 67108 12000
rect 64275 11252 64341 11253
rect 60782 11190 61026 11250
rect 60966 11117 61026 11190
rect 64275 11188 64276 11252
rect 64340 11188 64341 11252
rect 64275 11187 64341 11188
rect 60779 11116 60845 11117
rect 60779 11052 60780 11116
rect 60844 11052 60845 11116
rect 60779 11051 60845 11052
rect 60963 11116 61029 11117
rect 60963 11052 60964 11116
rect 61028 11052 61029 11116
rect 60963 11051 61029 11052
rect 60782 10573 60842 11051
rect 66788 10912 67108 11936
rect 66788 10848 66796 10912
rect 66860 10848 66876 10912
rect 66940 10848 66956 10912
rect 67020 10848 67036 10912
rect 67100 10848 67108 10912
rect 60779 10572 60845 10573
rect 60779 10508 60780 10572
rect 60844 10508 60845 10572
rect 60779 10507 60845 10508
rect 56915 10300 56981 10301
rect 56915 10236 56916 10300
rect 56980 10236 56981 10300
rect 56915 10235 56981 10236
rect 55814 9216 55822 9280
rect 55886 9216 55902 9280
rect 55966 9216 55982 9280
rect 56046 9216 56062 9280
rect 56126 9216 56134 9280
rect 55814 8192 56134 9216
rect 55814 8128 55822 8192
rect 55886 8128 55902 8192
rect 55966 8128 55982 8192
rect 56046 8128 56062 8192
rect 56126 8128 56134 8192
rect 55814 7104 56134 8128
rect 55814 7040 55822 7104
rect 55886 7040 55902 7104
rect 55966 7040 55982 7104
rect 56046 7040 56062 7104
rect 56126 7040 56134 7104
rect 55814 6016 56134 7040
rect 55814 5952 55822 6016
rect 55886 5952 55902 6016
rect 55966 5952 55982 6016
rect 56046 5952 56062 6016
rect 56126 5952 56134 6016
rect 55814 4928 56134 5952
rect 55814 4864 55822 4928
rect 55886 4864 55902 4928
rect 55966 4864 55982 4928
rect 56046 4864 56062 4928
rect 56126 4864 56134 4928
rect 55814 3840 56134 4864
rect 55814 3776 55822 3840
rect 55886 3776 55902 3840
rect 55966 3776 55982 3840
rect 56046 3776 56062 3840
rect 56126 3776 56134 3840
rect 55814 2752 56134 3776
rect 55814 2688 55822 2752
rect 55886 2688 55902 2752
rect 55966 2688 55982 2752
rect 56046 2688 56062 2752
rect 56126 2688 56134 2752
rect 55814 2128 56134 2688
rect 66788 9824 67108 10848
rect 66788 9760 66796 9824
rect 66860 9760 66876 9824
rect 66940 9760 66956 9824
rect 67020 9760 67036 9824
rect 67100 9760 67108 9824
rect 66788 8736 67108 9760
rect 66788 8672 66796 8736
rect 66860 8672 66876 8736
rect 66940 8672 66956 8736
rect 67020 8672 67036 8736
rect 67100 8672 67108 8736
rect 66788 7648 67108 8672
rect 66788 7584 66796 7648
rect 66860 7584 66876 7648
rect 66940 7584 66956 7648
rect 67020 7584 67036 7648
rect 67100 7584 67108 7648
rect 66788 6560 67108 7584
rect 66788 6496 66796 6560
rect 66860 6496 66876 6560
rect 66940 6496 66956 6560
rect 67020 6496 67036 6560
rect 67100 6496 67108 6560
rect 66788 5472 67108 6496
rect 66788 5408 66796 5472
rect 66860 5408 66876 5472
rect 66940 5408 66956 5472
rect 67020 5408 67036 5472
rect 67100 5408 67108 5472
rect 66788 4384 67108 5408
rect 66788 4320 66796 4384
rect 66860 4320 66876 4384
rect 66940 4320 66956 4384
rect 67020 4320 67036 4384
rect 67100 4320 67108 4384
rect 66788 3296 67108 4320
rect 66788 3232 66796 3296
rect 66860 3232 66876 3296
rect 66940 3232 66956 3296
rect 67020 3232 67036 3296
rect 67100 3232 67108 3296
rect 66788 2208 67108 3232
rect 66788 2144 66796 2208
rect 66860 2144 66876 2208
rect 66940 2144 66956 2208
rect 67020 2144 67036 2208
rect 67100 2144 67108 2208
rect 66788 2128 67108 2144
rect 77762 27776 78082 27792
rect 77762 27712 77770 27776
rect 77834 27712 77850 27776
rect 77914 27712 77930 27776
rect 77994 27712 78010 27776
rect 78074 27712 78082 27776
rect 77762 26688 78082 27712
rect 77762 26624 77770 26688
rect 77834 26624 77850 26688
rect 77914 26624 77930 26688
rect 77994 26624 78010 26688
rect 78074 26624 78082 26688
rect 77762 25600 78082 26624
rect 77762 25536 77770 25600
rect 77834 25536 77850 25600
rect 77914 25536 77930 25600
rect 77994 25536 78010 25600
rect 78074 25536 78082 25600
rect 77762 24512 78082 25536
rect 77762 24448 77770 24512
rect 77834 24448 77850 24512
rect 77914 24448 77930 24512
rect 77994 24448 78010 24512
rect 78074 24448 78082 24512
rect 77762 23424 78082 24448
rect 77762 23360 77770 23424
rect 77834 23360 77850 23424
rect 77914 23360 77930 23424
rect 77994 23360 78010 23424
rect 78074 23360 78082 23424
rect 77762 22336 78082 23360
rect 77762 22272 77770 22336
rect 77834 22272 77850 22336
rect 77914 22272 77930 22336
rect 77994 22272 78010 22336
rect 78074 22272 78082 22336
rect 77762 21248 78082 22272
rect 77762 21184 77770 21248
rect 77834 21184 77850 21248
rect 77914 21184 77930 21248
rect 77994 21184 78010 21248
rect 78074 21184 78082 21248
rect 77762 20160 78082 21184
rect 77762 20096 77770 20160
rect 77834 20096 77850 20160
rect 77914 20096 77930 20160
rect 77994 20096 78010 20160
rect 78074 20096 78082 20160
rect 77762 19072 78082 20096
rect 77762 19008 77770 19072
rect 77834 19008 77850 19072
rect 77914 19008 77930 19072
rect 77994 19008 78010 19072
rect 78074 19008 78082 19072
rect 77762 17984 78082 19008
rect 77762 17920 77770 17984
rect 77834 17920 77850 17984
rect 77914 17920 77930 17984
rect 77994 17920 78010 17984
rect 78074 17920 78082 17984
rect 77762 16896 78082 17920
rect 77762 16832 77770 16896
rect 77834 16832 77850 16896
rect 77914 16832 77930 16896
rect 77994 16832 78010 16896
rect 78074 16832 78082 16896
rect 77762 15808 78082 16832
rect 77762 15744 77770 15808
rect 77834 15744 77850 15808
rect 77914 15744 77930 15808
rect 77994 15744 78010 15808
rect 78074 15744 78082 15808
rect 77762 14720 78082 15744
rect 77762 14656 77770 14720
rect 77834 14656 77850 14720
rect 77914 14656 77930 14720
rect 77994 14656 78010 14720
rect 78074 14656 78082 14720
rect 77762 13632 78082 14656
rect 77762 13568 77770 13632
rect 77834 13568 77850 13632
rect 77914 13568 77930 13632
rect 77994 13568 78010 13632
rect 78074 13568 78082 13632
rect 77762 12544 78082 13568
rect 77762 12480 77770 12544
rect 77834 12480 77850 12544
rect 77914 12480 77930 12544
rect 77994 12480 78010 12544
rect 78074 12480 78082 12544
rect 77762 11456 78082 12480
rect 77762 11392 77770 11456
rect 77834 11392 77850 11456
rect 77914 11392 77930 11456
rect 77994 11392 78010 11456
rect 78074 11392 78082 11456
rect 77762 10368 78082 11392
rect 77762 10304 77770 10368
rect 77834 10304 77850 10368
rect 77914 10304 77930 10368
rect 77994 10304 78010 10368
rect 78074 10304 78082 10368
rect 77762 9280 78082 10304
rect 77762 9216 77770 9280
rect 77834 9216 77850 9280
rect 77914 9216 77930 9280
rect 77994 9216 78010 9280
rect 78074 9216 78082 9280
rect 77762 8192 78082 9216
rect 77762 8128 77770 8192
rect 77834 8128 77850 8192
rect 77914 8128 77930 8192
rect 77994 8128 78010 8192
rect 78074 8128 78082 8192
rect 77762 7104 78082 8128
rect 77762 7040 77770 7104
rect 77834 7040 77850 7104
rect 77914 7040 77930 7104
rect 77994 7040 78010 7104
rect 78074 7040 78082 7104
rect 77762 6016 78082 7040
rect 77762 5952 77770 6016
rect 77834 5952 77850 6016
rect 77914 5952 77930 6016
rect 77994 5952 78010 6016
rect 78074 5952 78082 6016
rect 77762 4928 78082 5952
rect 77762 4864 77770 4928
rect 77834 4864 77850 4928
rect 77914 4864 77930 4928
rect 77994 4864 78010 4928
rect 78074 4864 78082 4928
rect 77762 3840 78082 4864
rect 77762 3776 77770 3840
rect 77834 3776 77850 3840
rect 77914 3776 77930 3840
rect 77994 3776 78010 3840
rect 78074 3776 78082 3840
rect 77762 2752 78082 3776
rect 77762 2688 77770 2752
rect 77834 2688 77850 2752
rect 77914 2688 77930 2752
rect 77994 2688 78010 2752
rect 78074 2688 78082 2752
rect 77762 2128 78082 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1649977179
transform 1 0 55936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1649977179
transform 1 0 56580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1649977179
transform -1 0 87860 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1649977179
transform 1 0 2116 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1649977179
transform 1 0 2208 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1649977179
transform 1 0 23368 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1649977179
transform 1 0 52900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1649977179
transform -1 0 87860 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1649977179
transform 1 0 19412 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1649977179
transform -1 0 87308 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1649977179
transform -1 0 86572 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1649977179
transform 1 0 65412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1649977179
transform 1 0 86664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1649977179
transform 1 0 1840 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1649977179
transform -1 0 41400 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1649977179
transform -1 0 87860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1649977179
transform -1 0 87860 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1649977179
transform -1 0 87032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1649977179
transform -1 0 87860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1649977179
transform -1 0 32936 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1649977179
transform 1 0 75072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1649977179
transform 1 0 81328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1649977179
transform 1 0 70748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1649977179
transform 1 0 30820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1649977179
transform 1 0 77004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1649977179
transform 1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1649977179
transform 1 0 81512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1649977179
transform -1 0 87860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1649977179
transform -1 0 87860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1649977179
transform -1 0 87860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1649977179
transform 1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1649977179
transform -1 0 86940 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1649977179
transform -1 0 24012 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1649977179
transform -1 0 23368 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1649977179
transform 1 0 41308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1649977179
transform -1 0 27968 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1649977179
transform 1 0 55936 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1649977179
transform 1 0 70840 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1649977179
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1649977179
transform 1 0 33488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1649977179
transform 1 0 51060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1649977179
transform 1 0 87308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1649977179
transform 1 0 86572 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1649977179
transform 1 0 25944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1649977179
transform 1 0 50232 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1649977179
transform 1 0 48300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1649977179
transform 1 0 55752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1649977179
transform 1 0 19688 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1649977179
transform 1 0 34684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1649977179
transform 1 0 35972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1649977179
transform 1 0 35604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1649977179
transform 1 0 34224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1649977179
transform 1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1649977179
transform 1 0 34224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1649977179
transform 1 0 77096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1649977179
transform 1 0 20792 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1649977179
transform 1 0 63480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1649977179
transform 1 0 84088 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_61
timestamp 1649977179
transform 1 0 78660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_62
timestamp 1649977179
transform 1 0 26772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_63
timestamp 1649977179
transform 1 0 38548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_64
timestamp 1649977179
transform 1 0 27416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_65
timestamp 1649977179
transform 1 0 57040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_66
timestamp 1649977179
transform 1 0 76728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_67
timestamp 1649977179
transform 1 0 38916 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_68
timestamp 1649977179
transform 1 0 24564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_69
timestamp 1649977179
transform 1 0 49312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_70
timestamp 1649977179
transform 1 0 9568 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_71
timestamp 1649977179
transform 1 0 1840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_72
timestamp 1649977179
transform 1 0 58696 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_73
timestamp 1649977179
transform 1 0 79764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_74
timestamp 1649977179
transform 1 0 55568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14
timestamp 1649977179
transform 1 0 2392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25
timestamp 1649977179
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36
timestamp 1649977179
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42
timestamp 1649977179
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71
timestamp 1649977179
transform 1 0 7636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1649977179
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_124
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_155
timestamp 1649977179
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1649977179
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_207
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_211
timestamp 1649977179
transform 1 0 20516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_215
timestamp 1649977179
transform 1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_231
timestamp 1649977179
transform 1 0 22356 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_239
timestamp 1649977179
transform 1 0 23092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1649977179
transform 1 0 23552 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1649977179
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_272
timestamp 1649977179
transform 1 0 26128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_288
timestamp 1649977179
transform 1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1649977179
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_314
timestamp 1649977179
transform 1 0 29992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_320
timestamp 1649977179
transform 1 0 30544 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_328
timestamp 1649977179
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_343
timestamp 1649977179
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1649977179
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_368 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp 1649977179
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_383
timestamp 1649977179
transform 1 0 36340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1649977179
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_398
timestamp 1649977179
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_406
timestamp 1649977179
transform 1 0 38456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1649977179
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_437
timestamp 1649977179
transform 1 0 41308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_441
timestamp 1649977179
transform 1 0 41676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1649977179
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_454
timestamp 1649977179
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_461
timestamp 1649977179
transform 1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_467
timestamp 1649977179
transform 1 0 44068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1649977179
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_482
timestamp 1649977179
transform 1 0 45448 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_490
timestamp 1649977179
transform 1 0 46184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1649977179
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_514
timestamp 1649977179
transform 1 0 48392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_520
timestamp 1649977179
transform 1 0 48944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_524
timestamp 1649977179
transform 1 0 49312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1649977179
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_542
timestamp 1649977179
transform 1 0 50968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_549
timestamp 1649977179
transform 1 0 51612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_555
timestamp 1649977179
transform 1 0 52164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1649977179
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_561
timestamp 1649977179
transform 1 0 52716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_568
timestamp 1649977179
transform 1 0 53360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_576
timestamp 1649977179
transform 1 0 54096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_580
timestamp 1649977179
transform 1 0 54464 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_598
timestamp 1649977179
transform 1 0 56120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_604
timestamp 1649977179
transform 1 0 56672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_610
timestamp 1649977179
transform 1 0 57224 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_626
timestamp 1649977179
transform 1 0 58696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_632
timestamp 1649977179
transform 1 0 59248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_638
timestamp 1649977179
transform 1 0 59800 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_648
timestamp 1649977179
transform 1 0 60720 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_657
timestamp 1649977179
transform 1 0 61548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_664
timestamp 1649977179
transform 1 0 62192 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_673
timestamp 1649977179
transform 1 0 63020 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1649977179
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_704
timestamp 1649977179
transform 1 0 65872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_710
timestamp 1649977179
transform 1 0 66424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_716
timestamp 1649977179
transform 1 0 66976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_722
timestamp 1649977179
transform 1 0 67528 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_732
timestamp 1649977179
transform 1 0 68448 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_741
timestamp 1649977179
transform 1 0 69276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_748
timestamp 1649977179
transform 1 0 69920 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_760
timestamp 1649977179
transform 1 0 71024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_766
timestamp 1649977179
transform 1 0 71576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_772
timestamp 1649977179
transform 1 0 72128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_777
timestamp 1649977179
transform 1 0 72588 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_783
timestamp 1649977179
transform 1 0 73140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_788
timestamp 1649977179
transform 1 0 73600 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_797
timestamp 1649977179
transform 1 0 74428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_805
timestamp 1649977179
transform 1 0 75164 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_811
timestamp 1649977179
transform 1 0 75716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_816
timestamp 1649977179
transform 1 0 76176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_823
timestamp 1649977179
transform 1 0 76820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_827
timestamp 1649977179
transform 1 0 77188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_832
timestamp 1649977179
transform 1 0 77648 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_841
timestamp 1649977179
transform 1 0 78476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_845
timestamp 1649977179
transform 1 0 78844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_853
timestamp 1649977179
transform 1 0 79580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_863
timestamp 1649977179
transform 1 0 80500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_869
timestamp 1649977179
transform 1 0 81052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_874
timestamp 1649977179
transform 1 0 81512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_879
timestamp 1649977179
transform 1 0 81972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_889
timestamp 1649977179
transform 1 0 82892 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_895
timestamp 1649977179
transform 1 0 83444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_900
timestamp 1649977179
transform 1 0 83904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_904
timestamp 1649977179
transform 1 0 84272 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_909
timestamp 1649977179
transform 1 0 84732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_917
timestamp 1649977179
transform 1 0 85468 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_923
timestamp 1649977179
transform 1 0 86020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_928
timestamp 1649977179
transform 1 0 86480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_935
timestamp 1649977179
transform 1 0 87124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_941
timestamp 1649977179
transform 1 0 87676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_948
timestamp 1649977179
transform 1 0 88320 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_7
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_23
timestamp 1649977179
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_29
timestamp 1649977179
transform 1 0 3772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_37
timestamp 1649977179
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_45
timestamp 1649977179
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_66
timestamp 1649977179
transform 1 0 7176 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_78
timestamp 1649977179
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_86
timestamp 1649977179
transform 1 0 9016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_91
timestamp 1649977179
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_97
timestamp 1649977179
transform 1 0 10028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1649977179
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_121
timestamp 1649977179
transform 1 0 12236 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_133
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_139
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_151
timestamp 1649977179
transform 1 0 14996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_200
timestamp 1649977179
transform 1 0 19504 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_204
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_209
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_233
timestamp 1649977179
transform 1 0 22540 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_239
timestamp 1649977179
transform 1 0 23092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_251
timestamp 1649977179
transform 1 0 24196 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_259
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_265
timestamp 1649977179
transform 1 0 25484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_271
timestamp 1649977179
transform 1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1649977179
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_287
timestamp 1649977179
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1649977179
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_315
timestamp 1649977179
transform 1 0 30084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_321
timestamp 1649977179
transform 1 0 30636 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_329
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1649977179
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_358
timestamp 1649977179
transform 1 0 34040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_362
timestamp 1649977179
transform 1 0 34408 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_367
timestamp 1649977179
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_379
timestamp 1649977179
transform 1 0 35972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_409
timestamp 1649977179
transform 1 0 38732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_413
timestamp 1649977179
transform 1 0 39100 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_420
timestamp 1649977179
transform 1 0 39744 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_426
timestamp 1649977179
transform 1 0 40296 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_445
timestamp 1649977179
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_464
timestamp 1649977179
transform 1 0 43792 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_476
timestamp 1649977179
transform 1 0 44896 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_488
timestamp 1649977179
transform 1 0 46000 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_496
timestamp 1649977179
transform 1 0 46736 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_501
timestamp 1649977179
transform 1 0 47196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_524
timestamp 1649977179
transform 1 0 49312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1649977179
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_550
timestamp 1649977179
transform 1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_556
timestamp 1649977179
transform 1 0 52256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1649977179
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_565
timestamp 1649977179
transform 1 0 53084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_573
timestamp 1649977179
transform 1 0 53820 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_577
timestamp 1649977179
transform 1 0 54188 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_589
timestamp 1649977179
transform 1 0 55292 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_596
timestamp 1649977179
transform 1 0 55936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_608
timestamp 1649977179
transform 1 0 57040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_626
timestamp 1649977179
transform 1 0 58696 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_638
timestamp 1649977179
transform 1 0 59800 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_650
timestamp 1649977179
transform 1 0 60904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_656
timestamp 1649977179
transform 1 0 61456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_662
timestamp 1649977179
transform 1 0 62008 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_670
timestamp 1649977179
transform 1 0 62744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_676
timestamp 1649977179
transform 1 0 63296 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_683
timestamp 1649977179
transform 1 0 63940 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_699
timestamp 1649977179
transform 1 0 65412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_711
timestamp 1649977179
transform 1 0 66516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_723
timestamp 1649977179
transform 1 0 67620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1649977179
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1649977179
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_736
timestamp 1649977179
transform 1 0 68816 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_748
timestamp 1649977179
transform 1 0 69920 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_760
timestamp 1649977179
transform 1 0 71024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_767
timestamp 1649977179
transform 1 0 71668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_773
timestamp 1649977179
transform 1 0 72220 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_781
timestamp 1649977179
transform 1 0 72956 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1649977179
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1649977179
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1649977179
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_821
timestamp 1649977179
transform 1 0 76636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_824
timestamp 1649977179
transform 1 0 76912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_828
timestamp 1649977179
transform 1 0 77280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_835
timestamp 1649977179
transform 1 0 77924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1649977179
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_844
timestamp 1649977179
transform 1 0 78752 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_856
timestamp 1649977179
transform 1 0 79856 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_868
timestamp 1649977179
transform 1 0 80960 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_876
timestamp 1649977179
transform 1 0 81696 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_881
timestamp 1649977179
transform 1 0 82156 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_893
timestamp 1649977179
transform 1 0 83260 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1649977179
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1649977179
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_921
timestamp 1649977179
transform 1 0 85836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_925
timestamp 1649977179
transform 1 0 86204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_934
timestamp 1649977179
transform 1 0 87032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_940
timestamp 1649977179
transform 1 0 87584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_6
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_12
timestamp 1649977179
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1649977179
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_258
timestamp 1649977179
transform 1 0 24840 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_266
timestamp 1649977179
transform 1 0 25576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_272
timestamp 1649977179
transform 1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_279
timestamp 1649977179
transform 1 0 26772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_287
timestamp 1649977179
transform 1 0 27508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_298
timestamp 1649977179
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1649977179
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_325
timestamp 1649977179
transform 1 0 31004 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_332
timestamp 1649977179
transform 1 0 31648 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_344
timestamp 1649977179
transform 1 0 32752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_348
timestamp 1649977179
transform 1 0 33120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1649977179
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1649977179
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1649977179
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_497
timestamp 1649977179
transform 1 0 46828 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_509
timestamp 1649977179
transform 1 0 47932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_524
timestamp 1649977179
transform 1 0 49312 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_540
timestamp 1649977179
transform 1 0 50784 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_564
timestamp 1649977179
transform 1 0 52992 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_576
timestamp 1649977179
transform 1 0 54096 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1649977179
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1649977179
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1649977179
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1649977179
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1649977179
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1649977179
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1649977179
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1649977179
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1649977179
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1649977179
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1649977179
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1649977179
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1649977179
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1649977179
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1649977179
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1649977179
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1649977179
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1649977179
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1649977179
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1649977179
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1649977179
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1649977179
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1649977179
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1649977179
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1649977179
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1649977179
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1649977179
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1649977179
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1649977179
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1649977179
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1649977179
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1649977179
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1649977179
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1649977179
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_925
timestamp 1649977179
transform 1 0 86204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_930
timestamp 1649977179
transform 1 0 86664 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_934
timestamp 1649977179
transform 1 0 87032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_939
timestamp 1649977179
transform 1 0 87492 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_946
timestamp 1649977179
transform 1 0 88136 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_528
timestamp 1649977179
transform 1 0 49680 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_540
timestamp 1649977179
transform 1 0 50784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_544
timestamp 1649977179
transform 1 0 51152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_554
timestamp 1649977179
transform 1 0 52072 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_629
timestamp 1649977179
transform 1 0 58972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_633
timestamp 1649977179
transform 1 0 59340 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_640
timestamp 1649977179
transform 1 0 59984 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_652
timestamp 1649977179
transform 1 0 61088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_664
timestamp 1649977179
transform 1 0 62192 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1649977179
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1649977179
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1649977179
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_753
timestamp 1649977179
transform 1 0 70380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_759
timestamp 1649977179
transform 1 0 70932 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_766
timestamp 1649977179
transform 1 0 71576 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_778
timestamp 1649977179
transform 1 0 72680 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1649977179
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1649977179
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1649977179
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1649977179
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1649977179
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1649977179
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1649977179
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1649977179
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1649977179
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1649977179
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1649977179
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1649977179
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1649977179
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1649977179
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_921
timestamp 1649977179
transform 1 0 85836 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_931
timestamp 1649977179
transform 1 0 86756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_936
timestamp 1649977179
transform 1 0 87216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_942
timestamp 1649977179
transform 1 0 87768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_948
timestamp 1649977179
transform 1 0 88320 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6
timestamp 1649977179
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_18
timestamp 1649977179
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1649977179
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_262
timestamp 1649977179
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_268
timestamp 1649977179
transform 1 0 25760 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_291
timestamp 1649977179
transform 1 0 27876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 1649977179
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_341
timestamp 1649977179
transform 1 0 32476 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_349
timestamp 1649977179
transform 1 0 33212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp 1649977179
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_594
timestamp 1649977179
transform 1 0 55752 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_598
timestamp 1649977179
transform 1 0 56120 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_610
timestamp 1649977179
transform 1 0 57224 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_622
timestamp 1649977179
transform 1 0 58328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_634
timestamp 1649977179
transform 1 0 59432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_642
timestamp 1649977179
transform 1 0 60168 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1649977179
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1649977179
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1649977179
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1649977179
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1649977179
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1649977179
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1649977179
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1649977179
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1649977179
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1649977179
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1649977179
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1649977179
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1649977179
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1649977179
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1649977179
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1649977179
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1649977179
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1649977179
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1649977179
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1649977179
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1649977179
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1649977179
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1649977179
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1649977179
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1649977179
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1649977179
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1649977179
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1649977179
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_937
timestamp 1649977179
transform 1 0 87308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_943
timestamp 1649977179
transform 1 0 87860 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_948
timestamp 1649977179
transform 1 0 88320 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_260
timestamp 1649977179
transform 1 0 25024 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_272
timestamp 1649977179
transform 1 0 26128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_286
timestamp 1649977179
transform 1 0 27416 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_290
timestamp 1649977179
transform 1 0 27784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_302
timestamp 1649977179
transform 1 0 28888 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_310
timestamp 1649977179
transform 1 0 29624 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_318
timestamp 1649977179
transform 1 0 30360 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_330
timestamp 1649977179
transform 1 0 31464 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1649977179
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1649977179
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1649977179
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1649977179
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1649977179
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1649977179
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1649977179
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1649977179
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1649977179
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1649977179
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1649977179
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1649977179
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1649977179
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1649977179
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1649977179
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1649977179
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1649977179
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1649977179
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1649977179
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1649977179
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1649977179
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1649977179
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1649977179
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1649977179
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1649977179
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1649977179
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_933
timestamp 1649977179
transform 1 0 86940 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_943
timestamp 1649977179
transform 1 0 87860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_948
timestamp 1649977179
transform 1 0 88320 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6
timestamp 1649977179
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_18
timestamp 1649977179
transform 1 0 2760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1649977179
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_262
timestamp 1649977179
transform 1 0 25208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_266
timestamp 1649977179
transform 1 0 25576 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_284
timestamp 1649977179
transform 1 0 27232 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_296
timestamp 1649977179
transform 1 0 28336 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_605
timestamp 1649977179
transform 1 0 56764 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_616
timestamp 1649977179
transform 1 0 57776 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_628
timestamp 1649977179
transform 1 0 58880 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_640
timestamp 1649977179
transform 1 0 59984 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1649977179
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1649977179
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1649977179
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1649977179
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1649977179
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1649977179
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1649977179
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1649977179
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1649977179
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1649977179
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1649977179
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1649977179
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1649977179
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1649977179
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1649977179
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1649977179
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1649977179
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1649977179
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1649977179
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1649977179
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1649977179
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1649977179
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_937
timestamp 1649977179
transform 1 0 87308 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_943
timestamp 1649977179
transform 1 0 87860 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_948
timestamp 1649977179
transform 1 0 88320 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_12
timestamp 1649977179
transform 1 0 2208 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_24
timestamp 1649977179
transform 1 0 3312 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_36
timestamp 1649977179
transform 1 0 4416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1649977179
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_593
timestamp 1649977179
transform 1 0 55660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_613
timestamp 1649977179
transform 1 0 57500 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1649977179
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1649977179
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1649977179
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1649977179
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1649977179
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1649977179
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1649977179
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1649977179
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1649977179
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1649977179
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1649977179
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1649977179
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1649977179
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1649977179
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1649977179
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1649977179
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1649977179
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1649977179
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1649977179
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1649977179
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1649977179
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_933
timestamp 1649977179
transform 1 0 86940 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_937
timestamp 1649977179
transform 1 0 87308 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_948
timestamp 1649977179
transform 1 0 88320 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_269
timestamp 1649977179
transform 1 0 25852 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_276
timestamp 1649977179
transform 1 0 26496 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_288
timestamp 1649977179
transform 1 0 27600 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_300
timestamp 1649977179
transform 1 0 28704 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_409
timestamp 1649977179
transform 1 0 38732 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_416
timestamp 1649977179
transform 1 0 39376 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_606
timestamp 1649977179
transform 1 0 56856 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_618
timestamp 1649977179
transform 1 0 57960 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_630
timestamp 1649977179
transform 1 0 59064 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_642
timestamp 1649977179
transform 1 0 60168 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1649977179
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1649977179
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1649977179
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1649977179
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1649977179
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1649977179
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1649977179
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1649977179
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1649977179
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1649977179
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1649977179
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1649977179
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1649977179
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1649977179
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1649977179
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1649977179
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1649977179
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1649977179
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1649977179
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1649977179
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1649977179
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1649977179
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1649977179
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_949
timestamp 1649977179
transform 1 0 88412 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6
timestamp 1649977179
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_18
timestamp 1649977179
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_30
timestamp 1649977179
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_42
timestamp 1649977179
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_411
timestamp 1649977179
transform 1 0 38916 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_432
timestamp 1649977179
transform 1 0 40848 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_444
timestamp 1649977179
transform 1 0 41952 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1649977179
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1649977179
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1649977179
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1649977179
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1649977179
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1649977179
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1649977179
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1649977179
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_821
timestamp 1649977179
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1649977179
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1649977179
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1649977179
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1649977179
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_865
timestamp 1649977179
transform 1 0 80684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_877
timestamp 1649977179
transform 1 0 81788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_889
timestamp 1649977179
transform 1 0 82892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_895
timestamp 1649977179
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1649977179
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1649977179
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_921
timestamp 1649977179
transform 1 0 85836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_933
timestamp 1649977179
transform 1 0 86940 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_941
timestamp 1649977179
transform 1 0 87676 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_948
timestamp 1649977179
transform 1 0 88320 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_444
timestamp 1649977179
transform 1 0 41952 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_456
timestamp 1649977179
transform 1 0 43056 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_468
timestamp 1649977179
transform 1 0 44160 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_496
timestamp 1649977179
transform 1 0 46736 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_508
timestamp 1649977179
transform 1 0 47840 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_520
timestamp 1649977179
transform 1 0 48944 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1649977179
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1649977179
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1649977179
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1649977179
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1649977179
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1649977179
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1649977179
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1649977179
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1649977179
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_813
timestamp 1649977179
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_825
timestamp 1649977179
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_837
timestamp 1649977179
transform 1 0 78108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_849
timestamp 1649977179
transform 1 0 79212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_861
timestamp 1649977179
transform 1 0 80316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_867
timestamp 1649977179
transform 1 0 80868 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_869
timestamp 1649977179
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_881
timestamp 1649977179
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_893
timestamp 1649977179
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_905
timestamp 1649977179
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_917
timestamp 1649977179
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_923
timestamp 1649977179
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_925
timestamp 1649977179
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_937
timestamp 1649977179
transform 1 0 87308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_943
timestamp 1649977179
transform 1 0 87860 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_948
timestamp 1649977179
transform 1 0 88320 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_13
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_25
timestamp 1649977179
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_37
timestamp 1649977179
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1649977179
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_404
timestamp 1649977179
transform 1 0 38272 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_416
timestamp 1649977179
transform 1 0 39376 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_428
timestamp 1649977179
transform 1 0 40480 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_436
timestamp 1649977179
transform 1 0 41216 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_443
timestamp 1649977179
transform 1 0 41860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_462
timestamp 1649977179
transform 1 0 43608 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_474
timestamp 1649977179
transform 1 0 44712 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_486
timestamp 1649977179
transform 1 0 45816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_498
timestamp 1649977179
transform 1 0 46920 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_521
timestamp 1649977179
transform 1 0 49036 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_531
timestamp 1649977179
transform 1 0 49956 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_537
timestamp 1649977179
transform 1 0 50508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_549
timestamp 1649977179
transform 1 0 51612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_557
timestamp 1649977179
transform 1 0 52348 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_570
timestamp 1649977179
transform 1 0 53544 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_582
timestamp 1649977179
transform 1 0 54648 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_594
timestamp 1649977179
transform 1 0 55752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_606
timestamp 1649977179
transform 1 0 56856 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1649977179
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1649977179
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1649977179
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1649977179
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1649977179
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1649977179
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1649977179
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1649977179
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1649977179
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1649977179
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_821
timestamp 1649977179
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1649977179
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1649977179
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_841
timestamp 1649977179
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_853
timestamp 1649977179
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_865
timestamp 1649977179
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_877
timestamp 1649977179
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1649977179
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1649977179
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_897
timestamp 1649977179
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_909
timestamp 1649977179
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_921
timestamp 1649977179
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_933
timestamp 1649977179
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_948
timestamp 1649977179
transform 1 0 88320 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_6
timestamp 1649977179
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_18
timestamp 1649977179
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_381
timestamp 1649977179
transform 1 0 36156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_391
timestamp 1649977179
transform 1 0 37076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_400
timestamp 1649977179
transform 1 0 37904 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_411
timestamp 1649977179
transform 1 0 38916 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_449
timestamp 1649977179
transform 1 0 42412 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_468
timestamp 1649977179
transform 1 0 44160 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_485
timestamp 1649977179
transform 1 0 45724 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_508
timestamp 1649977179
transform 1 0 47840 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_520
timestamp 1649977179
transform 1 0 48944 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_552
timestamp 1649977179
transform 1 0 51888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_558
timestamp 1649977179
transform 1 0 52440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_577
timestamp 1649977179
transform 1 0 54188 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_585
timestamp 1649977179
transform 1 0 54924 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_592
timestamp 1649977179
transform 1 0 55568 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_604
timestamp 1649977179
transform 1 0 56672 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_616
timestamp 1649977179
transform 1 0 57776 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_628
timestamp 1649977179
transform 1 0 58880 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_640
timestamp 1649977179
transform 1 0 59984 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_738
timestamp 1649977179
transform 1 0 69000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_750
timestamp 1649977179
transform 1 0 70104 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1649977179
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1649977179
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1649977179
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1649977179
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1649977179
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1649977179
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_813
timestamp 1649977179
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_825
timestamp 1649977179
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_837
timestamp 1649977179
transform 1 0 78108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_849
timestamp 1649977179
transform 1 0 79212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_861
timestamp 1649977179
transform 1 0 80316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_867
timestamp 1649977179
transform 1 0 80868 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_869
timestamp 1649977179
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_881
timestamp 1649977179
transform 1 0 82156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_893
timestamp 1649977179
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_905
timestamp 1649977179
transform 1 0 84364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1649977179
transform 1 0 85468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1649977179
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_925
timestamp 1649977179
transform 1 0 86204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_937
timestamp 1649977179
transform 1 0 87308 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_948
timestamp 1649977179
transform 1 0 88320 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_320
timestamp 1649977179
transform 1 0 30544 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1649977179
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_345
timestamp 1649977179
transform 1 0 32844 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_357
timestamp 1649977179
transform 1 0 33948 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_369
timestamp 1649977179
transform 1 0 35052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_386
timestamp 1649977179
transform 1 0 36616 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_399
timestamp 1649977179
transform 1 0 37812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_423
timestamp 1649977179
transform 1 0 40020 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_442
timestamp 1649977179
transform 1 0 41768 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_456
timestamp 1649977179
transform 1 0 43056 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_468
timestamp 1649977179
transform 1 0 44160 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_476
timestamp 1649977179
transform 1 0 44896 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_481
timestamp 1649977179
transform 1 0 45356 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_501
timestamp 1649977179
transform 1 0 47196 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_524
timestamp 1649977179
transform 1 0 49312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_543
timestamp 1649977179
transform 1 0 51060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_549
timestamp 1649977179
transform 1 0 51612 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_557
timestamp 1649977179
transform 1 0 52348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_577
timestamp 1649977179
transform 1 0 54188 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_583
timestamp 1649977179
transform 1 0 54740 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_595
timestamp 1649977179
transform 1 0 55844 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_607
timestamp 1649977179
transform 1 0 56948 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_611
timestamp 1649977179
transform 1 0 57316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_633
timestamp 1649977179
transform 1 0 59340 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_650
timestamp 1649977179
transform 1 0 60904 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_662
timestamp 1649977179
transform 1 0 62008 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_670
timestamp 1649977179
transform 1 0 62744 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_691
timestamp 1649977179
transform 1 0 64676 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_703
timestamp 1649977179
transform 1 0 65780 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_715
timestamp 1649977179
transform 1 0 66884 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_732
timestamp 1649977179
transform 1 0 68448 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_754
timestamp 1649977179
transform 1 0 70472 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_766
timestamp 1649977179
transform 1 0 71576 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_778
timestamp 1649977179
transform 1 0 72680 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1649977179
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1649977179
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1649977179
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_821
timestamp 1649977179
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1649977179
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1649977179
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_841
timestamp 1649977179
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_853
timestamp 1649977179
transform 1 0 79580 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_865
timestamp 1649977179
transform 1 0 80684 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_877
timestamp 1649977179
transform 1 0 81788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_889
timestamp 1649977179
transform 1 0 82892 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_895
timestamp 1649977179
transform 1 0 83444 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_897
timestamp 1649977179
transform 1 0 83628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_909
timestamp 1649977179
transform 1 0 84732 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_921
timestamp 1649977179
transform 1 0 85836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_933
timestamp 1649977179
transform 1 0 86940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_945
timestamp 1649977179
transform 1 0 88044 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_6
timestamp 1649977179
transform 1 0 1656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_18
timestamp 1649977179
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_259
timestamp 1649977179
transform 1 0 24932 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_263
timestamp 1649977179
transform 1 0 25300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_275
timestamp 1649977179
transform 1 0 26404 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_287
timestamp 1649977179
transform 1 0 27508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_299
timestamp 1649977179
transform 1 0 28612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1649977179
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_326
timestamp 1649977179
transform 1 0 31096 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_338
timestamp 1649977179
transform 1 0 32200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_368
timestamp 1649977179
transform 1 0 34960 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_376
timestamp 1649977179
transform 1 0 35696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_380
timestamp 1649977179
transform 1 0 36064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_404
timestamp 1649977179
transform 1 0 38272 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1649977179
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_427
timestamp 1649977179
transform 1 0 40388 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_463
timestamp 1649977179
transform 1 0 43700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_496
timestamp 1649977179
transform 1 0 46736 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_504
timestamp 1649977179
transform 1 0 47472 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_516
timestamp 1649977179
transform 1 0 48576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_523
timestamp 1649977179
transform 1 0 49220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_529
timestamp 1649977179
transform 1 0 49772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_542
timestamp 1649977179
transform 1 0 50968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_548
timestamp 1649977179
transform 1 0 51520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_552
timestamp 1649977179
transform 1 0 51888 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_573
timestamp 1649977179
transform 1 0 53820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_585
timestamp 1649977179
transform 1 0 54924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_605
timestamp 1649977179
transform 1 0 56764 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_611
timestamp 1649977179
transform 1 0 57316 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_621
timestamp 1649977179
transform 1 0 58236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_628
timestamp 1649977179
transform 1 0 58880 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_635
timestamp 1649977179
transform 1 0 59524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_641
timestamp 1649977179
transform 1 0 60076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_654
timestamp 1649977179
transform 1 0 61272 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_660
timestamp 1649977179
transform 1 0 61824 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_666
timestamp 1649977179
transform 1 0 62376 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_678
timestamp 1649977179
transform 1 0 63480 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_686
timestamp 1649977179
transform 1 0 64216 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_694
timestamp 1649977179
transform 1 0 64952 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1649977179
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1649977179
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1649977179
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1649977179
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1649977179
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1649977179
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1649977179
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1649977179
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1649977179
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_813
timestamp 1649977179
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_825
timestamp 1649977179
transform 1 0 77004 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_837
timestamp 1649977179
transform 1 0 78108 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_849
timestamp 1649977179
transform 1 0 79212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_861
timestamp 1649977179
transform 1 0 80316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_867
timestamp 1649977179
transform 1 0 80868 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_869
timestamp 1649977179
transform 1 0 81052 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_881
timestamp 1649977179
transform 1 0 82156 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_893
timestamp 1649977179
transform 1 0 83260 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_905
timestamp 1649977179
transform 1 0 84364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_917
timestamp 1649977179
transform 1 0 85468 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_923
timestamp 1649977179
transform 1 0 86020 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_925
timestamp 1649977179
transform 1 0 86204 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_937
timestamp 1649977179
transform 1 0 87308 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_949
timestamp 1649977179
transform 1 0 88412 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_6
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_18
timestamp 1649977179
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_30
timestamp 1649977179
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_42
timestamp 1649977179
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_262
timestamp 1649977179
transform 1 0 25208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_266
timestamp 1649977179
transform 1 0 25576 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_296
timestamp 1649977179
transform 1 0 28336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_308
timestamp 1649977179
transform 1 0 29440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 1649977179
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_345
timestamp 1649977179
transform 1 0 32844 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_350
timestamp 1649977179
transform 1 0 33304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_357
timestamp 1649977179
transform 1 0 33948 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_363
timestamp 1649977179
transform 1 0 34500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_375
timestamp 1649977179
transform 1 0 35604 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_379
timestamp 1649977179
transform 1 0 35972 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1649977179
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_403
timestamp 1649977179
transform 1 0 38180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_407
timestamp 1649977179
transform 1 0 38548 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_427
timestamp 1649977179
transform 1 0 40388 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_434
timestamp 1649977179
transform 1 0 41032 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1649977179
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_456
timestamp 1649977179
transform 1 0 43056 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_463
timestamp 1649977179
transform 1 0 43700 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_472
timestamp 1649977179
transform 1 0 44528 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_482
timestamp 1649977179
transform 1 0 45448 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_501
timestamp 1649977179
transform 1 0 47196 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1649977179
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_516
timestamp 1649977179
transform 1 0 48576 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_537
timestamp 1649977179
transform 1 0 50508 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_545
timestamp 1649977179
transform 1 0 51244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_557
timestamp 1649977179
transform 1 0 52348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_564
timestamp 1649977179
transform 1 0 52992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_570
timestamp 1649977179
transform 1 0 53544 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_578
timestamp 1649977179
transform 1 0 54280 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_595
timestamp 1649977179
transform 1 0 55844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_601
timestamp 1649977179
transform 1 0 56396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_607
timestamp 1649977179
transform 1 0 56948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_613
timestamp 1649977179
transform 1 0 57500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_621
timestamp 1649977179
transform 1 0 58236 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_637
timestamp 1649977179
transform 1 0 59708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_658
timestamp 1649977179
transform 1 0 61640 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_662
timestamp 1649977179
transform 1 0 62008 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_666
timestamp 1649977179
transform 1 0 62376 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_678
timestamp 1649977179
transform 1 0 63480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_697
timestamp 1649977179
transform 1 0 65228 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_716
timestamp 1649977179
transform 1 0 66976 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1649977179
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1649977179
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1649977179
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1649977179
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1649977179
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1649977179
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1649977179
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1649977179
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_821
timestamp 1649977179
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1649977179
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1649977179
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_841
timestamp 1649977179
transform 1 0 78476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_853
timestamp 1649977179
transform 1 0 79580 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_865
timestamp 1649977179
transform 1 0 80684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_877
timestamp 1649977179
transform 1 0 81788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_889
timestamp 1649977179
transform 1 0 82892 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_895
timestamp 1649977179
transform 1 0 83444 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_897
timestamp 1649977179
transform 1 0 83628 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_909
timestamp 1649977179
transform 1 0 84732 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_921
timestamp 1649977179
transform 1 0 85836 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_933
timestamp 1649977179
transform 1 0 86940 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_943
timestamp 1649977179
transform 1 0 87860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_948
timestamp 1649977179
transform 1 0 88320 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_6
timestamp 1649977179
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1649977179
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_158
timestamp 1649977179
transform 1 0 15640 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_170
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_182
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_259
timestamp 1649977179
transform 1 0 24932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_285
timestamp 1649977179
transform 1 0 27324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_291
timestamp 1649977179
transform 1 0 27876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_299
timestamp 1649977179
transform 1 0 28612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1649977179
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_325
timestamp 1649977179
transform 1 0 31004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_338
timestamp 1649977179
transform 1 0 32200 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_344
timestamp 1649977179
transform 1 0 32752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1649977179
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_370
timestamp 1649977179
transform 1 0 35144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_374
timestamp 1649977179
transform 1 0 35512 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_381
timestamp 1649977179
transform 1 0 36156 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_385
timestamp 1649977179
transform 1 0 36524 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_396
timestamp 1649977179
transform 1 0 37536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_406
timestamp 1649977179
transform 1 0 38456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_416
timestamp 1649977179
transform 1 0 39376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_427
timestamp 1649977179
transform 1 0 40388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_438
timestamp 1649977179
transform 1 0 41400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_451
timestamp 1649977179
transform 1 0 42596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_463
timestamp 1649977179
transform 1 0 43700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_467
timestamp 1649977179
transform 1 0 44068 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_473
timestamp 1649977179
transform 1 0 44620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_480
timestamp 1649977179
transform 1 0 45264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_490
timestamp 1649977179
transform 1 0 46184 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_499
timestamp 1649977179
transform 1 0 47012 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_506
timestamp 1649977179
transform 1 0 47656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_518
timestamp 1649977179
transform 1 0 48760 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_524
timestamp 1649977179
transform 1 0 49312 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_529
timestamp 1649977179
transform 1 0 49772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_541
timestamp 1649977179
transform 1 0 50876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_560
timestamp 1649977179
transform 1 0 52624 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_570
timestamp 1649977179
transform 1 0 53544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_582
timestamp 1649977179
transform 1 0 54648 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_592
timestamp 1649977179
transform 1 0 55568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_599
timestamp 1649977179
transform 1 0 56212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_619
timestamp 1649977179
transform 1 0 58052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_638
timestamp 1649977179
transform 1 0 59800 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_648
timestamp 1649977179
transform 1 0 60720 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_660
timestamp 1649977179
transform 1 0 61824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_664
timestamp 1649977179
transform 1 0 62192 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_675
timestamp 1649977179
transform 1 0 63204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_683
timestamp 1649977179
transform 1 0 63940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_692
timestamp 1649977179
transform 1 0 64768 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_722
timestamp 1649977179
transform 1 0 67528 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_741
timestamp 1649977179
transform 1 0 69276 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_753
timestamp 1649977179
transform 1 0 70380 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1649977179
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1649977179
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1649977179
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1649977179
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1649977179
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1649977179
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_813
timestamp 1649977179
transform 1 0 75900 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_825
timestamp 1649977179
transform 1 0 77004 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_837
timestamp 1649977179
transform 1 0 78108 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_849
timestamp 1649977179
transform 1 0 79212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_861
timestamp 1649977179
transform 1 0 80316 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_867
timestamp 1649977179
transform 1 0 80868 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_869
timestamp 1649977179
transform 1 0 81052 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_881
timestamp 1649977179
transform 1 0 82156 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_893
timestamp 1649977179
transform 1 0 83260 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_905
timestamp 1649977179
transform 1 0 84364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_917
timestamp 1649977179
transform 1 0 85468 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_923
timestamp 1649977179
transform 1 0 86020 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_925
timestamp 1649977179
transform 1 0 86204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_937
timestamp 1649977179
transform 1 0 87308 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_948
timestamp 1649977179
transform 1 0 88320 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_6
timestamp 1649977179
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_18
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_30
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_42
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_196
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_207
timestamp 1649977179
transform 1 0 20148 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1649977179
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_256
timestamp 1649977179
transform 1 0 24656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_265
timestamp 1649977179
transform 1 0 25484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1649977179
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_300
timestamp 1649977179
transform 1 0 28704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_315
timestamp 1649977179
transform 1 0 30084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_326
timestamp 1649977179
transform 1 0 31096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1649977179
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_344
timestamp 1649977179
transform 1 0 32752 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_366
timestamp 1649977179
transform 1 0 34776 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_372
timestamp 1649977179
transform 1 0 35328 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_379
timestamp 1649977179
transform 1 0 35972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_389
timestamp 1649977179
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_397
timestamp 1649977179
transform 1 0 37628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_410
timestamp 1649977179
transform 1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_420
timestamp 1649977179
transform 1 0 39744 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_428
timestamp 1649977179
transform 1 0 40480 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_434
timestamp 1649977179
transform 1 0 41032 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_445
timestamp 1649977179
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_472
timestamp 1649977179
transform 1 0 44528 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_491
timestamp 1649977179
transform 1 0 46276 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_500
timestamp 1649977179
transform 1 0 47104 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_511
timestamp 1649977179
transform 1 0 48116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_523
timestamp 1649977179
transform 1 0 49220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_532
timestamp 1649977179
transform 1 0 50048 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_551
timestamp 1649977179
transform 1 0 51796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_557
timestamp 1649977179
transform 1 0 52348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_567
timestamp 1649977179
transform 1 0 53268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_576
timestamp 1649977179
transform 1 0 54096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_580
timestamp 1649977179
transform 1 0 54464 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_592
timestamp 1649977179
transform 1 0 55568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_598
timestamp 1649977179
transform 1 0 56120 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_613
timestamp 1649977179
transform 1 0 57500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_622
timestamp 1649977179
transform 1 0 58328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_633
timestamp 1649977179
transform 1 0 59340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_642
timestamp 1649977179
transform 1 0 60168 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_648
timestamp 1649977179
transform 1 0 60720 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_685
timestamp 1649977179
transform 1 0 64124 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_692
timestamp 1649977179
transform 1 0 64768 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_704
timestamp 1649977179
transform 1 0 65872 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_712
timestamp 1649977179
transform 1 0 66608 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_718
timestamp 1649977179
transform 1 0 67160 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_726
timestamp 1649977179
transform 1 0 67896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_734
timestamp 1649977179
transform 1 0 68632 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_756
timestamp 1649977179
transform 1 0 70656 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_760
timestamp 1649977179
transform 1 0 71024 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_771
timestamp 1649977179
transform 1 0 72036 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1649977179
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1649977179
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1649977179
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_809
timestamp 1649977179
transform 1 0 75532 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_821
timestamp 1649977179
transform 1 0 76636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_833
timestamp 1649977179
transform 1 0 77740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_839
timestamp 1649977179
transform 1 0 78292 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_841
timestamp 1649977179
transform 1 0 78476 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_853
timestamp 1649977179
transform 1 0 79580 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_865
timestamp 1649977179
transform 1 0 80684 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_877
timestamp 1649977179
transform 1 0 81788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_889
timestamp 1649977179
transform 1 0 82892 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_895
timestamp 1649977179
transform 1 0 83444 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_897
timestamp 1649977179
transform 1 0 83628 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_909
timestamp 1649977179
transform 1 0 84732 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_921
timestamp 1649977179
transform 1 0 85836 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_933
timestamp 1649977179
transform 1 0 86940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_948
timestamp 1649977179
transform 1 0 88320 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_210
timestamp 1649977179
transform 1 0 20424 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_220
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_232
timestamp 1649977179
transform 1 0 22448 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_244
timestamp 1649977179
transform 1 0 23552 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_281
timestamp 1649977179
transform 1 0 26956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1649977179
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_325
timestamp 1649977179
transform 1 0 31004 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_334
timestamp 1649977179
transform 1 0 31832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_343
timestamp 1649977179
transform 1 0 32660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_347
timestamp 1649977179
transform 1 0 33028 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_353
timestamp 1649977179
transform 1 0 33580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 1649977179
transform 1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_372
timestamp 1649977179
transform 1 0 35328 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_380
timestamp 1649977179
transform 1 0 36064 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_398
timestamp 1649977179
transform 1 0 37720 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_417
timestamp 1649977179
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_430
timestamp 1649977179
transform 1 0 40664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_449
timestamp 1649977179
transform 1 0 42412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_462
timestamp 1649977179
transform 1 0 43608 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_471
timestamp 1649977179
transform 1 0 44436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_487
timestamp 1649977179
transform 1 0 45908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_498
timestamp 1649977179
transform 1 0 46920 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_506
timestamp 1649977179
transform 1 0 47656 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_511
timestamp 1649977179
transform 1 0 48116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_517
timestamp 1649977179
transform 1 0 48668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_529
timestamp 1649977179
transform 1 0 49772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_543
timestamp 1649977179
transform 1 0 51060 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_565
timestamp 1649977179
transform 1 0 53084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_572
timestamp 1649977179
transform 1 0 53728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_579
timestamp 1649977179
transform 1 0 54372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_585
timestamp 1649977179
transform 1 0 54924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_607
timestamp 1649977179
transform 1 0 56948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_616
timestamp 1649977179
transform 1 0 57776 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_628
timestamp 1649977179
transform 1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_641
timestamp 1649977179
transform 1 0 60076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_661
timestamp 1649977179
transform 1 0 61916 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_676
timestamp 1649977179
transform 1 0 63296 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_682
timestamp 1649977179
transform 1 0 63848 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_690
timestamp 1649977179
transform 1 0 64584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_697
timestamp 1649977179
transform 1 0 65228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_708
timestamp 1649977179
transform 1 0 66240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_727
timestamp 1649977179
transform 1 0 67988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_738
timestamp 1649977179
transform 1 0 69000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_746
timestamp 1649977179
transform 1 0 69736 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_753
timestamp 1649977179
transform 1 0 70380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_773
timestamp 1649977179
transform 1 0 72220 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_779
timestamp 1649977179
transform 1 0 72772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_791
timestamp 1649977179
transform 1 0 73876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_803
timestamp 1649977179
transform 1 0 74980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 1649977179
transform 1 0 75716 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_813
timestamp 1649977179
transform 1 0 75900 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_825
timestamp 1649977179
transform 1 0 77004 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_837
timestamp 1649977179
transform 1 0 78108 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_849
timestamp 1649977179
transform 1 0 79212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_861
timestamp 1649977179
transform 1 0 80316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_867
timestamp 1649977179
transform 1 0 80868 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_869
timestamp 1649977179
transform 1 0 81052 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_881
timestamp 1649977179
transform 1 0 82156 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_893
timestamp 1649977179
transform 1 0 83260 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_905
timestamp 1649977179
transform 1 0 84364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_917
timestamp 1649977179
transform 1 0 85468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_923
timestamp 1649977179
transform 1 0 86020 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_925
timestamp 1649977179
transform 1 0 86204 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_937
timestamp 1649977179
transform 1 0 87308 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_949
timestamp 1649977179
transform 1 0 88412 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_25
timestamp 1649977179
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_37
timestamp 1649977179
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_196
timestamp 1649977179
transform 1 0 19136 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_202
timestamp 1649977179
transform 1 0 19688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_209
timestamp 1649977179
transform 1 0 20332 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1649977179
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_250
timestamp 1649977179
transform 1 0 24104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_256
timestamp 1649977179
transform 1 0 24656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_265
timestamp 1649977179
transform 1 0 25484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1649977179
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1649977179
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_288
timestamp 1649977179
transform 1 0 27600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_296
timestamp 1649977179
transform 1 0 28336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_320
timestamp 1649977179
transform 1 0 30544 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_326
timestamp 1649977179
transform 1 0 31096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1649977179
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_344
timestamp 1649977179
transform 1 0 32752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_351
timestamp 1649977179
transform 1 0 33396 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_360
timestamp 1649977179
transform 1 0 34224 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_370
timestamp 1649977179
transform 1 0 35144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_381
timestamp 1649977179
transform 1 0 36156 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1649977179
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_403
timestamp 1649977179
transform 1 0 38180 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_409
timestamp 1649977179
transform 1 0 38732 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_432
timestamp 1649977179
transform 1 0 40848 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_436
timestamp 1649977179
transform 1 0 41216 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_443
timestamp 1649977179
transform 1 0 41860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_459
timestamp 1649977179
transform 1 0 43332 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_469
timestamp 1649977179
transform 1 0 44252 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_476
timestamp 1649977179
transform 1 0 44896 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_480
timestamp 1649977179
transform 1 0 45264 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_488
timestamp 1649977179
transform 1 0 46000 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_500
timestamp 1649977179
transform 1 0 47104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_514
timestamp 1649977179
transform 1 0 48392 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_521
timestamp 1649977179
transform 1 0 49036 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_545
timestamp 1649977179
transform 1 0 51244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_555
timestamp 1649977179
transform 1 0 52164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_567
timestamp 1649977179
transform 1 0 53268 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_574
timestamp 1649977179
transform 1 0 53912 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_580
timestamp 1649977179
transform 1 0 54464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_601
timestamp 1649977179
transform 1 0 56396 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_611
timestamp 1649977179
transform 1 0 57316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_627
timestamp 1649977179
transform 1 0 58788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_634
timestamp 1649977179
transform 1 0 59432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_658
timestamp 1649977179
transform 1 0 61640 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_667
timestamp 1649977179
transform 1 0 62468 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_689
timestamp 1649977179
transform 1 0 64492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_699
timestamp 1649977179
transform 1 0 65412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_707
timestamp 1649977179
transform 1 0 66148 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_715
timestamp 1649977179
transform 1 0 66884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_724
timestamp 1649977179
transform 1 0 67712 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_729
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_736
timestamp 1649977179
transform 1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_744
timestamp 1649977179
transform 1 0 69552 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_763
timestamp 1649977179
transform 1 0 71300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_771
timestamp 1649977179
transform 1 0 72036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 1649977179
transform 1 0 72588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1649977179
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1649977179
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_797
timestamp 1649977179
transform 1 0 74428 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_809
timestamp 1649977179
transform 1 0 75532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_821
timestamp 1649977179
transform 1 0 76636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_833
timestamp 1649977179
transform 1 0 77740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_839
timestamp 1649977179
transform 1 0 78292 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_841
timestamp 1649977179
transform 1 0 78476 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_853
timestamp 1649977179
transform 1 0 79580 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_865
timestamp 1649977179
transform 1 0 80684 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_877
timestamp 1649977179
transform 1 0 81788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_889
timestamp 1649977179
transform 1 0 82892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_895
timestamp 1649977179
transform 1 0 83444 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_897
timestamp 1649977179
transform 1 0 83628 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_909
timestamp 1649977179
transform 1 0 84732 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_921
timestamp 1649977179
transform 1 0 85836 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_929
timestamp 1649977179
transform 1 0 86572 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_934
timestamp 1649977179
transform 1 0 87032 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_942
timestamp 1649977179
transform 1 0 87768 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_948
timestamp 1649977179
transform 1 0 88320 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_6
timestamp 1649977179
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1649977179
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1649977179
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_154
timestamp 1649977179
transform 1 0 15272 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_166
timestamp 1649977179
transform 1 0 16376 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_182
timestamp 1649977179
transform 1 0 17848 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1649977179
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_206
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_214
timestamp 1649977179
transform 1 0 20792 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_242
timestamp 1649977179
transform 1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1649977179
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_257
timestamp 1649977179
transform 1 0 24748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_263
timestamp 1649977179
transform 1 0 25300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_273
timestamp 1649977179
transform 1 0 26220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_284
timestamp 1649977179
transform 1 0 27232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_293
timestamp 1649977179
transform 1 0 28060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_297
timestamp 1649977179
transform 1 0 28428 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1649977179
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_312
timestamp 1649977179
transform 1 0 29808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_319
timestamp 1649977179
transform 1 0 30452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_328
timestamp 1649977179
transform 1 0 31280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_341
timestamp 1649977179
transform 1 0 32476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_350
timestamp 1649977179
transform 1 0 33304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_354
timestamp 1649977179
transform 1 0 33672 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_381
timestamp 1649977179
transform 1 0 36156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_404
timestamp 1649977179
transform 1 0 38272 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_410
timestamp 1649977179
transform 1 0 38824 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_417
timestamp 1649977179
transform 1 0 39468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_431
timestamp 1649977179
transform 1 0 40756 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_437
timestamp 1649977179
transform 1 0 41308 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_443
timestamp 1649977179
transform 1 0 41860 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_463
timestamp 1649977179
transform 1 0 43700 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_473
timestamp 1649977179
transform 1 0 44620 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_483
timestamp 1649977179
transform 1 0 45540 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_502
timestamp 1649977179
transform 1 0 47288 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_515
timestamp 1649977179
transform 1 0 48484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_526
timestamp 1649977179
transform 1 0 49496 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_539
timestamp 1649977179
transform 1 0 50692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_554
timestamp 1649977179
transform 1 0 52072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_567
timestamp 1649977179
transform 1 0 53268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_574
timestamp 1649977179
transform 1 0 53912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_592
timestamp 1649977179
transform 1 0 55568 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_598
timestamp 1649977179
transform 1 0 56120 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_605
timestamp 1649977179
transform 1 0 56764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_618
timestamp 1649977179
transform 1 0 57960 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_631
timestamp 1649977179
transform 1 0 59156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_641
timestamp 1649977179
transform 1 0 60076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_653
timestamp 1649977179
transform 1 0 61180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_661
timestamp 1649977179
transform 1 0 61916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_680
timestamp 1649977179
transform 1 0 63664 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_687
timestamp 1649977179
transform 1 0 64308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1649977179
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1649977179
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_704
timestamp 1649977179
transform 1 0 65872 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_716
timestamp 1649977179
transform 1 0 66976 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_722
timestamp 1649977179
transform 1 0 67528 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_727
timestamp 1649977179
transform 1 0 67988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_734
timestamp 1649977179
transform 1 0 68632 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_744
timestamp 1649977179
transform 1 0 69552 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_753
timestamp 1649977179
transform 1 0 70380 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_773
timestamp 1649977179
transform 1 0 72220 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_785
timestamp 1649977179
transform 1 0 73324 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_797
timestamp 1649977179
transform 1 0 74428 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_809
timestamp 1649977179
transform 1 0 75532 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_813
timestamp 1649977179
transform 1 0 75900 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_825
timestamp 1649977179
transform 1 0 77004 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_837
timestamp 1649977179
transform 1 0 78108 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_849
timestamp 1649977179
transform 1 0 79212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_861
timestamp 1649977179
transform 1 0 80316 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_867
timestamp 1649977179
transform 1 0 80868 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_869
timestamp 1649977179
transform 1 0 81052 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_881
timestamp 1649977179
transform 1 0 82156 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_893
timestamp 1649977179
transform 1 0 83260 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_905
timestamp 1649977179
transform 1 0 84364 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_917
timestamp 1649977179
transform 1 0 85468 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_923
timestamp 1649977179
transform 1 0 86020 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_925
timestamp 1649977179
transform 1 0 86204 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_937
timestamp 1649977179
transform 1 0 87308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_948
timestamp 1649977179
transform 1 0 88320 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_6
timestamp 1649977179
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_18
timestamp 1649977179
transform 1 0 2760 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_22
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_34
timestamp 1649977179
transform 1 0 4232 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1649977179
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_191
timestamp 1649977179
transform 1 0 18676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_200
timestamp 1649977179
transform 1 0 19504 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_209
timestamp 1649977179
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_213
timestamp 1649977179
transform 1 0 20700 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_231
timestamp 1649977179
transform 1 0 22356 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_241
timestamp 1649977179
transform 1 0 23276 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1649977179
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_255
timestamp 1649977179
transform 1 0 24564 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_259
timestamp 1649977179
transform 1 0 24932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_267
timestamp 1649977179
transform 1 0 25668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1649977179
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_290
timestamp 1649977179
transform 1 0 27784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_299
timestamp 1649977179
transform 1 0 28612 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_308
timestamp 1649977179
transform 1 0 29440 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_320
timestamp 1649977179
transform 1 0 30544 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_326
timestamp 1649977179
transform 1 0 31096 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1649977179
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_344
timestamp 1649977179
transform 1 0 32752 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_348
timestamp 1649977179
transform 1 0 33120 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_355
timestamp 1649977179
transform 1 0 33764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_359
timestamp 1649977179
transform 1 0 34132 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_363
timestamp 1649977179
transform 1 0 34500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_367
timestamp 1649977179
transform 1 0 34868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_377
timestamp 1649977179
transform 1 0 35788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_381
timestamp 1649977179
transform 1 0 36156 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_389
timestamp 1649977179
transform 1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_401
timestamp 1649977179
transform 1 0 37996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_409
timestamp 1649977179
transform 1 0 38732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_420
timestamp 1649977179
transform 1 0 39744 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_426
timestamp 1649977179
transform 1 0 40296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_438
timestamp 1649977179
transform 1 0 41400 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1649977179
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_480
timestamp 1649977179
transform 1 0 45264 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_488
timestamp 1649977179
transform 1 0 46000 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_495
timestamp 1649977179
transform 1 0 46644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_501
timestamp 1649977179
transform 1 0 47196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_525
timestamp 1649977179
transform 1 0 49404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_545
timestamp 1649977179
transform 1 0 51244 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_579
timestamp 1649977179
transform 1 0 54372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_590
timestamp 1649977179
transform 1 0 55384 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_603
timestamp 1649977179
transform 1 0 56580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_607
timestamp 1649977179
transform 1 0 56948 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_613
timestamp 1649977179
transform 1 0 57500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_621
timestamp 1649977179
transform 1 0 58236 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_637
timestamp 1649977179
transform 1 0 59708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_655
timestamp 1649977179
transform 1 0 61364 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_666
timestamp 1649977179
transform 1 0 62376 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_679
timestamp 1649977179
transform 1 0 63572 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_688
timestamp 1649977179
transform 1 0 64400 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_696
timestamp 1649977179
transform 1 0 65136 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_708
timestamp 1649977179
transform 1 0 66240 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_720
timestamp 1649977179
transform 1 0 67344 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_725
timestamp 1649977179
transform 1 0 67804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_737
timestamp 1649977179
transform 1 0 68908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_741
timestamp 1649977179
transform 1 0 69276 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_758
timestamp 1649977179
transform 1 0 70840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_768
timestamp 1649977179
transform 1 0 71760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 1649977179
transform 1 0 72588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 1649977179
transform 1 0 73140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_785
timestamp 1649977179
transform 1 0 73324 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_792
timestamp 1649977179
transform 1 0 73968 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_804
timestamp 1649977179
transform 1 0 75072 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_816
timestamp 1649977179
transform 1 0 76176 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_828
timestamp 1649977179
transform 1 0 77280 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_841
timestamp 1649977179
transform 1 0 78476 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_853
timestamp 1649977179
transform 1 0 79580 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_865
timestamp 1649977179
transform 1 0 80684 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_877
timestamp 1649977179
transform 1 0 81788 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_889
timestamp 1649977179
transform 1 0 82892 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_895
timestamp 1649977179
transform 1 0 83444 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_897
timestamp 1649977179
transform 1 0 83628 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_909
timestamp 1649977179
transform 1 0 84732 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_921
timestamp 1649977179
transform 1 0 85836 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_933
timestamp 1649977179
transform 1 0 86940 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_948
timestamp 1649977179
transform 1 0 88320 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_6
timestamp 1649977179
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_214
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_224
timestamp 1649977179
transform 1 0 21712 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_235
timestamp 1649977179
transform 1 0 22724 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_260
timestamp 1649977179
transform 1 0 25024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_269
timestamp 1649977179
transform 1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_275
timestamp 1649977179
transform 1 0 26404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_295
timestamp 1649977179
transform 1 0 28244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1649977179
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_317
timestamp 1649977179
transform 1 0 30268 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_324
timestamp 1649977179
transform 1 0 30912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_352
timestamp 1649977179
transform 1 0 33488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_358
timestamp 1649977179
transform 1 0 34040 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1649977179
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_373
timestamp 1649977179
transform 1 0 35420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_381
timestamp 1649977179
transform 1 0 36156 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1649977179
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_394
timestamp 1649977179
transform 1 0 37352 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_409
timestamp 1649977179
transform 1 0 38732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_417
timestamp 1649977179
transform 1 0 39468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_437
timestamp 1649977179
transform 1 0 41308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_450
timestamp 1649977179
transform 1 0 42504 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_462
timestamp 1649977179
transform 1 0 43608 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_470
timestamp 1649977179
transform 1 0 44344 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_480
timestamp 1649977179
transform 1 0 45264 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_486
timestamp 1649977179
transform 1 0 45816 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_492
timestamp 1649977179
transform 1 0 46368 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_504
timestamp 1649977179
transform 1 0 47472 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_508
timestamp 1649977179
transform 1 0 47840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_516
timestamp 1649977179
transform 1 0 48576 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_529
timestamp 1649977179
transform 1 0 49772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_540
timestamp 1649977179
transform 1 0 50784 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_546
timestamp 1649977179
transform 1 0 51336 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_552
timestamp 1649977179
transform 1 0 51888 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_570
timestamp 1649977179
transform 1 0 53544 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_583
timestamp 1649977179
transform 1 0 54740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_608
timestamp 1649977179
transform 1 0 57040 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_615
timestamp 1649977179
transform 1 0 57684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_622
timestamp 1649977179
transform 1 0 58328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_641
timestamp 1649977179
transform 1 0 60076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_653
timestamp 1649977179
transform 1 0 61180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_662
timestamp 1649977179
transform 1 0 62008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_671
timestamp 1649977179
transform 1 0 62836 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_685
timestamp 1649977179
transform 1 0 64124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_695
timestamp 1649977179
transform 1 0 65044 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1649977179
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_701
timestamp 1649977179
transform 1 0 65596 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_709
timestamp 1649977179
transform 1 0 66332 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_726
timestamp 1649977179
transform 1 0 67896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_730
timestamp 1649977179
transform 1 0 68264 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_734
timestamp 1649977179
transform 1 0 68632 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_753
timestamp 1649977179
transform 1 0 70380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_766
timestamp 1649977179
transform 1 0 71576 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_774
timestamp 1649977179
transform 1 0 72312 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_786
timestamp 1649977179
transform 1 0 73416 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_798
timestamp 1649977179
transform 1 0 74520 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_810
timestamp 1649977179
transform 1 0 75624 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_813
timestamp 1649977179
transform 1 0 75900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_825
timestamp 1649977179
transform 1 0 77004 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_837
timestamp 1649977179
transform 1 0 78108 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_849
timestamp 1649977179
transform 1 0 79212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_861
timestamp 1649977179
transform 1 0 80316 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_867
timestamp 1649977179
transform 1 0 80868 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_869
timestamp 1649977179
transform 1 0 81052 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_881
timestamp 1649977179
transform 1 0 82156 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_893
timestamp 1649977179
transform 1 0 83260 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_905
timestamp 1649977179
transform 1 0 84364 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_917
timestamp 1649977179
transform 1 0 85468 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_923
timestamp 1649977179
transform 1 0 86020 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_925
timestamp 1649977179
transform 1 0 86204 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_937
timestamp 1649977179
transform 1 0 87308 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_943
timestamp 1649977179
transform 1 0 87860 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_948
timestamp 1649977179
transform 1 0 88320 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_196
timestamp 1649977179
transform 1 0 19136 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_204
timestamp 1649977179
transform 1 0 19872 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_212
timestamp 1649977179
transform 1 0 20608 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_232
timestamp 1649977179
transform 1 0 22448 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_241
timestamp 1649977179
transform 1 0 23276 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_255
timestamp 1649977179
transform 1 0 24564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_259
timestamp 1649977179
transform 1 0 24932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1649977179
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_290
timestamp 1649977179
transform 1 0 27784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_294
timestamp 1649977179
transform 1 0 28152 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_302
timestamp 1649977179
transform 1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_315
timestamp 1649977179
transform 1 0 30084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_321
timestamp 1649977179
transform 1 0 30636 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1649977179
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_346
timestamp 1649977179
transform 1 0 32936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_355
timestamp 1649977179
transform 1 0 33764 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_367
timestamp 1649977179
transform 1 0 34868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_375
timestamp 1649977179
transform 1 0 35604 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_409
timestamp 1649977179
transform 1 0 38732 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_415
timestamp 1649977179
transform 1 0 39284 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_432
timestamp 1649977179
transform 1 0 40848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_438
timestamp 1649977179
transform 1 0 41400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_445
timestamp 1649977179
transform 1 0 42044 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_453
timestamp 1649977179
transform 1 0 42780 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_466
timestamp 1649977179
transform 1 0 43976 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_475
timestamp 1649977179
transform 1 0 44804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_481
timestamp 1649977179
transform 1 0 45356 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_494
timestamp 1649977179
transform 1 0 46552 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_502
timestamp 1649977179
transform 1 0 47288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_509
timestamp 1649977179
transform 1 0 47932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1649977179
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_520
timestamp 1649977179
transform 1 0 48944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_524
timestamp 1649977179
transform 1 0 49312 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_548
timestamp 1649977179
transform 1 0 51520 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_556
timestamp 1649977179
transform 1 0 52256 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_571
timestamp 1649977179
transform 1 0 53636 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_577
timestamp 1649977179
transform 1 0 54188 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_583
timestamp 1649977179
transform 1 0 54740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_590
timestamp 1649977179
transform 1 0 55384 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_607
timestamp 1649977179
transform 1 0 56948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_613
timestamp 1649977179
transform 1 0 57500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_629
timestamp 1649977179
transform 1 0 58972 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_637
timestamp 1649977179
transform 1 0 59708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_655
timestamp 1649977179
transform 1 0 61364 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_661
timestamp 1649977179
transform 1 0 61916 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_669
timestamp 1649977179
transform 1 0 62652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_673
timestamp 1649977179
transform 1 0 63020 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_683
timestamp 1649977179
transform 1 0 63940 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_703
timestamp 1649977179
transform 1 0 65780 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_712
timestamp 1649977179
transform 1 0 66608 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1649977179
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1649977179
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_729
timestamp 1649977179
transform 1 0 68172 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_742
timestamp 1649977179
transform 1 0 69368 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_764
timestamp 1649977179
transform 1 0 71392 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_771
timestamp 1649977179
transform 1 0 72036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 1649977179
transform 1 0 73140 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_785
timestamp 1649977179
transform 1 0 73324 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_797
timestamp 1649977179
transform 1 0 74428 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_809
timestamp 1649977179
transform 1 0 75532 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_821
timestamp 1649977179
transform 1 0 76636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_833
timestamp 1649977179
transform 1 0 77740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_839
timestamp 1649977179
transform 1 0 78292 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_841
timestamp 1649977179
transform 1 0 78476 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_853
timestamp 1649977179
transform 1 0 79580 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_865
timestamp 1649977179
transform 1 0 80684 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_877
timestamp 1649977179
transform 1 0 81788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_889
timestamp 1649977179
transform 1 0 82892 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_895
timestamp 1649977179
transform 1 0 83444 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_897
timestamp 1649977179
transform 1 0 83628 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_909
timestamp 1649977179
transform 1 0 84732 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_921
timestamp 1649977179
transform 1 0 85836 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_933
timestamp 1649977179
transform 1 0 86940 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_945
timestamp 1649977179
transform 1 0 88044 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1649977179
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_215
timestamp 1649977179
transform 1 0 20884 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_227
timestamp 1649977179
transform 1 0 21988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_242
timestamp 1649977179
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1649977179
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_259
timestamp 1649977179
transform 1 0 24932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_263
timestamp 1649977179
transform 1 0 25300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_283
timestamp 1649977179
transform 1 0 27140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_295
timestamp 1649977179
transform 1 0 28244 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1649977179
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_319
timestamp 1649977179
transform 1 0 30452 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_341
timestamp 1649977179
transform 1 0 32476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1649977179
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_373
timestamp 1649977179
transform 1 0 35420 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_379
timestamp 1649977179
transform 1 0 35972 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_397
timestamp 1649977179
transform 1 0 37628 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_409
timestamp 1649977179
transform 1 0 38732 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_417
timestamp 1649977179
transform 1 0 39468 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_440
timestamp 1649977179
transform 1 0 41584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_449
timestamp 1649977179
transform 1 0 42412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_468
timestamp 1649977179
transform 1 0 44160 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_482
timestamp 1649977179
transform 1 0 45448 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_510
timestamp 1649977179
transform 1 0 48024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_519
timestamp 1649977179
transform 1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_526
timestamp 1649977179
transform 1 0 49496 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_537
timestamp 1649977179
transform 1 0 50508 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_546
timestamp 1649977179
transform 1 0 51336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_553
timestamp 1649977179
transform 1 0 51980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_566
timestamp 1649977179
transform 1 0 53176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_579
timestamp 1649977179
transform 1 0 54372 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_593
timestamp 1649977179
transform 1 0 55660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_606
timestamp 1649977179
transform 1 0 56856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_622
timestamp 1649977179
transform 1 0 58328 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_641
timestamp 1649977179
transform 1 0 60076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_645
timestamp 1649977179
transform 1 0 60444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_656
timestamp 1649977179
transform 1 0 61456 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_666
timestamp 1649977179
transform 1 0 62376 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_688
timestamp 1649977179
transform 1 0 64400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_694
timestamp 1649977179
transform 1 0 64952 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_707
timestamp 1649977179
transform 1 0 66148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_719
timestamp 1649977179
transform 1 0 67252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_728
timestamp 1649977179
transform 1 0 68080 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_734
timestamp 1649977179
transform 1 0 68632 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_753
timestamp 1649977179
transform 1 0 70380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_766
timestamp 1649977179
transform 1 0 71576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_772
timestamp 1649977179
transform 1 0 72128 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_778
timestamp 1649977179
transform 1 0 72680 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_790
timestamp 1649977179
transform 1 0 73784 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_802
timestamp 1649977179
transform 1 0 74888 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_810
timestamp 1649977179
transform 1 0 75624 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_813
timestamp 1649977179
transform 1 0 75900 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_825
timestamp 1649977179
transform 1 0 77004 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_837
timestamp 1649977179
transform 1 0 78108 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_849
timestamp 1649977179
transform 1 0 79212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_861
timestamp 1649977179
transform 1 0 80316 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_867
timestamp 1649977179
transform 1 0 80868 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_869
timestamp 1649977179
transform 1 0 81052 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_881
timestamp 1649977179
transform 1 0 82156 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_893
timestamp 1649977179
transform 1 0 83260 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_905
timestamp 1649977179
transform 1 0 84364 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_917
timestamp 1649977179
transform 1 0 85468 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_923
timestamp 1649977179
transform 1 0 86020 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_925
timestamp 1649977179
transform 1 0 86204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_937
timestamp 1649977179
transform 1 0 87308 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_943
timestamp 1649977179
transform 1 0 87860 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_948
timestamp 1649977179
transform 1 0 88320 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_19
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_23
timestamp 1649977179
transform 1 0 3220 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_35
timestamp 1649977179
transform 1 0 4324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1649977179
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_121
timestamp 1649977179
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_129
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_141
timestamp 1649977179
transform 1 0 14076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_153
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1649977179
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_231
timestamp 1649977179
transform 1 0 22356 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1649977179
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_247
timestamp 1649977179
transform 1 0 23828 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_257
timestamp 1649977179
transform 1 0 24748 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1649977179
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_298
timestamp 1649977179
transform 1 0 28520 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_306
timestamp 1649977179
transform 1 0 29256 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_314
timestamp 1649977179
transform 1 0 29992 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_320
timestamp 1649977179
transform 1 0 30544 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_327
timestamp 1649977179
transform 1 0 31188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1649977179
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_347
timestamp 1649977179
transform 1 0 33028 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_366
timestamp 1649977179
transform 1 0 34776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_372
timestamp 1649977179
transform 1 0 35328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1649977179
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_399
timestamp 1649977179
transform 1 0 37812 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_411
timestamp 1649977179
transform 1 0 38916 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_423
timestamp 1649977179
transform 1 0 40020 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_435
timestamp 1649977179
transform 1 0 41124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_442
timestamp 1649977179
transform 1 0 41768 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_459
timestamp 1649977179
transform 1 0 43332 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_470
timestamp 1649977179
transform 1 0 44344 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_479
timestamp 1649977179
transform 1 0 45172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_483
timestamp 1649977179
transform 1 0 45540 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_487
timestamp 1649977179
transform 1 0 45908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_499
timestamp 1649977179
transform 1 0 47012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_509
timestamp 1649977179
transform 1 0 47932 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_516
timestamp 1649977179
transform 1 0 48576 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_528
timestamp 1649977179
transform 1 0 49680 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_536
timestamp 1649977179
transform 1 0 50416 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_544
timestamp 1649977179
transform 1 0 51152 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_551
timestamp 1649977179
transform 1 0 51796 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_569
timestamp 1649977179
transform 1 0 53452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_583
timestamp 1649977179
transform 1 0 54740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_603
timestamp 1649977179
transform 1 0 56580 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_610
timestamp 1649977179
transform 1 0 57224 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_623
timestamp 1649977179
transform 1 0 58420 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_634
timestamp 1649977179
transform 1 0 59432 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_643
timestamp 1649977179
transform 1 0 60260 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_659
timestamp 1649977179
transform 1 0 61732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_666
timestamp 1649977179
transform 1 0 62376 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_678
timestamp 1649977179
transform 1 0 63480 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_684
timestamp 1649977179
transform 1 0 64032 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_688
timestamp 1649977179
transform 1 0 64400 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_696
timestamp 1649977179
transform 1 0 65136 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_705
timestamp 1649977179
transform 1 0 65964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_717
timestamp 1649977179
transform 1 0 67068 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_725
timestamp 1649977179
transform 1 0 67804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_729
timestamp 1649977179
transform 1 0 68172 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_735
timestamp 1649977179
transform 1 0 68724 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_739
timestamp 1649977179
transform 1 0 69092 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_744
timestamp 1649977179
transform 1 0 69552 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_763
timestamp 1649977179
transform 1 0 71300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_775
timestamp 1649977179
transform 1 0 72404 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 1649977179
transform 1 0 73140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_785
timestamp 1649977179
transform 1 0 73324 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_791
timestamp 1649977179
transform 1 0 73876 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_803
timestamp 1649977179
transform 1 0 74980 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_815
timestamp 1649977179
transform 1 0 76084 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_827
timestamp 1649977179
transform 1 0 77188 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_839
timestamp 1649977179
transform 1 0 78292 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_841
timestamp 1649977179
transform 1 0 78476 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_853
timestamp 1649977179
transform 1 0 79580 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_865
timestamp 1649977179
transform 1 0 80684 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_877
timestamp 1649977179
transform 1 0 81788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_889
timestamp 1649977179
transform 1 0 82892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_895
timestamp 1649977179
transform 1 0 83444 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_897
timestamp 1649977179
transform 1 0 83628 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_909
timestamp 1649977179
transform 1 0 84732 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_921
timestamp 1649977179
transform 1 0 85836 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_933
timestamp 1649977179
transform 1 0 86940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_948
timestamp 1649977179
transform 1 0 88320 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_6
timestamp 1649977179
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1649977179
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1649977179
transform 1 0 20608 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_216
timestamp 1649977179
transform 1 0 20976 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_224
timestamp 1649977179
transform 1 0 21712 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_236
timestamp 1649977179
transform 1 0 22816 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1649977179
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_268
timestamp 1649977179
transform 1 0 25760 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_288
timestamp 1649977179
transform 1 0 27600 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_294
timestamp 1649977179
transform 1 0 28152 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_300
timestamp 1649977179
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_324
timestamp 1649977179
transform 1 0 30912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_343
timestamp 1649977179
transform 1 0 32660 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_347
timestamp 1649977179
transform 1 0 33028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_371
timestamp 1649977179
transform 1 0 35236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_375
timestamp 1649977179
transform 1 0 35604 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_387
timestamp 1649977179
transform 1 0 36708 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_399
timestamp 1649977179
transform 1 0 37812 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_404
timestamp 1649977179
transform 1 0 38272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_410
timestamp 1649977179
transform 1 0 38824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1649977179
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_426
timestamp 1649977179
transform 1 0 40296 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_434
timestamp 1649977179
transform 1 0 41032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_440
timestamp 1649977179
transform 1 0 41584 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_459
timestamp 1649977179
transform 1 0 43332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_468
timestamp 1649977179
transform 1 0 44160 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_493
timestamp 1649977179
transform 1 0 46460 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_498
timestamp 1649977179
transform 1 0 46920 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_509
timestamp 1649977179
transform 1 0 47932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_521
timestamp 1649977179
transform 1 0 49036 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_529
timestamp 1649977179
transform 1 0 49772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_549
timestamp 1649977179
transform 1 0 51612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_565
timestamp 1649977179
transform 1 0 53084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_575
timestamp 1649977179
transform 1 0 54004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_584
timestamp 1649977179
transform 1 0 54832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_605
timestamp 1649977179
transform 1 0 56764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_611
timestamp 1649977179
transform 1 0 57316 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_615
timestamp 1649977179
transform 1 0 57684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_620
timestamp 1649977179
transform 1 0 58144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_627
timestamp 1649977179
transform 1 0 58788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_634
timestamp 1649977179
transform 1 0 59432 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_641
timestamp 1649977179
transform 1 0 60076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_649
timestamp 1649977179
transform 1 0 60812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_662
timestamp 1649977179
transform 1 0 62008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_671
timestamp 1649977179
transform 1 0 62836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_678
timestamp 1649977179
transform 1 0 63480 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_685
timestamp 1649977179
transform 1 0 64124 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_697
timestamp 1649977179
transform 1 0 65228 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_717
timestamp 1649977179
transform 1 0 67068 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_729
timestamp 1649977179
transform 1 0 68172 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_747
timestamp 1649977179
transform 1 0 69828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_753
timestamp 1649977179
transform 1 0 70380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_757
timestamp 1649977179
transform 1 0 70748 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_766
timestamp 1649977179
transform 1 0 71576 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_778
timestamp 1649977179
transform 1 0 72680 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_790
timestamp 1649977179
transform 1 0 73784 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_802
timestamp 1649977179
transform 1 0 74888 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_810
timestamp 1649977179
transform 1 0 75624 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_813
timestamp 1649977179
transform 1 0 75900 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_825
timestamp 1649977179
transform 1 0 77004 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_837
timestamp 1649977179
transform 1 0 78108 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_849
timestamp 1649977179
transform 1 0 79212 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_861
timestamp 1649977179
transform 1 0 80316 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_867
timestamp 1649977179
transform 1 0 80868 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_869
timestamp 1649977179
transform 1 0 81052 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_881
timestamp 1649977179
transform 1 0 82156 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_893
timestamp 1649977179
transform 1 0 83260 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_905
timestamp 1649977179
transform 1 0 84364 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_917
timestamp 1649977179
transform 1 0 85468 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_923
timestamp 1649977179
transform 1 0 86020 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_925
timestamp 1649977179
transform 1 0 86204 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_937
timestamp 1649977179
transform 1 0 87308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_948
timestamp 1649977179
transform 1 0 88320 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_10
timestamp 1649977179
transform 1 0 2024 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_22
timestamp 1649977179
transform 1 0 3128 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_34
timestamp 1649977179
transform 1 0 4232 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_46
timestamp 1649977179
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_242
timestamp 1649977179
transform 1 0 23368 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_253
timestamp 1649977179
transform 1 0 24380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_260
timestamp 1649977179
transform 1 0 25024 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_268
timestamp 1649977179
transform 1 0 25760 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1649977179
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_301
timestamp 1649977179
transform 1 0 28796 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_313
timestamp 1649977179
transform 1 0 29900 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_325
timestamp 1649977179
transform 1 0 31004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1649977179
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_346
timestamp 1649977179
transform 1 0 32936 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_350
timestamp 1649977179
transform 1 0 33304 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_357
timestamp 1649977179
transform 1 0 33948 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_369
timestamp 1649977179
transform 1 0 35052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1649977179
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_400
timestamp 1649977179
transform 1 0 37904 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_406
timestamp 1649977179
transform 1 0 38456 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_434
timestamp 1649977179
transform 1 0 41032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_438
timestamp 1649977179
transform 1 0 41400 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_445
timestamp 1649977179
transform 1 0 42044 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_458
timestamp 1649977179
transform 1 0 43240 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_465
timestamp 1649977179
transform 1 0 43884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_491
timestamp 1649977179
transform 1 0 46276 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1649977179
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_521
timestamp 1649977179
transform 1 0 49036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_525
timestamp 1649977179
transform 1 0 49404 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_532
timestamp 1649977179
transform 1 0 50048 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_536
timestamp 1649977179
transform 1 0 50416 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_543
timestamp 1649977179
transform 1 0 51060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_549
timestamp 1649977179
transform 1 0 51612 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_557
timestamp 1649977179
transform 1 0 52348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_566
timestamp 1649977179
transform 1 0 53176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_592
timestamp 1649977179
transform 1 0 55568 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_596
timestamp 1649977179
transform 1 0 55936 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_603
timestamp 1649977179
transform 1 0 56580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1649977179
transform 1 0 58236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_625
timestamp 1649977179
transform 1 0 58604 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_632
timestamp 1649977179
transform 1 0 59248 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_640
timestamp 1649977179
transform 1 0 59984 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_659
timestamp 1649977179
transform 1 0 61732 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_666
timestamp 1649977179
transform 1 0 62376 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_673
timestamp 1649977179
transform 1 0 63020 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_680
timestamp 1649977179
transform 1 0 63664 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_686
timestamp 1649977179
transform 1 0 64216 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_690
timestamp 1649977179
transform 1 0 64584 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_697
timestamp 1649977179
transform 1 0 65228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_701
timestamp 1649977179
transform 1 0 65596 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_712
timestamp 1649977179
transform 1 0 66608 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_718
timestamp 1649977179
transform 1 0 67160 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_726
timestamp 1649977179
transform 1 0 67896 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_729
timestamp 1649977179
transform 1 0 68172 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_738
timestamp 1649977179
transform 1 0 69000 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_744
timestamp 1649977179
transform 1 0 69552 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_764
timestamp 1649977179
transform 1 0 71392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_776
timestamp 1649977179
transform 1 0 72496 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_785
timestamp 1649977179
transform 1 0 73324 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_791
timestamp 1649977179
transform 1 0 73876 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_803
timestamp 1649977179
transform 1 0 74980 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_815
timestamp 1649977179
transform 1 0 76084 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_827
timestamp 1649977179
transform 1 0 77188 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_839
timestamp 1649977179
transform 1 0 78292 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_841
timestamp 1649977179
transform 1 0 78476 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_853
timestamp 1649977179
transform 1 0 79580 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_865
timestamp 1649977179
transform 1 0 80684 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_877
timestamp 1649977179
transform 1 0 81788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_889
timestamp 1649977179
transform 1 0 82892 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_895
timestamp 1649977179
transform 1 0 83444 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_897
timestamp 1649977179
transform 1 0 83628 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_909
timestamp 1649977179
transform 1 0 84732 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_921
timestamp 1649977179
transform 1 0 85836 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_933
timestamp 1649977179
transform 1 0 86940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_948
timestamp 1649977179
transform 1 0 88320 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_260
timestamp 1649977179
transform 1 0 25024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_282
timestamp 1649977179
transform 1 0 27048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1649977179
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_329
timestamp 1649977179
transform 1 0 31372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_341
timestamp 1649977179
transform 1 0 32476 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_349
timestamp 1649977179
transform 1 0 33212 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_382
timestamp 1649977179
transform 1 0 36248 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1649977179
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_425
timestamp 1649977179
transform 1 0 40204 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_435
timestamp 1649977179
transform 1 0 41124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_455
timestamp 1649977179
transform 1 0 42964 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_460
timestamp 1649977179
transform 1 0 43424 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 1649977179
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_481
timestamp 1649977179
transform 1 0 45356 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_488
timestamp 1649977179
transform 1 0 46000 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_496
timestamp 1649977179
transform 1 0 46736 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_506
timestamp 1649977179
transform 1 0 47656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_515
timestamp 1649977179
transform 1 0 48484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_524
timestamp 1649977179
transform 1 0 49312 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_539
timestamp 1649977179
transform 1 0 50692 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_551
timestamp 1649977179
transform 1 0 51796 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_563
timestamp 1649977179
transform 1 0 52900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_571
timestamp 1649977179
transform 1 0 53636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_580
timestamp 1649977179
transform 1 0 54464 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_594
timestamp 1649977179
transform 1 0 55752 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_602
timestamp 1649977179
transform 1 0 56488 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_608
timestamp 1649977179
transform 1 0 57040 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_620
timestamp 1649977179
transform 1 0 58144 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_633
timestamp 1649977179
transform 1 0 59340 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_637
timestamp 1649977179
transform 1 0 59708 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_641
timestamp 1649977179
transform 1 0 60076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_645
timestamp 1649977179
transform 1 0 60444 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_652
timestamp 1649977179
transform 1 0 61088 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_659
timestamp 1649977179
transform 1 0 61732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_663
timestamp 1649977179
transform 1 0 62100 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_670
timestamp 1649977179
transform 1 0 62744 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_682
timestamp 1649977179
transform 1 0 63848 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_697
timestamp 1649977179
transform 1 0 65228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_717
timestamp 1649977179
transform 1 0 67068 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_725
timestamp 1649977179
transform 1 0 67804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_729
timestamp 1649977179
transform 1 0 68172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_752
timestamp 1649977179
transform 1 0 70288 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_760
timestamp 1649977179
transform 1 0 71024 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_772
timestamp 1649977179
transform 1 0 72128 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_784
timestamp 1649977179
transform 1 0 73232 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_796
timestamp 1649977179
transform 1 0 74336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_808
timestamp 1649977179
transform 1 0 75440 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_813
timestamp 1649977179
transform 1 0 75900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_825
timestamp 1649977179
transform 1 0 77004 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_837
timestamp 1649977179
transform 1 0 78108 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_849
timestamp 1649977179
transform 1 0 79212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_861
timestamp 1649977179
transform 1 0 80316 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_867
timestamp 1649977179
transform 1 0 80868 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_869
timestamp 1649977179
transform 1 0 81052 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_881
timestamp 1649977179
transform 1 0 82156 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_893
timestamp 1649977179
transform 1 0 83260 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_905
timestamp 1649977179
transform 1 0 84364 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_917
timestamp 1649977179
transform 1 0 85468 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_923
timestamp 1649977179
transform 1 0 86020 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_925
timestamp 1649977179
transform 1 0 86204 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_937
timestamp 1649977179
transform 1 0 87308 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_949
timestamp 1649977179
transform 1 0 88412 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_6
timestamp 1649977179
transform 1 0 1656 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_18
timestamp 1649977179
transform 1 0 2760 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_30
timestamp 1649977179
transform 1 0 3864 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_42
timestamp 1649977179
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_245
timestamp 1649977179
transform 1 0 23644 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_260
timestamp 1649977179
transform 1 0 25024 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_266
timestamp 1649977179
transform 1 0 25576 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1649977179
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_285
timestamp 1649977179
transform 1 0 27324 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_289
timestamp 1649977179
transform 1 0 27692 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_301
timestamp 1649977179
transform 1 0 28796 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_307
timestamp 1649977179
transform 1 0 29348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_319
timestamp 1649977179
transform 1 0 30452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1649977179
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_354
timestamp 1649977179
transform 1 0 33672 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_366
timestamp 1649977179
transform 1 0 34776 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_372
timestamp 1649977179
transform 1 0 35328 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_376
timestamp 1649977179
transform 1 0 35696 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1649977179
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_444
timestamp 1649977179
transform 1 0 41952 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_478
timestamp 1649977179
transform 1 0 45080 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_490
timestamp 1649977179
transform 1 0 46184 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_502
timestamp 1649977179
transform 1 0 47288 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_511
timestamp 1649977179
transform 1 0 48116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_522
timestamp 1649977179
transform 1 0 49128 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_526
timestamp 1649977179
transform 1 0 49496 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_538
timestamp 1649977179
transform 1 0 50600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_550
timestamp 1649977179
transform 1 0 51704 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_558
timestamp 1649977179
transform 1 0 52440 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_582
timestamp 1649977179
transform 1 0 54648 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_591
timestamp 1649977179
transform 1 0 55476 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_600
timestamp 1649977179
transform 1 0 56304 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_612
timestamp 1649977179
transform 1 0 57408 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1649977179
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1649977179
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1649977179
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1649977179
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1649977179
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1649977179
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1649977179
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1649977179
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_709
timestamp 1649977179
transform 1 0 66332 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_715
timestamp 1649977179
transform 1 0 66884 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_725
timestamp 1649977179
transform 1 0 67804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_729
timestamp 1649977179
transform 1 0 68172 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_737
timestamp 1649977179
transform 1 0 68908 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_747
timestamp 1649977179
transform 1 0 69828 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_759
timestamp 1649977179
transform 1 0 70932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_771
timestamp 1649977179
transform 1 0 72036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 1649977179
transform 1 0 73140 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_785
timestamp 1649977179
transform 1 0 73324 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_797
timestamp 1649977179
transform 1 0 74428 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_809
timestamp 1649977179
transform 1 0 75532 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_821
timestamp 1649977179
transform 1 0 76636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_833
timestamp 1649977179
transform 1 0 77740 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_839
timestamp 1649977179
transform 1 0 78292 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_841
timestamp 1649977179
transform 1 0 78476 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_853
timestamp 1649977179
transform 1 0 79580 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_865
timestamp 1649977179
transform 1 0 80684 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_877
timestamp 1649977179
transform 1 0 81788 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_889
timestamp 1649977179
transform 1 0 82892 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_895
timestamp 1649977179
transform 1 0 83444 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_897
timestamp 1649977179
transform 1 0 83628 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_909
timestamp 1649977179
transform 1 0 84732 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_921
timestamp 1649977179
transform 1 0 85836 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_933
timestamp 1649977179
transform 1 0 86940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_945
timestamp 1649977179
transform 1 0 88044 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_6
timestamp 1649977179
transform 1 0 1656 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_10
timestamp 1649977179
transform 1 0 2024 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1649977179
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_261
timestamp 1649977179
transform 1 0 25116 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_273
timestamp 1649977179
transform 1 0 26220 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_285
timestamp 1649977179
transform 1 0 27324 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_297
timestamp 1649977179
transform 1 0 28428 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_305
timestamp 1649977179
transform 1 0 29164 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_382
timestamp 1649977179
transform 1 0 36248 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_394
timestamp 1649977179
transform 1 0 37352 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_406
timestamp 1649977179
transform 1 0 38456 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_418
timestamp 1649977179
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_508
timestamp 1649977179
transform 1 0 47840 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_520
timestamp 1649977179
transform 1 0 48944 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_610
timestamp 1649977179
transform 1 0 57224 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_622
timestamp 1649977179
transform 1 0 58328 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_634
timestamp 1649977179
transform 1 0 59432 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_642
timestamp 1649977179
transform 1 0 60168 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1649977179
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1649977179
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1649977179
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1649977179
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1649977179
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1649977179
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1649977179
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1649977179
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_725
timestamp 1649977179
transform 1 0 67804 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_737
timestamp 1649977179
transform 1 0 68908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 1649977179
transform 1 0 70012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 1649977179
transform 1 0 70564 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_757
timestamp 1649977179
transform 1 0 70748 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_769
timestamp 1649977179
transform 1 0 71852 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_781
timestamp 1649977179
transform 1 0 72956 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_793
timestamp 1649977179
transform 1 0 74060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 1649977179
transform 1 0 75164 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 1649977179
transform 1 0 75716 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_813
timestamp 1649977179
transform 1 0 75900 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_825
timestamp 1649977179
transform 1 0 77004 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_837
timestamp 1649977179
transform 1 0 78108 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_849
timestamp 1649977179
transform 1 0 79212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_861
timestamp 1649977179
transform 1 0 80316 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_867
timestamp 1649977179
transform 1 0 80868 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_869
timestamp 1649977179
transform 1 0 81052 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_881
timestamp 1649977179
transform 1 0 82156 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_893
timestamp 1649977179
transform 1 0 83260 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_905
timestamp 1649977179
transform 1 0 84364 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_917
timestamp 1649977179
transform 1 0 85468 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_923
timestamp 1649977179
transform 1 0 86020 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_925
timestamp 1649977179
transform 1 0 86204 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_937
timestamp 1649977179
transform 1 0 87308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_948
timestamp 1649977179
transform 1 0 88320 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_10
timestamp 1649977179
transform 1 0 2024 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_22
timestamp 1649977179
transform 1 0 3128 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_34
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_46
timestamp 1649977179
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1649977179
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1649977179
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_591
timestamp 1649977179
transform 1 0 55476 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_594
timestamp 1649977179
transform 1 0 55752 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_598
timestamp 1649977179
transform 1 0 56120 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_606
timestamp 1649977179
transform 1 0 56856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_610
timestamp 1649977179
transform 1 0 57224 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1649977179
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1649977179
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1649977179
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1649977179
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1649977179
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1649977179
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1649977179
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1649977179
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1649977179
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1649977179
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1649977179
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_729
timestamp 1649977179
transform 1 0 68172 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_741
timestamp 1649977179
transform 1 0 69276 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_753
timestamp 1649977179
transform 1 0 70380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_765
timestamp 1649977179
transform 1 0 71484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 1649977179
transform 1 0 72588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 1649977179
transform 1 0 73140 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_785
timestamp 1649977179
transform 1 0 73324 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_797
timestamp 1649977179
transform 1 0 74428 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_809
timestamp 1649977179
transform 1 0 75532 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_821
timestamp 1649977179
transform 1 0 76636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_833
timestamp 1649977179
transform 1 0 77740 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_839
timestamp 1649977179
transform 1 0 78292 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_841
timestamp 1649977179
transform 1 0 78476 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_853
timestamp 1649977179
transform 1 0 79580 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_865
timestamp 1649977179
transform 1 0 80684 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_877
timestamp 1649977179
transform 1 0 81788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_889
timestamp 1649977179
transform 1 0 82892 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_895
timestamp 1649977179
transform 1 0 83444 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_897
timestamp 1649977179
transform 1 0 83628 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_909
timestamp 1649977179
transform 1 0 84732 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_921
timestamp 1649977179
transform 1 0 85836 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_933
timestamp 1649977179
transform 1 0 86940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_948
timestamp 1649977179
transform 1 0 88320 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1649977179
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1649977179
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1649977179
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1649977179
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1649977179
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1649977179
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1649977179
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1649977179
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1649977179
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1649977179
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1649977179
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1649977179
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_725
timestamp 1649977179
transform 1 0 67804 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_737
timestamp 1649977179
transform 1 0 68908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 1649977179
transform 1 0 70012 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 1649977179
transform 1 0 70564 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_757
timestamp 1649977179
transform 1 0 70748 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_769
timestamp 1649977179
transform 1 0 71852 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_781
timestamp 1649977179
transform 1 0 72956 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_793
timestamp 1649977179
transform 1 0 74060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 1649977179
transform 1 0 75164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 1649977179
transform 1 0 75716 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_813
timestamp 1649977179
transform 1 0 75900 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_825
timestamp 1649977179
transform 1 0 77004 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_837
timestamp 1649977179
transform 1 0 78108 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_849
timestamp 1649977179
transform 1 0 79212 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_861
timestamp 1649977179
transform 1 0 80316 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_867
timestamp 1649977179
transform 1 0 80868 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_869
timestamp 1649977179
transform 1 0 81052 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_881
timestamp 1649977179
transform 1 0 82156 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_893
timestamp 1649977179
transform 1 0 83260 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_905
timestamp 1649977179
transform 1 0 84364 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_917
timestamp 1649977179
transform 1 0 85468 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_923
timestamp 1649977179
transform 1 0 86020 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_925
timestamp 1649977179
transform 1 0 86204 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_937
timestamp 1649977179
transform 1 0 87308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_943
timestamp 1649977179
transform 1 0 87860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_948
timestamp 1649977179
transform 1 0 88320 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_235
timestamp 1649977179
transform 1 0 22724 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_247
timestamp 1649977179
transform 1 0 23828 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_259
timestamp 1649977179
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1649977179
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_311
timestamp 1649977179
transform 1 0 29716 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_319
timestamp 1649977179
transform 1 0 30452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_331
timestamp 1649977179
transform 1 0 31556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1649977179
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1649977179
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1649977179
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1649977179
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1649977179
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1649977179
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1649977179
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1649977179
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1649977179
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1649977179
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1649977179
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_729
timestamp 1649977179
transform 1 0 68172 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_741
timestamp 1649977179
transform 1 0 69276 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_753
timestamp 1649977179
transform 1 0 70380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_765
timestamp 1649977179
transform 1 0 71484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_777
timestamp 1649977179
transform 1 0 72588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_783
timestamp 1649977179
transform 1 0 73140 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_785
timestamp 1649977179
transform 1 0 73324 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_797
timestamp 1649977179
transform 1 0 74428 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_809
timestamp 1649977179
transform 1 0 75532 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_821
timestamp 1649977179
transform 1 0 76636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_833
timestamp 1649977179
transform 1 0 77740 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_839
timestamp 1649977179
transform 1 0 78292 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_841
timestamp 1649977179
transform 1 0 78476 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_853
timestamp 1649977179
transform 1 0 79580 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_865
timestamp 1649977179
transform 1 0 80684 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_877
timestamp 1649977179
transform 1 0 81788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_889
timestamp 1649977179
transform 1 0 82892 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_895
timestamp 1649977179
transform 1 0 83444 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_897
timestamp 1649977179
transform 1 0 83628 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_909
timestamp 1649977179
transform 1 0 84732 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_921
timestamp 1649977179
transform 1 0 85836 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_933
timestamp 1649977179
transform 1 0 86940 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_945
timestamp 1649977179
transform 1 0 88044 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_6
timestamp 1649977179
transform 1 0 1656 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_10
timestamp 1649977179
transform 1 0 2024 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1649977179
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1649977179
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1649977179
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1649977179
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1649977179
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1649977179
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1649977179
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1649977179
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1649977179
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1649977179
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1649977179
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1649977179
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_725
timestamp 1649977179
transform 1 0 67804 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_737
timestamp 1649977179
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 1649977179
transform 1 0 70012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 1649977179
transform 1 0 70564 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_757
timestamp 1649977179
transform 1 0 70748 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_769
timestamp 1649977179
transform 1 0 71852 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_781
timestamp 1649977179
transform 1 0 72956 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_793
timestamp 1649977179
transform 1 0 74060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 1649977179
transform 1 0 75164 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 1649977179
transform 1 0 75716 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_813
timestamp 1649977179
transform 1 0 75900 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_825
timestamp 1649977179
transform 1 0 77004 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_837
timestamp 1649977179
transform 1 0 78108 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_849
timestamp 1649977179
transform 1 0 79212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_861
timestamp 1649977179
transform 1 0 80316 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_867
timestamp 1649977179
transform 1 0 80868 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_869
timestamp 1649977179
transform 1 0 81052 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_881
timestamp 1649977179
transform 1 0 82156 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_893
timestamp 1649977179
transform 1 0 83260 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_905
timestamp 1649977179
transform 1 0 84364 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_917
timestamp 1649977179
transform 1 0 85468 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_923
timestamp 1649977179
transform 1 0 86020 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_925
timestamp 1649977179
transform 1 0 86204 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_937
timestamp 1649977179
transform 1 0 87308 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_948
timestamp 1649977179
transform 1 0 88320 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_7
timestamp 1649977179
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_19
timestamp 1649977179
transform 1 0 2852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_34
timestamp 1649977179
transform 1 0 4232 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1649977179
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1649977179
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1649977179
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1649977179
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1649977179
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1649977179
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1649977179
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1649977179
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1649977179
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1649977179
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1649977179
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1649977179
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1649977179
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_729
timestamp 1649977179
transform 1 0 68172 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_741
timestamp 1649977179
transform 1 0 69276 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_753
timestamp 1649977179
transform 1 0 70380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_765
timestamp 1649977179
transform 1 0 71484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 1649977179
transform 1 0 72588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 1649977179
transform 1 0 73140 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_785
timestamp 1649977179
transform 1 0 73324 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_797
timestamp 1649977179
transform 1 0 74428 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_809
timestamp 1649977179
transform 1 0 75532 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_821
timestamp 1649977179
transform 1 0 76636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_833
timestamp 1649977179
transform 1 0 77740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_839
timestamp 1649977179
transform 1 0 78292 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_841
timestamp 1649977179
transform 1 0 78476 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_853
timestamp 1649977179
transform 1 0 79580 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_865
timestamp 1649977179
transform 1 0 80684 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_877
timestamp 1649977179
transform 1 0 81788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_889
timestamp 1649977179
transform 1 0 82892 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_895
timestamp 1649977179
transform 1 0 83444 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_897
timestamp 1649977179
transform 1 0 83628 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_909
timestamp 1649977179
transform 1 0 84732 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_921
timestamp 1649977179
transform 1 0 85836 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_933
timestamp 1649977179
transform 1 0 86940 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_943
timestamp 1649977179
transform 1 0 87860 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_948
timestamp 1649977179
transform 1 0 88320 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_6
timestamp 1649977179
transform 1 0 1656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_18
timestamp 1649977179
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1649977179
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1649977179
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1649977179
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1649977179
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1649977179
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1649977179
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1649977179
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1649977179
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1649977179
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1649977179
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1649977179
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1649977179
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1649977179
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_725
timestamp 1649977179
transform 1 0 67804 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_737
timestamp 1649977179
transform 1 0 68908 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 1649977179
transform 1 0 70012 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 1649977179
transform 1 0 70564 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_757
timestamp 1649977179
transform 1 0 70748 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_769
timestamp 1649977179
transform 1 0 71852 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_781
timestamp 1649977179
transform 1 0 72956 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_793
timestamp 1649977179
transform 1 0 74060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 1649977179
transform 1 0 75164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 1649977179
transform 1 0 75716 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_813
timestamp 1649977179
transform 1 0 75900 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_825
timestamp 1649977179
transform 1 0 77004 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_837
timestamp 1649977179
transform 1 0 78108 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_849
timestamp 1649977179
transform 1 0 79212 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_861
timestamp 1649977179
transform 1 0 80316 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_867
timestamp 1649977179
transform 1 0 80868 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_869
timestamp 1649977179
transform 1 0 81052 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_881
timestamp 1649977179
transform 1 0 82156 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_893
timestamp 1649977179
transform 1 0 83260 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_905
timestamp 1649977179
transform 1 0 84364 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_917
timestamp 1649977179
transform 1 0 85468 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_923
timestamp 1649977179
transform 1 0 86020 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_925
timestamp 1649977179
transform 1 0 86204 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_937
timestamp 1649977179
transform 1 0 87308 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_943
timestamp 1649977179
transform 1 0 87860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_948
timestamp 1649977179
transform 1 0 88320 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_6
timestamp 1649977179
transform 1 0 1656 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_18
timestamp 1649977179
transform 1 0 2760 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_30
timestamp 1649977179
transform 1 0 3864 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_42
timestamp 1649977179
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1649977179
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1649977179
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1649977179
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1649977179
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1649977179
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1649977179
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1649977179
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1649977179
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1649977179
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1649977179
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1649977179
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1649977179
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_729
timestamp 1649977179
transform 1 0 68172 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_741
timestamp 1649977179
transform 1 0 69276 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_753
timestamp 1649977179
transform 1 0 70380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_765
timestamp 1649977179
transform 1 0 71484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 1649977179
transform 1 0 72588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 1649977179
transform 1 0 73140 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_788
timestamp 1649977179
transform 1 0 73600 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_800
timestamp 1649977179
transform 1 0 74704 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_812
timestamp 1649977179
transform 1 0 75808 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_824
timestamp 1649977179
transform 1 0 76912 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_836
timestamp 1649977179
transform 1 0 78016 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_841
timestamp 1649977179
transform 1 0 78476 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_853
timestamp 1649977179
transform 1 0 79580 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_865
timestamp 1649977179
transform 1 0 80684 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_877
timestamp 1649977179
transform 1 0 81788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_889
timestamp 1649977179
transform 1 0 82892 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_895
timestamp 1649977179
transform 1 0 83444 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_897
timestamp 1649977179
transform 1 0 83628 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_909
timestamp 1649977179
transform 1 0 84732 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_921
timestamp 1649977179
transform 1 0 85836 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_933
timestamp 1649977179
transform 1 0 86940 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_941
timestamp 1649977179
transform 1 0 87676 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_948
timestamp 1649977179
transform 1 0 88320 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1649977179
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1649977179
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1649977179
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1649977179
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1649977179
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1649977179
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1649977179
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1649977179
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1649977179
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1649977179
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1649977179
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_725
timestamp 1649977179
transform 1 0 67804 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_737
timestamp 1649977179
transform 1 0 68908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 1649977179
transform 1 0 70012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 1649977179
transform 1 0 70564 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_757
timestamp 1649977179
transform 1 0 70748 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_769
timestamp 1649977179
transform 1 0 71852 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_781
timestamp 1649977179
transform 1 0 72956 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_793
timestamp 1649977179
transform 1 0 74060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 1649977179
transform 1 0 75164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 1649977179
transform 1 0 75716 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_813
timestamp 1649977179
transform 1 0 75900 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_825
timestamp 1649977179
transform 1 0 77004 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_837
timestamp 1649977179
transform 1 0 78108 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_849
timestamp 1649977179
transform 1 0 79212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_861
timestamp 1649977179
transform 1 0 80316 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_867
timestamp 1649977179
transform 1 0 80868 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_869
timestamp 1649977179
transform 1 0 81052 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_881
timestamp 1649977179
transform 1 0 82156 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_893
timestamp 1649977179
transform 1 0 83260 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_905
timestamp 1649977179
transform 1 0 84364 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_917
timestamp 1649977179
transform 1 0 85468 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_923
timestamp 1649977179
transform 1 0 86020 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_925
timestamp 1649977179
transform 1 0 86204 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_937
timestamp 1649977179
transform 1 0 87308 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_949
timestamp 1649977179
transform 1 0 88412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_10
timestamp 1649977179
transform 1 0 2024 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_22
timestamp 1649977179
transform 1 0 3128 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_34
timestamp 1649977179
transform 1 0 4232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_46
timestamp 1649977179
transform 1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1649977179
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_228
timestamp 1649977179
transform 1 0 22080 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_240
timestamp 1649977179
transform 1 0 23184 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_252
timestamp 1649977179
transform 1 0 24288 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_264
timestamp 1649977179
transform 1 0 25392 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1649977179
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1649977179
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1649977179
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1649977179
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1649977179
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1649977179
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1649977179
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1649977179
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1649977179
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1649977179
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1649977179
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1649977179
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_729
timestamp 1649977179
transform 1 0 68172 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_741
timestamp 1649977179
transform 1 0 69276 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_753
timestamp 1649977179
transform 1 0 70380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_765
timestamp 1649977179
transform 1 0 71484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 1649977179
transform 1 0 72588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 1649977179
transform 1 0 73140 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_785
timestamp 1649977179
transform 1 0 73324 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_797
timestamp 1649977179
transform 1 0 74428 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_809
timestamp 1649977179
transform 1 0 75532 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_821
timestamp 1649977179
transform 1 0 76636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_833
timestamp 1649977179
transform 1 0 77740 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_839
timestamp 1649977179
transform 1 0 78292 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_841
timestamp 1649977179
transform 1 0 78476 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_853
timestamp 1649977179
transform 1 0 79580 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_865
timestamp 1649977179
transform 1 0 80684 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_877
timestamp 1649977179
transform 1 0 81788 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_889
timestamp 1649977179
transform 1 0 82892 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_895
timestamp 1649977179
transform 1 0 83444 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_897
timestamp 1649977179
transform 1 0 83628 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_909
timestamp 1649977179
transform 1 0 84732 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_921
timestamp 1649977179
transform 1 0 85836 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_929
timestamp 1649977179
transform 1 0 86572 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_934
timestamp 1649977179
transform 1 0 87032 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_942
timestamp 1649977179
transform 1 0 87768 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_948
timestamp 1649977179
transform 1 0 88320 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1649977179
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1649977179
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1649977179
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1649977179
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1649977179
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1649977179
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1649977179
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1649977179
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1649977179
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1649977179
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1649977179
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_725
timestamp 1649977179
transform 1 0 67804 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_737
timestamp 1649977179
transform 1 0 68908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 1649977179
transform 1 0 70012 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 1649977179
transform 1 0 70564 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_757
timestamp 1649977179
transform 1 0 70748 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_769
timestamp 1649977179
transform 1 0 71852 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_781
timestamp 1649977179
transform 1 0 72956 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_793
timestamp 1649977179
transform 1 0 74060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 1649977179
transform 1 0 75164 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 1649977179
transform 1 0 75716 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_813
timestamp 1649977179
transform 1 0 75900 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_825
timestamp 1649977179
transform 1 0 77004 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_837
timestamp 1649977179
transform 1 0 78108 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_849
timestamp 1649977179
transform 1 0 79212 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_861
timestamp 1649977179
transform 1 0 80316 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_867
timestamp 1649977179
transform 1 0 80868 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_869
timestamp 1649977179
transform 1 0 81052 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_881
timestamp 1649977179
transform 1 0 82156 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_893
timestamp 1649977179
transform 1 0 83260 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_905
timestamp 1649977179
transform 1 0 84364 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_917
timestamp 1649977179
transform 1 0 85468 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_923
timestamp 1649977179
transform 1 0 86020 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_925
timestamp 1649977179
transform 1 0 86204 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_937
timestamp 1649977179
transform 1 0 87308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_948
timestamp 1649977179
transform 1 0 88320 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_13
timestamp 1649977179
transform 1 0 2300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_25
timestamp 1649977179
transform 1 0 3404 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_37
timestamp 1649977179
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1649977179
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1649977179
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1649977179
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1649977179
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1649977179
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1649977179
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1649977179
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1649977179
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1649977179
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1649977179
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1649977179
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1649977179
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_729
timestamp 1649977179
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_741
timestamp 1649977179
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_753
timestamp 1649977179
transform 1 0 70380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_765
timestamp 1649977179
transform 1 0 71484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 1649977179
transform 1 0 72588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 1649977179
transform 1 0 73140 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_785
timestamp 1649977179
transform 1 0 73324 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_797
timestamp 1649977179
transform 1 0 74428 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_809
timestamp 1649977179
transform 1 0 75532 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_821
timestamp 1649977179
transform 1 0 76636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_833
timestamp 1649977179
transform 1 0 77740 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_839
timestamp 1649977179
transform 1 0 78292 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_841
timestamp 1649977179
transform 1 0 78476 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_853
timestamp 1649977179
transform 1 0 79580 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_865
timestamp 1649977179
transform 1 0 80684 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_877
timestamp 1649977179
transform 1 0 81788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_889
timestamp 1649977179
transform 1 0 82892 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_895
timestamp 1649977179
transform 1 0 83444 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_897
timestamp 1649977179
transform 1 0 83628 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_909
timestamp 1649977179
transform 1 0 84732 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_921
timestamp 1649977179
transform 1 0 85836 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_933
timestamp 1649977179
transform 1 0 86940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_948
timestamp 1649977179
transform 1 0 88320 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_13
timestamp 1649977179
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1649977179
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1649977179
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1649977179
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1649977179
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1649977179
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1649977179
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1649977179
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1649977179
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1649977179
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1649977179
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1649977179
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1649977179
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_725
timestamp 1649977179
transform 1 0 67804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_737
timestamp 1649977179
transform 1 0 68908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 1649977179
transform 1 0 70012 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 1649977179
transform 1 0 70564 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_757
timestamp 1649977179
transform 1 0 70748 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_769
timestamp 1649977179
transform 1 0 71852 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_781
timestamp 1649977179
transform 1 0 72956 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_793
timestamp 1649977179
transform 1 0 74060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 1649977179
transform 1 0 75164 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 1649977179
transform 1 0 75716 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_813
timestamp 1649977179
transform 1 0 75900 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_825
timestamp 1649977179
transform 1 0 77004 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_837
timestamp 1649977179
transform 1 0 78108 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_849
timestamp 1649977179
transform 1 0 79212 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_861
timestamp 1649977179
transform 1 0 80316 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_867
timestamp 1649977179
transform 1 0 80868 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_869
timestamp 1649977179
transform 1 0 81052 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_881
timestamp 1649977179
transform 1 0 82156 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_893
timestamp 1649977179
transform 1 0 83260 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_905
timestamp 1649977179
transform 1 0 84364 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_917
timestamp 1649977179
transform 1 0 85468 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_923
timestamp 1649977179
transform 1 0 86020 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_925
timestamp 1649977179
transform 1 0 86204 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_937
timestamp 1649977179
transform 1 0 87308 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_941
timestamp 1649977179
transform 1 0 87676 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_948
timestamp 1649977179
transform 1 0 88320 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_6
timestamp 1649977179
transform 1 0 1656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_10
timestamp 1649977179
transform 1 0 2024 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_13
timestamp 1649977179
transform 1 0 2300 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_21
timestamp 1649977179
transform 1 0 3036 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_33
timestamp 1649977179
transform 1 0 4140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_45
timestamp 1649977179
transform 1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1649977179
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_288
timestamp 1649977179
transform 1 0 27600 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_292
timestamp 1649977179
transform 1 0 27968 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_304
timestamp 1649977179
transform 1 0 29072 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_316
timestamp 1649977179
transform 1 0 30176 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_328
timestamp 1649977179
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_467
timestamp 1649977179
transform 1 0 44068 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_479
timestamp 1649977179
transform 1 0 45172 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_491
timestamp 1649977179
transform 1 0 46276 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1649977179
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1649977179
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1649977179
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1649977179
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1649977179
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1649977179
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1649977179
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1649977179
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1649977179
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1649977179
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1649977179
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_729
timestamp 1649977179
transform 1 0 68172 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_741
timestamp 1649977179
transform 1 0 69276 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_753
timestamp 1649977179
transform 1 0 70380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_765
timestamp 1649977179
transform 1 0 71484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 1649977179
transform 1 0 72588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 1649977179
transform 1 0 73140 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_785
timestamp 1649977179
transform 1 0 73324 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_797
timestamp 1649977179
transform 1 0 74428 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_809
timestamp 1649977179
transform 1 0 75532 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_821
timestamp 1649977179
transform 1 0 76636 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_833
timestamp 1649977179
transform 1 0 77740 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_839
timestamp 1649977179
transform 1 0 78292 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_841
timestamp 1649977179
transform 1 0 78476 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_853
timestamp 1649977179
transform 1 0 79580 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_865
timestamp 1649977179
transform 1 0 80684 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_877
timestamp 1649977179
transform 1 0 81788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_889
timestamp 1649977179
transform 1 0 82892 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_895
timestamp 1649977179
transform 1 0 83444 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_897
timestamp 1649977179
transform 1 0 83628 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_909
timestamp 1649977179
transform 1 0 84732 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_921
timestamp 1649977179
transform 1 0 85836 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_929
timestamp 1649977179
transform 1 0 86572 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_933
timestamp 1649977179
transform 1 0 86940 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_937
timestamp 1649977179
transform 1 0 87308 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_942
timestamp 1649977179
transform 1 0 87768 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_948
timestamp 1649977179
transform 1 0 88320 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_13
timestamp 1649977179
transform 1 0 2300 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_22
timestamp 1649977179
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_32
timestamp 1649977179
transform 1 0 4048 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_44
timestamp 1649977179
transform 1 0 5152 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_56
timestamp 1649977179
transform 1 0 6256 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_68
timestamp 1649977179
transform 1 0 7360 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1649977179
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_281
timestamp 1649977179
transform 1 0 26956 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_287
timestamp 1649977179
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1649977179
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_314
timestamp 1649977179
transform 1 0 29992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_318
timestamp 1649977179
transform 1 0 30360 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_322
timestamp 1649977179
transform 1 0 30728 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_335
timestamp 1649977179
transform 1 0 31924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_347
timestamp 1649977179
transform 1 0 33028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1649977179
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_434
timestamp 1649977179
transform 1 0 41032 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_446
timestamp 1649977179
transform 1 0 42136 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_458
timestamp 1649977179
transform 1 0 43240 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_470
timestamp 1649977179
transform 1 0 44344 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1649977179
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1649977179
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1649977179
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1649977179
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1649977179
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1649977179
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1649977179
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1649977179
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1649977179
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1649977179
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1649977179
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_725
timestamp 1649977179
transform 1 0 67804 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_737
timestamp 1649977179
transform 1 0 68908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 1649977179
transform 1 0 70012 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 1649977179
transform 1 0 70564 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_757
timestamp 1649977179
transform 1 0 70748 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_769
timestamp 1649977179
transform 1 0 71852 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_781
timestamp 1649977179
transform 1 0 72956 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_793
timestamp 1649977179
transform 1 0 74060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 1649977179
transform 1 0 75164 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 1649977179
transform 1 0 75716 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_813
timestamp 1649977179
transform 1 0 75900 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_825
timestamp 1649977179
transform 1 0 77004 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_837
timestamp 1649977179
transform 1 0 78108 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_849
timestamp 1649977179
transform 1 0 79212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_861
timestamp 1649977179
transform 1 0 80316 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_867
timestamp 1649977179
transform 1 0 80868 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_869
timestamp 1649977179
transform 1 0 81052 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_881
timestamp 1649977179
transform 1 0 82156 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_893
timestamp 1649977179
transform 1 0 83260 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_905
timestamp 1649977179
transform 1 0 84364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_917
timestamp 1649977179
transform 1 0 85468 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_923
timestamp 1649977179
transform 1 0 86020 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_925
timestamp 1649977179
transform 1 0 86204 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_931
timestamp 1649977179
transform 1 0 86756 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_935
timestamp 1649977179
transform 1 0 87124 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_941
timestamp 1649977179
transform 1 0 87676 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_948
timestamp 1649977179
transform 1 0 88320 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_10
timestamp 1649977179
transform 1 0 2024 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_14
timestamp 1649977179
transform 1 0 2392 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_19
timestamp 1649977179
transform 1 0 2852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_25
timestamp 1649977179
transform 1 0 3404 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_34
timestamp 1649977179
transform 1 0 4232 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_46
timestamp 1649977179
transform 1 0 5336 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1649977179
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_64
timestamp 1649977179
transform 1 0 6992 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_70
timestamp 1649977179
transform 1 0 7544 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_82
timestamp 1649977179
transform 1 0 8648 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_94
timestamp 1649977179
transform 1 0 9752 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_100
timestamp 1649977179
transform 1 0 10304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1649977179
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_121
timestamp 1649977179
transform 1 0 12236 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_126
timestamp 1649977179
transform 1 0 12696 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_134
timestamp 1649977179
transform 1 0 13432 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_139
timestamp 1649977179
transform 1 0 13892 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_145
timestamp 1649977179
transform 1 0 14444 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_174
timestamp 1649977179
transform 1 0 17112 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_186
timestamp 1649977179
transform 1 0 18216 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_198
timestamp 1649977179
transform 1 0 19320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_201
timestamp 1649977179
transform 1 0 19596 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_206
timestamp 1649977179
transform 1 0 20056 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_212
timestamp 1649977179
transform 1 0 20608 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_245
timestamp 1649977179
transform 1 0 23644 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_251
timestamp 1649977179
transform 1 0 24196 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_263
timestamp 1649977179
transform 1 0 25300 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_271
timestamp 1649977179
transform 1 0 26036 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1649977179
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_285
timestamp 1649977179
transform 1 0 27324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_291
timestamp 1649977179
transform 1 0 27876 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_297
timestamp 1649977179
transform 1 0 28428 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_306
timestamp 1649977179
transform 1 0 29256 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_328
timestamp 1649977179
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_342
timestamp 1649977179
transform 1 0 32568 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_399
timestamp 1649977179
transform 1 0 37812 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_406
timestamp 1649977179
transform 1 0 38456 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_418
timestamp 1649977179
transform 1 0 39560 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_427
timestamp 1649977179
transform 1 0 40388 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_433
timestamp 1649977179
transform 1 0 40940 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_445
timestamp 1649977179
transform 1 0 42044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_455
timestamp 1649977179
transform 1 0 42964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_467
timestamp 1649977179
transform 1 0 44068 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_477
timestamp 1649977179
transform 1 0 44988 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_489
timestamp 1649977179
transform 1 0 46092 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_501
timestamp 1649977179
transform 1 0 47196 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_525
timestamp 1649977179
transform 1 0 49404 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_531
timestamp 1649977179
transform 1 0 49956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_543
timestamp 1649977179
transform 1 0 51060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_555
timestamp 1649977179
transform 1 0 52164 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_566
timestamp 1649977179
transform 1 0 53176 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_570
timestamp 1649977179
transform 1 0 53544 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_574
timestamp 1649977179
transform 1 0 53912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_587
timestamp 1649977179
transform 1 0 55108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_595
timestamp 1649977179
transform 1 0 55844 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_601
timestamp 1649977179
transform 1 0 56396 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_613
timestamp 1649977179
transform 1 0 57500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_624
timestamp 1649977179
transform 1 0 58512 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_630
timestamp 1649977179
transform 1 0 59064 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_642
timestamp 1649977179
transform 1 0 60168 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_646
timestamp 1649977179
transform 1 0 60536 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_650
timestamp 1649977179
transform 1 0 60904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_662
timestamp 1649977179
transform 1 0 62008 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_670
timestamp 1649977179
transform 1 0 62744 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1649977179
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_685
timestamp 1649977179
transform 1 0 64124 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_690
timestamp 1649977179
transform 1 0 64584 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_696
timestamp 1649977179
transform 1 0 65136 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_702
timestamp 1649977179
transform 1 0 65688 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_714
timestamp 1649977179
transform 1 0 66792 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_726
timestamp 1649977179
transform 1 0 67896 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_729
timestamp 1649977179
transform 1 0 68172 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_735
timestamp 1649977179
transform 1 0 68724 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_739
timestamp 1649977179
transform 1 0 69092 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_747
timestamp 1649977179
transform 1 0 69828 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_753
timestamp 1649977179
transform 1 0 70380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_765
timestamp 1649977179
transform 1 0 71484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 1649977179
transform 1 0 72588 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 1649977179
transform 1 0 73140 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_788
timestamp 1649977179
transform 1 0 73600 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_796
timestamp 1649977179
transform 1 0 74336 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_802
timestamp 1649977179
transform 1 0 74888 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_806
timestamp 1649977179
transform 1 0 75256 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_811
timestamp 1649977179
transform 1 0 75716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_823
timestamp 1649977179
transform 1 0 76820 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_832
timestamp 1649977179
transform 1 0 77648 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_841
timestamp 1649977179
transform 1 0 78476 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_853
timestamp 1649977179
transform 1 0 79580 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_857
timestamp 1649977179
transform 1 0 79948 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_869
timestamp 1649977179
transform 1 0 81052 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_881
timestamp 1649977179
transform 1 0 82156 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_893
timestamp 1649977179
transform 1 0 83260 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_897
timestamp 1649977179
transform 1 0 83628 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_905
timestamp 1649977179
transform 1 0 84364 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_909
timestamp 1649977179
transform 1 0 84732 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_913
timestamp 1649977179
transform 1 0 85100 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_918
timestamp 1649977179
transform 1 0 85560 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_929
timestamp 1649977179
transform 1 0 86572 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_935
timestamp 1649977179
transform 1 0 87124 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_948
timestamp 1649977179
transform 1 0 88320 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_7
timestamp 1649977179
transform 1 0 1748 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1649977179
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1649977179
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_33
timestamp 1649977179
transform 1 0 4140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_37
timestamp 1649977179
transform 1 0 4508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_42
timestamp 1649977179
transform 1 0 4968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_48
timestamp 1649977179
transform 1 0 5520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_67
timestamp 1649977179
transform 1 0 7268 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_71
timestamp 1649977179
transform 1 0 7636 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_75
timestamp 1649977179
transform 1 0 8004 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1649977179
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_90
timestamp 1649977179
transform 1 0 9384 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_94
timestamp 1649977179
transform 1 0 9752 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_98
timestamp 1649977179
transform 1 0 10120 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_113
timestamp 1649977179
transform 1 0 11500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_124
timestamp 1649977179
transform 1 0 12512 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1649977179
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_146
timestamp 1649977179
transform 1 0 14536 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_160
timestamp 1649977179
transform 1 0 15824 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_179
timestamp 1649977179
transform 1 0 17572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_183
timestamp 1649977179
transform 1 0 17940 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_187
timestamp 1649977179
transform 1 0 18308 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1649977179
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_202
timestamp 1649977179
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_215
timestamp 1649977179
transform 1 0 20884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_225
timestamp 1649977179
transform 1 0 21804 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_230
timestamp 1649977179
transform 1 0 22264 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_236
timestamp 1649977179
transform 1 0 22816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1649977179
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1649977179
transform 1 0 24840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_262
timestamp 1649977179
transform 1 0 25208 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_266
timestamp 1649977179
transform 1 0 25576 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_273
timestamp 1649977179
transform 1 0 26220 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_279
timestamp 1649977179
transform 1 0 26772 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_281
timestamp 1649977179
transform 1 0 26956 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_286
timestamp 1649977179
transform 1 0 27416 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_293
timestamp 1649977179
transform 1 0 28060 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_299
timestamp 1649977179
transform 1 0 28612 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_305
timestamp 1649977179
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_314
timestamp 1649977179
transform 1 0 29992 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_322
timestamp 1649977179
transform 1 0 30728 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_347
timestamp 1649977179
transform 1 0 33028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_351
timestamp 1649977179
transform 1 0 33396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_355
timestamp 1649977179
transform 1 0 33764 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1649977179
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_370
timestamp 1649977179
transform 1 0 35144 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_383
timestamp 1649977179
transform 1 0 36340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_393
timestamp 1649977179
transform 1 0 37260 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_398
timestamp 1649977179
transform 1 0 37720 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_405
timestamp 1649977179
transform 1 0 38364 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_412
timestamp 1649977179
transform 1 0 39008 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_424
timestamp 1649977179
transform 1 0 40112 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_439
timestamp 1649977179
transform 1 0 41492 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_449
timestamp 1649977179
transform 1 0 42412 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_454
timestamp 1649977179
transform 1 0 42872 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_461
timestamp 1649977179
transform 1 0 43516 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_467
timestamp 1649977179
transform 1 0 44068 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_473
timestamp 1649977179
transform 1 0 44620 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_482
timestamp 1649977179
transform 1 0 45448 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_496
timestamp 1649977179
transform 1 0 46736 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_505
timestamp 1649977179
transform 1 0 47564 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_517
timestamp 1649977179
transform 1 0 48668 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_524
timestamp 1649977179
transform 1 0 49312 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_540
timestamp 1649977179
transform 1 0 50784 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_546
timestamp 1649977179
transform 1 0 51336 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_552
timestamp 1649977179
transform 1 0 51888 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_564
timestamp 1649977179
transform 1 0 52992 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_580
timestamp 1649977179
transform 1 0 54464 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_597
timestamp 1649977179
transform 1 0 56028 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_608
timestamp 1649977179
transform 1 0 57040 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_620
timestamp 1649977179
transform 1 0 58144 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_630
timestamp 1649977179
transform 1 0 59064 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_636
timestamp 1649977179
transform 1 0 59616 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_648
timestamp 1649977179
transform 1 0 60720 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_658
timestamp 1649977179
transform 1 0 61640 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_664
timestamp 1649977179
transform 1 0 62192 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_676
timestamp 1649977179
transform 1 0 63296 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_692
timestamp 1649977179
transform 1 0 64768 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_704
timestamp 1649977179
transform 1 0 65872 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_710
timestamp 1649977179
transform 1 0 66424 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_716
timestamp 1649977179
transform 1 0 66976 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_722
timestamp 1649977179
transform 1 0 67528 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_729
timestamp 1649977179
transform 1 0 68172 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_736
timestamp 1649977179
transform 1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_742
timestamp 1649977179
transform 1 0 69368 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_748
timestamp 1649977179
transform 1 0 69920 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_760
timestamp 1649977179
transform 1 0 71024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_766
timestamp 1649977179
transform 1 0 71576 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_772
timestamp 1649977179
transform 1 0 72128 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_778
timestamp 1649977179
transform 1 0 72680 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_785
timestamp 1649977179
transform 1 0 73324 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_792
timestamp 1649977179
transform 1 0 73968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_798
timestamp 1649977179
transform 1 0 74520 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_804
timestamp 1649977179
transform 1 0 75072 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_813
timestamp 1649977179
transform 1 0 75900 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_820
timestamp 1649977179
transform 1 0 76544 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_826
timestamp 1649977179
transform 1 0 77096 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_832
timestamp 1649977179
transform 1 0 77648 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_841
timestamp 1649977179
transform 1 0 78476 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_848
timestamp 1649977179
transform 1 0 79120 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_855
timestamp 1649977179
transform 1 0 79764 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_862
timestamp 1649977179
transform 1 0 80408 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_869
timestamp 1649977179
transform 1 0 81052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_876
timestamp 1649977179
transform 1 0 81696 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_882
timestamp 1649977179
transform 1 0 82248 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_889
timestamp 1649977179
transform 1 0 82892 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_895
timestamp 1649977179
transform 1 0 83444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_900
timestamp 1649977179
transform 1 0 83904 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_906
timestamp 1649977179
transform 1 0 84456 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_912
timestamp 1649977179
transform 1 0 85008 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_917
timestamp 1649977179
transform 1 0 85468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_923
timestamp 1649977179
transform 1 0 86020 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_928
timestamp 1649977179
transform 1 0 86480 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_935
timestamp 1649977179
transform 1 0 87124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_948
timestamp 1649977179
transform 1 0 88320 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 88872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 88872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 88872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 88872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 88872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 88872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 88872 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 88872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 88872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 88872 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 88872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 88872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 88872 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 88872 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 88872 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 88872 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 88872 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 88872 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 88872 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 88872 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 88872 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 88872 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 88872 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 88872 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 88872 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 88872 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 88872 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 88872 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 88872 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 88872 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 88872 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 88872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 88872 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 88872 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 88872 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 88872 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 88872 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 88872 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 88872 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 88872 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 88872 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 88872 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 88872 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 88872 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 88872 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 88872 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 88872 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 80960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 86112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 83536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 80960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 86112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 83536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 80960 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 86112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 83536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 80960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 86112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 83536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 80960 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 86112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 83536 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 80960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 86112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 83536 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 80960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 86112 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 83536 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 70656 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 75808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 80960 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 86112 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 73232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 78384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 83536 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 70656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 75808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 80960 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 86112 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 73232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 78384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 83536 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 70656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 75808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 80960 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 86112 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 73232 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 78384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 83536 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 70656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 75808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 80960 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 86112 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 73232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 78384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 83536 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 70656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 75808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 80960 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 86112 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 73232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 78384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 83536 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 70656 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 75808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 80960 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 86112 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 73232 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 78384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 83536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 70656 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 75808 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 80960 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 86112 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 73232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 78384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 83536 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 70656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 75808 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 80960 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 86112 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 73232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 78384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 83536 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 70656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 75808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 80960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 86112 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 73232 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 78384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 83536 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 32016 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 37168 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 42320 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 47472 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 52624 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 57776 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 62928 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 68080 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 70656 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 73232 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 75808 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 78384 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 80960 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 83536 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 86112 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0534_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 48024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0535_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 48208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0536_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0537_
timestamp 1649977179
transform 1 0 52808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0538_
timestamp 1649977179
transform 1 0 37904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0539_
timestamp 1649977179
transform 1 0 61088 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0540_
timestamp 1649977179
transform 1 0 60444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0541_
timestamp 1649977179
transform 1 0 37536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0542_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 49496 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0543_
timestamp 1649977179
transform 1 0 45448 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0544_
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0545_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0546_
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0547_
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0548_
timestamp 1649977179
transform 1 0 31556 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0549_
timestamp 1649977179
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0550_
timestamp 1649977179
transform 1 0 35880 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0551_
timestamp 1649977179
transform 1 0 48852 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0552_
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1649977179
transform 1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0554_
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0555_
timestamp 1649977179
transform 1 0 28520 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0556_
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0557_
timestamp 1649977179
transform 1 0 20056 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0558_
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0559_
timestamp 1649977179
transform 1 0 30084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0560_
timestamp 1649977179
transform 1 0 28244 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0561_
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0562_
timestamp 1649977179
transform 1 0 22172 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0563_
timestamp 1649977179
transform 1 0 29808 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0564_
timestamp 1649977179
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0565_
timestamp 1649977179
transform 1 0 21896 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0566_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0567_
timestamp 1649977179
transform 1 0 25852 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0568_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0569_
timestamp 1649977179
transform 1 0 38824 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0570_
timestamp 1649977179
transform 1 0 37904 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0571_
timestamp 1649977179
transform 1 0 39836 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0572_
timestamp 1649977179
transform 1 0 25944 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0573_
timestamp 1649977179
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0574_
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0575_
timestamp 1649977179
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0576_
timestamp 1649977179
transform 1 0 32476 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0577_
timestamp 1649977179
transform 1 0 20056 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0578_
timestamp 1649977179
transform 1 0 21160 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0579_
timestamp 1649977179
transform 1 0 32660 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0580_
timestamp 1649977179
transform 1 0 29900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0581_
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0582_
timestamp 1649977179
transform 1 0 30084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0583_
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0584_
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0585_
timestamp 1649977179
transform 1 0 18584 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0586_
timestamp 1649977179
transform 1 0 24932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0587_
timestamp 1649977179
transform 1 0 63112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0588_
timestamp 1649977179
transform 1 0 63572 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0589_
timestamp 1649977179
transform 1 0 46276 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0590_
timestamp 1649977179
transform 1 0 50416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0591_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0592_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38272 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0593_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37168 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0594_
timestamp 1649977179
transform 1 0 30728 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0595_
timestamp 1649977179
transform 1 0 59432 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0596_
timestamp 1649977179
transform 1 0 29624 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1649977179
transform 1 0 30360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0598_
timestamp 1649977179
transform 1 0 50324 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1649977179
transform 1 0 19228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0600_
timestamp 1649977179
transform 1 0 61548 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0601_
timestamp 1649977179
transform 1 0 63664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0602_
timestamp 1649977179
transform 1 0 43608 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0603_
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0604_
timestamp 1649977179
transform 1 0 40572 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0605_
timestamp 1649977179
transform 1 0 40664 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0606_
timestamp 1649977179
transform 1 0 33488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0607_
timestamp 1649977179
transform 1 0 27048 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1649977179
transform 1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0609_
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0610_
timestamp 1649977179
transform 1 0 31004 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0611_
timestamp 1649977179
transform 1 0 35604 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0612_
timestamp 1649977179
transform 1 0 39192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0613_
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1649977179
transform 1 0 14536 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0615_
timestamp 1649977179
transform 1 0 40020 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0616_
timestamp 1649977179
transform 1 0 40664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0617_
timestamp 1649977179
transform 1 0 29808 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0618_
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0619_
timestamp 1649977179
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0620_
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1649977179
transform 1 0 58236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0622_
timestamp 1649977179
transform 1 0 19688 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0623_
timestamp 1649977179
transform 1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0624_
timestamp 1649977179
transform 1 0 3772 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0625_
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0626_
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1649977179
transform 1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0628_
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0629_
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1649977179
transform 1 0 30452 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0631_
timestamp 1649977179
transform 1 0 77464 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0632_
timestamp 1649977179
transform 1 0 78476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0633_
timestamp 1649977179
transform 1 0 39284 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0634_
timestamp 1649977179
transform 1 0 41768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0635_
timestamp 1649977179
transform 1 0 77188 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1649977179
transform 1 0 79672 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0637_
timestamp 1649977179
transform 1 0 41400 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0638_
timestamp 1649977179
transform 1 0 41676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0639_
timestamp 1649977179
transform 1 0 28888 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0640_
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0641_
timestamp 1649977179
transform 1 0 26496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0642_
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1649977179
transform 1 0 55660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0644_
timestamp 1649977179
transform 1 0 71116 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1649977179
transform 1 0 71392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0646_
timestamp 1649977179
transform 1 0 28796 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0647_
timestamp 1649977179
transform 1 0 56120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0648_
timestamp 1649977179
transform 1 0 71116 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0649_
timestamp 1649977179
transform 1 0 73600 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0650_
timestamp 1649977179
transform 1 0 28520 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0651_
timestamp 1649977179
transform 1 0 26128 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1649977179
transform 1 0 27232 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0653_
timestamp 1649977179
transform 1 0 28244 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1649977179
transform 1 0 28980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0655_
timestamp 1649977179
transform 1 0 27416 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 1649977179
transform 1 0 28152 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0657_
timestamp 1649977179
transform 1 0 23552 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0658_
timestamp 1649977179
transform 1 0 17940 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0659_
timestamp 1649977179
transform 1 0 12512 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1649977179
transform 1 0 2944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0661_
timestamp 1649977179
transform 1 0 31188 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1649977179
transform 1 0 31464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0663_
timestamp 1649977179
transform 1 0 73508 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0664_
timestamp 1649977179
transform 1 0 74612 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0665_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 51152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0666_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 51060 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0667_
timestamp 1649977179
transform 1 0 55660 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0668_
timestamp 1649977179
transform 1 0 63940 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0669_
timestamp 1649977179
transform 1 0 41124 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0670_
timestamp 1649977179
transform 1 0 52624 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0671_
timestamp 1649977179
transform 1 0 54188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0672_
timestamp 1649977179
transform 1 0 46552 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1649977179
transform 1 0 41124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0674_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44528 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0675_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43884 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0676_
timestamp 1649977179
transform 1 0 58236 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0677_
timestamp 1649977179
transform 1 0 57224 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0678_
timestamp 1649977179
transform 1 0 49588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0679_
timestamp 1649977179
transform 1 0 49956 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0681_
timestamp 1649977179
transform 1 0 54556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0682_
timestamp 1649977179
transform 1 0 56672 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0683_
timestamp 1649977179
transform 1 0 57040 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0684_
timestamp 1649977179
transform 1 0 58328 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1649977179
transform 1 0 30360 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0686_
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _0687_
timestamp 1649977179
transform 1 0 54004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0688_
timestamp 1649977179
transform 1 0 59432 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0689_
timestamp 1649977179
transform 1 0 53360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0690_
timestamp 1649977179
transform 1 0 59616 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1649977179
transform 1 0 56672 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0692_
timestamp 1649977179
transform 1 0 55200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0693_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 58604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0694_
timestamp 1649977179
transform 1 0 53544 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1649977179
transform 1 0 48944 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0696_
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0697_
timestamp 1649977179
transform 1 0 52900 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0698_
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1649977179
transform 1 0 54648 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0700_
timestamp 1649977179
transform 1 0 53544 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0701_
timestamp 1649977179
transform 1 0 51428 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0702_
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0703_
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0704_
timestamp 1649977179
transform 1 0 53820 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0705_
timestamp 1649977179
transform 1 0 55016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1649977179
transform 1 0 49496 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0707_
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0708_
timestamp 1649977179
transform 1 0 51428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0709_
timestamp 1649977179
transform 1 0 60444 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0710_
timestamp 1649977179
transform 1 0 61916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1649977179
transform 1 0 62100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0712_
timestamp 1649977179
transform 1 0 48576 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0713_
timestamp 1649977179
transform 1 0 59708 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0714_
timestamp 1649977179
transform 1 0 64860 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0715_
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0716_
timestamp 1649977179
transform 1 0 62928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0717_
timestamp 1649977179
transform 1 0 63020 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0719_
timestamp 1649977179
transform 1 0 62284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0720_
timestamp 1649977179
transform 1 0 61640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0721_
timestamp 1649977179
transform 1 0 67160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1649977179
transform 1 0 68356 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0723_
timestamp 1649977179
transform 1 0 67620 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0724_
timestamp 1649977179
transform 1 0 66240 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0725_
timestamp 1649977179
transform 1 0 69828 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1649977179
transform 1 0 72312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0727_
timestamp 1649977179
transform 1 0 68264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0728_
timestamp 1649977179
transform 1 0 68908 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0729_
timestamp 1649977179
transform 1 0 59064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0730_
timestamp 1649977179
transform 1 0 72036 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0731_
timestamp 1649977179
transform 1 0 56672 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1649977179
transform 1 0 72404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0733_
timestamp 1649977179
transform 1 0 69184 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0734_
timestamp 1649977179
transform 1 0 68724 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0735_
timestamp 1649977179
transform 1 0 60444 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0736_
timestamp 1649977179
transform 1 0 61456 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1649977179
transform 1 0 35328 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0738_
timestamp 1649977179
transform 1 0 58052 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _0739_
timestamp 1649977179
transform 1 0 59064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0740_
timestamp 1649977179
transform 1 0 60444 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0741_
timestamp 1649977179
transform 1 0 60536 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0742_
timestamp 1649977179
transform 1 0 63388 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0744_
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0745_
timestamp 1649977179
transform 1 0 62008 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0746_
timestamp 1649977179
transform 1 0 66056 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1649977179
transform 1 0 55844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0748_
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0749_
timestamp 1649977179
transform 1 0 64400 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0750_
timestamp 1649977179
transform 1 0 65412 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1649977179
transform 1 0 41492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0752_
timestamp 1649977179
transform 1 0 58052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0753_
timestamp 1649977179
transform 1 0 64492 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0754_
timestamp 1649977179
transform 1 0 57960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0755_
timestamp 1649977179
transform 1 0 62284 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0756_
timestamp 1649977179
transform 1 0 57132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0758_
timestamp 1649977179
transform 1 0 57776 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0759_
timestamp 1649977179
transform 1 0 58696 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0760_
timestamp 1649977179
transform 1 0 57316 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0761_
timestamp 1649977179
transform 1 0 59708 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0763_
timestamp 1649977179
transform 1 0 56856 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0764_
timestamp 1649977179
transform 1 0 58420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0765_
timestamp 1649977179
transform 1 0 58696 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0766_
timestamp 1649977179
transform 1 0 51888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0767_
timestamp 1649977179
transform 1 0 51244 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1649977179
transform 1 0 56120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0769_
timestamp 1649977179
transform 1 0 55016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0770_
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0771_
timestamp 1649977179
transform 1 0 46552 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1649977179
transform 1 0 38180 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0773_
timestamp 1649977179
transform 1 0 46552 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0774_
timestamp 1649977179
transform 1 0 46920 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0775_
timestamp 1649977179
transform 1 0 47932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1649977179
transform 1 0 45080 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0777_
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0778_
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0779_
timestamp 1649977179
transform 1 0 49128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0780_
timestamp 1649977179
transform 1 0 43608 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0781_
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1649977179
transform 1 0 51336 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0783_
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0784_
timestamp 1649977179
transform 1 0 42596 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0785_
timestamp 1649977179
transform 1 0 55660 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0786_
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1649977179
transform 1 0 38548 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0788_
timestamp 1649977179
transform 1 0 52256 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _0789_
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0790_
timestamp 1649977179
transform 1 0 43608 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0791_
timestamp 1649977179
transform 1 0 51980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0792_
timestamp 1649977179
transform 1 0 53084 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0794_
timestamp 1649977179
transform 1 0 51612 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0795_
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0796_
timestamp 1649977179
transform 1 0 53912 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1649977179
transform 1 0 66884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0798_
timestamp 1649977179
transform 1 0 53268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0799_
timestamp 1649977179
transform 1 0 53452 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0800_
timestamp 1649977179
transform 1 0 47472 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1649977179
transform 1 0 68356 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0802_
timestamp 1649977179
transform 1 0 48208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0803_
timestamp 1649977179
transform 1 0 46276 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0804_
timestamp 1649977179
transform 1 0 54280 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0805_
timestamp 1649977179
transform 1 0 53544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1649977179
transform 1 0 68448 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0807_
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0808_
timestamp 1649977179
transform 1 0 53360 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0809_
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0810_
timestamp 1649977179
transform 1 0 42596 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0811_
timestamp 1649977179
transform 1 0 38916 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1649977179
transform 1 0 34040 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0813_
timestamp 1649977179
transform 1 0 41584 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _0814_
timestamp 1649977179
transform 1 0 35236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0815_
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0816_
timestamp 1649977179
transform 1 0 33672 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1649977179
transform 1 0 34592 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0818_
timestamp 1649977179
transform 1 0 33672 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0819_
timestamp 1649977179
transform 1 0 34500 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0820_
timestamp 1649977179
transform 1 0 36340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1649977179
transform 1 0 36432 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0822_
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0823_
timestamp 1649977179
transform 1 0 35052 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0824_
timestamp 1649977179
transform 1 0 35604 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1649977179
transform 1 0 35696 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0826_
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0827_
timestamp 1649977179
transform 1 0 35512 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0828_
timestamp 1649977179
transform 1 0 41308 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1649977179
transform 1 0 34224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0830_
timestamp 1649977179
transform 1 0 41676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0831_
timestamp 1649977179
transform 1 0 40020 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0832_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 54280 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  _0833_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0834_
timestamp 1649977179
transform 1 0 47564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0836_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 48760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _0837_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 68172 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0838_
timestamp 1649977179
transform 1 0 33856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0839_
timestamp 1649977179
transform 1 0 42688 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _0840_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43884 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _0841_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 85192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0842_
timestamp 1649977179
transform 1 0 71668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 1649977179
transform 1 0 71852 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0844_
timestamp 1649977179
transform 1 0 73324 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1649977179
transform 1 0 46920 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0846_
timestamp 1649977179
transform 1 0 45172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0847_
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1649977179
transform 1 0 40664 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0849_
timestamp 1649977179
transform 1 0 47288 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0850_
timestamp 1649977179
transform 1 0 37904 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0851_
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0852_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 46276 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0853_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 64768 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0854_
timestamp 1649977179
transform 1 0 43884 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0855_
timestamp 1649977179
transform 1 0 43608 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0856_
timestamp 1649977179
transform 1 0 63940 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0857_
timestamp 1649977179
transform 1 0 45356 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0858_
timestamp 1649977179
transform 1 0 45356 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0859_
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0860_
timestamp 1649977179
transform 1 0 36616 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0861_
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0862_
timestamp 1649977179
transform 1 0 36248 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _0863_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _0864_
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0865_
timestamp 1649977179
transform 1 0 38732 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0866_
timestamp 1649977179
transform 1 0 63296 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0867_
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0868_
timestamp 1649977179
transform 1 0 37812 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0869_
timestamp 1649977179
transform 1 0 39744 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0870_
timestamp 1649977179
transform 1 0 37352 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0871_
timestamp 1649977179
transform 1 0 36248 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0872_
timestamp 1649977179
transform 1 0 45540 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0873_
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0874_
timestamp 1649977179
transform 1 0 39100 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0875_
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0876_
timestamp 1649977179
transform 1 0 62008 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0877_
timestamp 1649977179
transform 1 0 64216 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0878_
timestamp 1649977179
transform 1 0 56856 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0879_
timestamp 1649977179
transform 1 0 58696 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0880_
timestamp 1649977179
transform 1 0 58328 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0881_
timestamp 1649977179
transform 1 0 61364 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0882_
timestamp 1649977179
transform 1 0 63112 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0883_
timestamp 1649977179
transform 1 0 62008 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0884_
timestamp 1649977179
transform 1 0 48484 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0885_
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0886_
timestamp 1649977179
transform 1 0 48760 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0887_
timestamp 1649977179
transform 1 0 62192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0888_
timestamp 1649977179
transform 1 0 63756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0889_
timestamp 1649977179
transform 1 0 63848 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0890_
timestamp 1649977179
transform 1 0 60812 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0891_
timestamp 1649977179
transform 1 0 64676 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1649977179
transform 1 0 66884 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0893_
timestamp 1649977179
transform 1 0 61732 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0894_
timestamp 1649977179
transform 1 0 65596 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0895_
timestamp 1649977179
transform 1 0 60720 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0896_
timestamp 1649977179
transform 1 0 62284 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0897_
timestamp 1649977179
transform 1 0 55936 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0898_
timestamp 1649977179
transform 1 0 55752 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0899_
timestamp 1649977179
transform 1 0 56304 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0900_
timestamp 1649977179
transform 1 0 56580 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 1649977179
transform 1 0 56396 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0902_
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0903_
timestamp 1649977179
transform 1 0 33396 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0904_
timestamp 1649977179
transform 1 0 34868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0905_
timestamp 1649977179
transform 1 0 33396 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0906_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 71116 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0907_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 69276 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0908_
timestamp 1649977179
transform 1 0 70012 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0909_
timestamp 1649977179
transform 1 0 68724 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0910_
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0911_
timestamp 1649977179
transform 1 0 68908 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0912_
timestamp 1649977179
transform 1 0 67252 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0913_
timestamp 1649977179
transform 1 0 64308 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0914_
timestamp 1649977179
transform 1 0 64216 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0915_
timestamp 1649977179
transform 1 0 64400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 1649977179
transform 1 0 63204 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0917_
timestamp 1649977179
transform 1 0 44804 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0918_
timestamp 1649977179
transform 1 0 47012 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0919_
timestamp 1649977179
transform 1 0 46460 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0920_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43976 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0922_
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0923_
timestamp 1649977179
transform 1 0 32660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0924_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27876 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0925_
timestamp 1649977179
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0926_
timestamp 1649977179
transform 1 0 51244 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0927_
timestamp 1649977179
transform 1 0 51428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0928_
timestamp 1649977179
transform 1 0 50140 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0929_
timestamp 1649977179
transform 1 0 49404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0930_
timestamp 1649977179
transform 1 0 38916 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1649977179
transform 1 0 37720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0932_
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0933_
timestamp 1649977179
transform 1 0 39192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0934_
timestamp 1649977179
transform 1 0 33856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0935_
timestamp 1649977179
transform 1 0 32384 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 1649977179
transform 1 0 29256 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1649977179
transform 1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 1649977179
transform 1 0 38548 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1649977179
transform 1 0 37996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 1649977179
transform 1 0 28612 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 1649977179
transform 1 0 29716 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1649977179
transform 1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0944_
timestamp 1649977179
transform 1 0 38640 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0945_
timestamp 1649977179
transform 1 0 38640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0946_
timestamp 1649977179
transform 1 0 33028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0947_
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0948_
timestamp 1649977179
transform 1 0 26128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0949_
timestamp 1649977179
transform 1 0 24380 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0950_
timestamp 1649977179
transform 1 0 25024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0951_
timestamp 1649977179
transform 1 0 24196 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0952_
timestamp 1649977179
transform 1 0 24748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0953_
timestamp 1649977179
transform 1 0 33396 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0955_
timestamp 1649977179
transform 1 0 33948 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0956_
timestamp 1649977179
transform 1 0 33396 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0957_
timestamp 1649977179
transform 1 0 31188 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0958_
timestamp 1649977179
transform 1 0 68172 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp 1649977179
transform 1 0 27968 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 1649977179
transform 1 0 27416 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0962_
timestamp 1649977179
transform 1 0 23920 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0963_
timestamp 1649977179
transform 1 0 25024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0964_
timestamp 1649977179
transform 1 0 66976 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 1649977179
transform 1 0 67896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0966_
timestamp 1649977179
transform 1 0 49128 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0967_
timestamp 1649977179
transform 1 0 50232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0968_
timestamp 1649977179
transform 1 0 32108 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0969_
timestamp 1649977179
transform 1 0 24196 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0970_
timestamp 1649977179
transform 1 0 24932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 1649977179
transform 1 0 56948 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0972_
timestamp 1649977179
transform 1 0 56580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0974_
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0975_
timestamp 1649977179
transform 1 0 23552 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0976_
timestamp 1649977179
transform 1 0 24748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0977_
timestamp 1649977179
transform 1 0 70104 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0978_
timestamp 1649977179
transform 1 0 70748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0979_
timestamp 1649977179
transform 1 0 32384 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0980_
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0981_
timestamp 1649977179
transform 1 0 25576 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0982_
timestamp 1649977179
transform 1 0 35604 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1649977179
transform 1 0 35052 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0984_
timestamp 1649977179
transform 1 0 27600 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1649977179
transform 1 0 29072 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0986_
timestamp 1649977179
transform 1 0 25668 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1649977179
transform 1 0 26036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0988_
timestamp 1649977179
transform 1 0 27416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp 1649977179
transform 1 0 27140 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1649977179
transform 1 0 27600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0992_
timestamp 1649977179
transform 1 0 47104 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1649977179
transform 1 0 46920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1649977179
transform 1 0 45540 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0995_
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1649977179
transform 1 0 24472 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0997_
timestamp 1649977179
transform 1 0 28612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0998_
timestamp 1649977179
transform 1 0 27784 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0999_
timestamp 1649977179
transform 1 0 27968 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1000_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25760 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1649977179
transform 1 0 27324 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1002_
timestamp 1649977179
transform 1 0 27508 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1003_
timestamp 1649977179
transform 1 0 25668 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1004_
timestamp 1649977179
transform 1 0 24932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1005_
timestamp 1649977179
transform 1 0 25760 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1649977179
transform 1 0 25024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1649977179
transform 1 0 28520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1008_
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1009_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26496 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1649977179
transform 1 0 25208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1649977179
transform 1 0 26312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1012_
timestamp 1649977179
transform 1 0 40756 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1013_
timestamp 1649977179
transform 1 0 25760 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1014_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1015_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1016_
timestamp 1649977179
transform 1 0 19872 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1017_
timestamp 1649977179
transform 1 0 20608 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _1018_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1649977179
transform 1 0 23092 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1020_
timestamp 1649977179
transform 1 0 23092 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1021_
timestamp 1649977179
transform 1 0 18952 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1022_
timestamp 1649977179
transform 1 0 20884 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _1023_
timestamp 1649977179
transform 1 0 20792 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1024_
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1025_
timestamp 1649977179
transform 1 0 18124 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1026_
timestamp 1649977179
transform 1 0 18584 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _1027_
timestamp 1649977179
transform 1 0 19412 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1028_
timestamp 1649977179
transform 1 0 22724 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1029_
timestamp 1649977179
transform 1 0 21988 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1030_
timestamp 1649977179
transform 1 0 22816 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _1031_
timestamp 1649977179
transform 1 0 23552 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1032_
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1649977179
transform 1 0 20516 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1034_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1649977179
transform 1 0 14996 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1649977179
transform 1 0 24380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1037_
timestamp 1649977179
transform 1 0 25944 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1649977179
transform 1 0 23736 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1649977179
transform 1 0 24656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1040_
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1041_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25208 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1649977179
transform 1 0 24288 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1044_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21988 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1045_
timestamp 1649977179
transform 1 0 24104 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1046_
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1047_
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _1048_
timestamp 1649977179
transform 1 0 23460 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1049_
timestamp 1649977179
transform 1 0 22448 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1050_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25576 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1051_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 46368 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1052_
timestamp 1649977179
transform 1 0 48392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1053_
timestamp 1649977179
transform 1 0 30912 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1054_
timestamp 1649977179
transform 1 0 31556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1055_
timestamp 1649977179
transform 1 0 54096 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1056_
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1057_
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1058_
timestamp 1649977179
transform 1 0 30912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1059_
timestamp 1649977179
transform 1 0 55016 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1060_
timestamp 1649977179
transform 1 0 54464 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1061_
timestamp 1649977179
transform 1 0 41216 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1062_
timestamp 1649977179
transform 1 0 43332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1063_
timestamp 1649977179
transform 1 0 48116 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1064_
timestamp 1649977179
transform 1 0 46460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1065_
timestamp 1649977179
transform 1 0 52440 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1066_
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1067_
timestamp 1649977179
transform 1 0 46092 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1649977179
transform 1 0 45816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1069_
timestamp 1649977179
transform 1 0 60996 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 1649977179
transform 1 0 62100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1071_
timestamp 1649977179
transform 1 0 42780 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1649977179
transform 1 0 40020 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1073_
timestamp 1649977179
transform 1 0 37628 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1074_
timestamp 1649977179
transform 1 0 70748 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1649977179
transform 1 0 67804 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1076_
timestamp 1649977179
transform 1 0 71208 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1077_
timestamp 1649977179
transform 1 0 72496 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1078_
timestamp 1649977179
transform 1 0 71576 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1079_
timestamp 1649977179
transform 1 0 71852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1080_
timestamp 1649977179
transform 1 0 33120 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1081_
timestamp 1649977179
transform 1 0 31464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1082_
timestamp 1649977179
transform 1 0 29716 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1083_
timestamp 1649977179
transform 1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1084_
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1085_
timestamp 1649977179
transform 1 0 51520 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1649977179
transform 1 0 53268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1087_
timestamp 1649977179
transform 1 0 40296 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1649977179
transform 1 0 40020 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1089_
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1091_
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1649977179
transform 1 0 59800 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1093_
timestamp 1649977179
transform 1 0 57408 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1649977179
transform 1 0 57040 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1095_
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1096_
timestamp 1649977179
transform 1 0 35880 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1097_
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1098_
timestamp 1649977179
transform 1 0 42780 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1099_
timestamp 1649977179
transform 1 0 42136 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1100_
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1101_
timestamp 1649977179
transform 1 0 52164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1102_
timestamp 1649977179
transform 1 0 35972 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1103_
timestamp 1649977179
transform 1 0 35972 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1104_
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1105_
timestamp 1649977179
transform 1 0 49036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1106_
timestamp 1649977179
transform 1 0 41860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1107_
timestamp 1649977179
transform 1 0 65780 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1108_
timestamp 1649977179
transform 1 0 64952 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1109_
timestamp 1649977179
transform 1 0 70748 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1110_
timestamp 1649977179
transform 1 0 70104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1111_
timestamp 1649977179
transform 1 0 69000 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1112_
timestamp 1649977179
transform 1 0 68724 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1113_
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1114_
timestamp 1649977179
transform 1 0 31464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1115_
timestamp 1649977179
transform 1 0 31648 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1116_
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1117_
timestamp 1649977179
transform 1 0 37904 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1118_
timestamp 1649977179
transform 1 0 37076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1119_
timestamp 1649977179
transform 1 0 36248 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1120_
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1121_
timestamp 1649977179
transform 1 0 33120 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1123_
timestamp 1649977179
transform 1 0 44160 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1124_
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1125_
timestamp 1649977179
transform 1 0 57040 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1126_
timestamp 1649977179
transform 1 0 55936 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1127_
timestamp 1649977179
transform 1 0 47564 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1128_
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1129_
timestamp 1649977179
transform 1 0 61456 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1130_
timestamp 1649977179
transform 1 0 64584 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1131_
timestamp 1649977179
transform 1 0 59064 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1132_
timestamp 1649977179
transform 1 0 57224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1133_
timestamp 1649977179
transform 1 0 50784 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1134_
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1135_
timestamp 1649977179
transform 1 0 51520 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1136_
timestamp 1649977179
transform 1 0 52072 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1137_
timestamp 1649977179
transform 1 0 50416 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1138_
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1139_
timestamp 1649977179
transform 1 0 59156 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1140_
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1141_
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1142_
timestamp 1649977179
transform 1 0 62192 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1143_
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1649977179
transform 1 0 66148 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1145_
timestamp 1649977179
transform 1 0 66884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1146_
timestamp 1649977179
transform 1 0 69092 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1147_
timestamp 1649977179
transform 1 0 67528 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1148_
timestamp 1649977179
transform 1 0 71576 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1649977179
transform 1 0 68540 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1150_
timestamp 1649977179
transform 1 0 58788 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1151_
timestamp 1649977179
transform 1 0 59248 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1152_
timestamp 1649977179
transform 1 0 55844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1153_
timestamp 1649977179
transform 1 0 63020 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1154_
timestamp 1649977179
transform 1 0 63756 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1155_
timestamp 1649977179
transform 1 0 64676 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1156_
timestamp 1649977179
transform 1 0 64676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1157_
timestamp 1649977179
transform 1 0 64768 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1158_
timestamp 1649977179
transform 1 0 64308 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1159_
timestamp 1649977179
transform 1 0 59524 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1160_
timestamp 1649977179
transform 1 0 59800 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1161_
timestamp 1649977179
transform 1 0 43056 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1162_
timestamp 1649977179
transform 1 0 57868 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1163_
timestamp 1649977179
transform 1 0 57224 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1164_
timestamp 1649977179
transform 1 0 50600 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1165_
timestamp 1649977179
transform 1 0 51336 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1166_
timestamp 1649977179
transform 1 0 44160 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1167_
timestamp 1649977179
transform 1 0 44804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1168_
timestamp 1649977179
transform 1 0 47656 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1649977179
transform 1 0 47564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1170_
timestamp 1649977179
transform 1 0 41584 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1171_
timestamp 1649977179
transform 1 0 41308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1172_
timestamp 1649977179
transform 1 0 45632 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1173_
timestamp 1649977179
transform 1 0 44344 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1174_
timestamp 1649977179
transform 1 0 45080 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1175_
timestamp 1649977179
transform 1 0 56120 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1176_
timestamp 1649977179
transform 1 0 57040 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1177_
timestamp 1649977179
transform 1 0 56028 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1178_
timestamp 1649977179
transform 1 0 56764 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1179_
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1180_
timestamp 1649977179
transform 1 0 45632 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1181_
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1182_
timestamp 1649977179
transform 1 0 54372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1183_
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1184_
timestamp 1649977179
transform 1 0 36432 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1185_
timestamp 1649977179
transform 1 0 38088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1186_
timestamp 1649977179
transform 1 0 33120 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1187_
timestamp 1649977179
transform 1 0 33028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1188_
timestamp 1649977179
transform 1 0 34960 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1189_
timestamp 1649977179
transform 1 0 34224 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1190_
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1191_
timestamp 1649977179
transform 1 0 33672 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1192_
timestamp 1649977179
transform 1 0 41400 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1193_
timestamp 1649977179
transform 1 0 42320 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1194_
timestamp 1649977179
transform 1 0 50232 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1195_
timestamp 1649977179
transform 1 0 51060 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1196_
timestamp 1649977179
transform 1 0 47932 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1197_
timestamp 1649977179
transform 1 0 47840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1198_
timestamp 1649977179
transform 1 0 45540 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1199_
timestamp 1649977179
transform 1 0 44344 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1200_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 70748 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1201_
timestamp 1649977179
transform 1 0 69184 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 1649977179
transform 1 0 67804 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp 1649977179
transform 1 0 65504 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1204_
timestamp 1649977179
transform 1 0 63756 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1205_
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp 1649977179
transform 1 0 45264 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp 1649977179
transform 1 0 42228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1208_
timestamp 1649977179
transform 1 0 27784 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1209_
timestamp 1649977179
transform 1 0 51520 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1210_
timestamp 1649977179
transform 1 0 49588 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1211_
timestamp 1649977179
transform 1 0 39376 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1212_
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1213_
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1214_
timestamp 1649977179
transform 1 0 40296 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1215_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1216_
timestamp 1649977179
transform 1 0 29716 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1217_
timestamp 1649977179
transform 1 0 38548 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1218_
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1219_
timestamp 1649977179
transform 1 0 25760 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1220_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25300 0 1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1221_
timestamp 1649977179
transform 1 0 32292 0 -1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1222_
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1223_
timestamp 1649977179
transform 1 0 68724 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1224_
timestamp 1649977179
transform 1 0 27324 0 1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1225_
timestamp 1649977179
transform 1 0 25024 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1226_
timestamp 1649977179
transform 1 0 68540 0 1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1227_
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1228_
timestamp 1649977179
transform 1 0 25668 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1229_
timestamp 1649977179
transform 1 0 55752 0 -1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1230_
timestamp 1649977179
transform 1 0 26128 0 1 4352
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1231_
timestamp 1649977179
transform 1 0 25576 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1232_
timestamp 1649977179
transform 1 0 69644 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1233_
timestamp 1649977179
transform 1 0 26680 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1234_
timestamp 1649977179
transform 1 0 36064 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1235_
timestamp 1649977179
transform 1 0 27232 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1236_
timestamp 1649977179
transform 1 0 26036 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1237_
timestamp 1649977179
transform 1 0 25024 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1238_
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1239_
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 1649977179
transform 1 0 45816 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 1649977179
transform 1 0 66424 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 1649977179
transform 1 0 32016 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 1649977179
transform 1 0 32752 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 1649977179
transform 1 0 54372 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 1649977179
transform 1 0 46368 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 1649977179
transform 1 0 52900 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 1649977179
transform 1 0 60812 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1649977179
transform 1 0 42228 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1649977179
transform 1 0 68908 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 1649977179
transform 1 0 70748 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 1649977179
transform 1 0 69828 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 1649977179
transform 1 0 33304 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 1649977179
transform 1 0 39560 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp 1649977179
transform 1 0 41492 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 1649977179
transform 1 0 59432 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 1649977179
transform 1 0 56580 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 1649977179
transform 1 0 36524 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 1649977179
transform 1 0 42688 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 1649977179
transform 1 0 52716 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 1649977179
transform 1 0 49588 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 1649977179
transform 1 0 65596 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 1649977179
transform 1 0 68908 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 1649977179
transform 1 0 68356 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp 1649977179
transform 1 0 31188 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp 1649977179
transform 1 0 31004 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp 1649977179
transform 1 0 35144 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp 1649977179
transform 1 0 32476 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1275_
timestamp 1649977179
transform 1 0 69644 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp 1649977179
transform 1 0 44804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1277_
timestamp 1649977179
transform 1 0 55476 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp 1649977179
transform 1 0 58328 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1280_
timestamp 1649977179
transform 1 0 51152 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1281_
timestamp 1649977179
transform 1 0 51612 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1649977179
transform 1 0 50324 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp 1649977179
transform 1 0 62192 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1649977179
transform 1 0 66516 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1286_
timestamp 1649977179
transform 1 0 69368 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1649977179
transform 1 0 69828 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1649977179
transform 1 0 58604 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp 1649977179
transform 1 0 62928 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1649977179
transform 1 0 64308 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1649977179
transform 1 0 65596 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp 1649977179
transform 1 0 60260 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp 1649977179
transform 1 0 58604 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp 1649977179
transform 1 0 44804 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1649977179
transform 1 0 41860 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp 1649977179
transform 1 0 42688 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1649977179
transform 1 0 55108 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1649977179
transform 1 0 45724 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1649977179
transform 1 0 54096 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1304_
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1305_
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1306_
timestamp 1649977179
transform 1 0 33304 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1307_
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1308_
timestamp 1649977179
transform 1 0 49404 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1309_
timestamp 1649977179
transform 1 0 47932 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1310_
timestamp 1649977179
transform 1 0 43792 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1321_
timestamp 1649977179
transform 1 0 42688 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1322_
timestamp 1649977179
transform 1 0 2852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1649977179
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1324_
timestamp 1649977179
transform 1 0 64308 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1325_
timestamp 1649977179
transform 1 0 25760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1649977179
transform 1 0 53912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1327_
timestamp 1649977179
transform 1 0 73600 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1328_
timestamp 1649977179
transform 1 0 57868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1329_
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1330_
timestamp 1649977179
transform 1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1649977179
transform 1 0 65412 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1332_
timestamp 1649977179
transform 1 0 53268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1333_
timestamp 1649977179
transform 1 0 85928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1334_
timestamp 1649977179
transform 1 0 19780 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1335_
timestamp 1649977179
transform 1 0 53636 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1336_
timestamp 1649977179
transform 1 0 38456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1337_
timestamp 1649977179
transform 1 0 86756 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1338_
timestamp 1649977179
transform 1 0 58420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1339_
timestamp 1649977179
transform 1 0 68540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1340_
timestamp 1649977179
transform 1 0 9752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1341_
timestamp 1649977179
transform 1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1342_
timestamp 1649977179
transform 1 0 86756 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1343_
timestamp 1649977179
transform 1 0 70104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1344_
timestamp 1649977179
transform 1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1345_
timestamp 1649977179
transform 1 0 26680 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1346_
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1347_
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1348_
timestamp 1649977179
transform 1 0 20332 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1349_
timestamp 1649977179
transform 1 0 86756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1649977179
transform 1 0 36432 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1649977179
transform 1 0 39008 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1649977179
transform 1 0 36432 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1649977179
transform 1 0 39008 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1649977179
transform 1 0 51980 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1649977179
transform 1 0 54556 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1649977179
transform 1 0 59800 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1649977179
transform 1 0 59800 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1649977179
transform 1 0 16652 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 71300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform 1 0 87400 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1649977179
transform 1 0 12788 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1649977179
transform 1 0 32936 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1649977179
transform 1 0 1656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 41768 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform 1 0 87400 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 69000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform 1 0 6624 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 60444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 38732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 55844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1649977179
transform 1 0 11592 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 48116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1649977179
transform 1 0 87400 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 88044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 84180 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform 1 0 23920 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 21160 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1649977179
transform 1 0 85100 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 4600 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1649977179
transform 1 0 87952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 45172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 51612 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1649977179
transform 1 0 87400 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1649977179
transform 1 0 30820 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform 1 0 54188 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1649977179
transform 1 0 80040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 48668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform 1 0 44344 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 70748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform 1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 67252 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform 1 0 49036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 53544 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform 1 0 87400 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform 1 0 88044 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform 1 0 36616 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform 1 0 28336 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 16836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1649977179
transform 1 0 82524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1649977179
transform 1 0 63204 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform 1 0 51980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1649977179
transform 1 0 86756 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1649977179
transform 1 0 1656 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input61
timestamp 1649977179
transform 1 0 85100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1649977179
transform 1 0 23092 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1649977179
transform 1 0 68448 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1649977179
transform 1 0 69092 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1649977179
transform 1 0 55292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1649977179
transform 1 0 87952 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input68
timestamp 1649977179
transform 1 0 79396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1649977179
transform 1 0 49404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1649977179
transform 1 0 30360 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1649977179
transform 1 0 80592 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1649977179
transform 1 0 32108 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input74
timestamp 1649977179
transform 1 0 87768 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1649977179
transform 1 0 12788 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1649977179
transform 1 0 51244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1649977179
transform 1 0 61272 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1649977179
transform 1 0 87952 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1649977179
transform 1 0 10212 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1649977179
transform 1 0 58696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input82
timestamp 1649977179
transform 1 0 87952 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1649977179
transform 1 0 6348 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1649977179
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input85
timestamp 1649977179
transform 1 0 72220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input87
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input88
timestamp 1649977179
transform 1 0 87768 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1649977179
transform 1 0 44344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1649977179
transform 1 0 48392 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1649977179
transform 1 0 82524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1649977179
transform 1 0 81328 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input94
timestamp 1649977179
transform 1 0 87400 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1649977179
transform 1 0 61272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input96
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1649977179
transform 1 0 87952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input98
timestamp 1649977179
transform 1 0 1472 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input99
timestamp 1649977179
transform 1 0 87952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1649977179
transform 1 0 78752 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input101
timestamp 1649977179
transform 1 0 64492 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1649977179
transform 1 0 76176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1649977179
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input105
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1649977179
transform 1 0 46276 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1649977179
transform 1 0 25852 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1649977179
transform 1 0 49680 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input111
timestamp 1649977179
transform 1 0 1656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input113
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input114
timestamp 1649977179
transform 1 0 63848 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1649977179
transform 1 0 50416 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1649977179
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 1649977179
transform 1 0 73600 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1649977179
transform 1 0 74796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input119
timestamp 1649977179
transform 1 0 12328 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1649977179
transform 1 0 87952 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input121
timestamp 1649977179
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input122
timestamp 1649977179
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input123
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  l1icache_32_318 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  l1icache_32_319
timestamp 1649977179
transform 1 0 84456 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  l1icache_32_320
timestamp 1649977179
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  l1icache_32_321
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  l1icache_32_322
timestamp 1649977179
transform 1 0 87860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  l1icache_32_323
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  l1icache_32_324
timestamp 1649977179
transform 1 0 74152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  l1icache_32_325
timestamp 1649977179
transform 1 0 8280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  l1icache_32_326
timestamp 1649977179
transform 1 0 59524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  l1icache_32_327
timestamp 1649977179
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output124
timestamp 1649977179
transform 1 0 5244 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output125
timestamp 1649977179
transform 1 0 88044 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output126
timestamp 1649977179
transform 1 0 35512 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output127
timestamp 1649977179
transform 1 0 88044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output128
timestamp 1649977179
transform 1 0 14904 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output129
timestamp 1649977179
transform 1 0 72404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output130
timestamp 1649977179
transform 1 0 56948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output131
timestamp 1649977179
transform 1 0 42596 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output132
timestamp 1649977179
transform 1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output133
timestamp 1649977179
transform 1 0 10396 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output134
timestamp 1649977179
transform 1 0 57868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output135
timestamp 1649977179
transform 1 0 52716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output136
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output137
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output138
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output139
timestamp 1649977179
transform 1 0 2576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output140
timestamp 1649977179
transform 1 0 61916 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output141
timestamp 1649977179
transform 1 0 45816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output142
timestamp 1649977179
transform 1 0 69644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output143
timestamp 1649977179
transform 1 0 88320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output144
timestamp 1649977179
transform 1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output145
timestamp 1649977179
transform 1 0 71852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output146
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output147
timestamp 1649977179
transform 1 0 33488 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output148
timestamp 1649977179
transform 1 0 20056 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output149
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output150
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output151
timestamp 1649977179
transform 1 0 65596 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output152
timestamp 1649977179
transform 1 0 7268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output153
timestamp 1649977179
transform 1 0 38732 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output154
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output155
timestamp 1649977179
transform 1 0 77372 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output156
timestamp 1649977179
transform 1 0 86940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output157
timestamp 1649977179
transform 1 0 36064 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output158
timestamp 1649977179
transform 1 0 88044 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output159
timestamp 1649977179
transform 1 0 81972 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output160
timestamp 1649977179
transform 1 0 88044 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output161
timestamp 1649977179
transform 1 0 83628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output162
timestamp 1649977179
transform 1 0 15548 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output163
timestamp 1649977179
transform 1 0 74244 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output164
timestamp 1649977179
transform 1 0 73324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output165
timestamp 1649977179
transform 1 0 87400 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output166
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output167
timestamp 1649977179
transform 1 0 74796 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output168
timestamp 1649977179
transform 1 0 88044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output169
timestamp 1649977179
transform 1 0 26312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output170
timestamp 1649977179
transform 1 0 43792 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output171
timestamp 1649977179
transform 1 0 66148 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output172
timestamp 1649977179
transform 1 0 88044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output173
timestamp 1649977179
transform 1 0 45172 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output174
timestamp 1649977179
transform 1 0 86204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output175
timestamp 1649977179
transform 1 0 9108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output176
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output177
timestamp 1649977179
transform 1 0 88044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output178
timestamp 1649977179
transform 1 0 73324 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output179
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output180
timestamp 1649977179
transform 1 0 88044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output181
timestamp 1649977179
transform 1 0 86848 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output182
timestamp 1649977179
transform 1 0 70748 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output183
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output184
timestamp 1649977179
transform 1 0 59340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output185
timestamp 1649977179
transform 1 0 88044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output186
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output187
timestamp 1649977179
transform 1 0 86848 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output188
timestamp 1649977179
transform 1 0 63020 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output189
timestamp 1649977179
transform 1 0 36616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output190
timestamp 1649977179
transform 1 0 61916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output191
timestamp 1649977179
transform 1 0 86388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output192
timestamp 1649977179
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output193
timestamp 1649977179
transform 1 0 51060 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output194
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output195
timestamp 1649977179
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output196
timestamp 1649977179
transform 1 0 34592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output197
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output198
timestamp 1649977179
transform 1 0 88044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output199
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output200
timestamp 1649977179
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output201
timestamp 1649977179
transform 1 0 21988 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output202
timestamp 1649977179
transform 1 0 88044 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output203
timestamp 1649977179
transform 1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output204
timestamp 1649977179
transform 1 0 51888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output205
timestamp 1649977179
transform 1 0 75440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output206
timestamp 1649977179
transform 1 0 80224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output207
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output208
timestamp 1649977179
transform 1 0 56764 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output209
timestamp 1649977179
transform 1 0 86204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output210
timestamp 1649977179
transform 1 0 81696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output211
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output212
timestamp 1649977179
transform 1 0 49036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output213
timestamp 1649977179
transform 1 0 88044 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output214
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output215
timestamp 1649977179
transform 1 0 66148 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output216
timestamp 1649977179
transform 1 0 60628 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output217
timestamp 1649977179
transform 1 0 63020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output218
timestamp 1649977179
transform 1 0 56120 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output219
timestamp 1649977179
transform 1 0 41216 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output220
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output221
timestamp 1649977179
transform 1 0 67252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output222
timestamp 1649977179
transform 1 0 84456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output223
timestamp 1649977179
transform 1 0 77372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output224
timestamp 1649977179
transform 1 0 37444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output225
timestamp 1649977179
transform 1 0 46460 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output226
timestamp 1649977179
transform 1 0 36064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output227
timestamp 1649977179
transform 1 0 43792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output228
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output229
timestamp 1649977179
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output230
timestamp 1649977179
transform 1 0 40020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output231
timestamp 1649977179
transform 1 0 76544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output232
timestamp 1649977179
transform 1 0 43240 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output233
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output234
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output235
timestamp 1649977179
transform 1 0 81880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output236
timestamp 1649977179
transform 1 0 34040 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output237
timestamp 1649977179
transform 1 0 14260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output238
timestamp 1649977179
transform 1 0 2668 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output239
timestamp 1649977179
transform 1 0 79304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output240
timestamp 1649977179
transform 1 0 88044 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output241
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output242
timestamp 1649977179
transform 1 0 32936 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output243
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output244
timestamp 1649977179
transform 1 0 88320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output245
timestamp 1649977179
transform 1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output246
timestamp 1649977179
transform 1 0 88044 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output247
timestamp 1649977179
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output248
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output249
timestamp 1649977179
transform 1 0 64860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output250
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output251
timestamp 1649977179
transform 1 0 54188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output252
timestamp 1649977179
transform 1 0 88044 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output253
timestamp 1649977179
transform 1 0 58420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output254
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output255
timestamp 1649977179
transform 1 0 18032 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output256
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output257
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output258
timestamp 1649977179
transform 1 0 88044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output259
timestamp 1649977179
transform 1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output260
timestamp 1649977179
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output261
timestamp 1649977179
transform 1 0 3956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output262
timestamp 1649977179
transform 1 0 79028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output263
timestamp 1649977179
transform 1 0 38088 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output264
timestamp 1649977179
transform 1 0 58788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output265
timestamp 1649977179
transform 1 0 66700 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output266
timestamp 1649977179
transform 1 0 53544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output267
timestamp 1649977179
transform 1 0 87308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output268
timestamp 1649977179
transform 1 0 18584 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output269
timestamp 1649977179
transform 1 0 52900 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output270
timestamp 1649977179
transform 1 0 41032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output271
timestamp 1649977179
transform 1 0 88044 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output272
timestamp 1649977179
transform 1 0 58972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output273
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output274
timestamp 1649977179
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output275
timestamp 1649977179
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output276
timestamp 1649977179
transform 1 0 60444 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output277
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output278
timestamp 1649977179
transform 1 0 2760 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output279
timestamp 1649977179
transform 1 0 21160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output280
timestamp 1649977179
transform 1 0 7728 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output281
timestamp 1649977179
transform 1 0 79948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output282
timestamp 1649977179
transform 1 0 43240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output283
timestamp 1649977179
transform 1 0 83628 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output284
timestamp 1649977179
transform 1 0 41768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output285
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output286
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output287
timestamp 1649977179
transform 1 0 56396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output288
timestamp 1649977179
transform 1 0 71944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output289
timestamp 1649977179
transform 1 0 57868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output290
timestamp 1649977179
transform 1 0 88044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output291
timestamp 1649977179
transform 1 0 25300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output292
timestamp 1649977179
transform 1 0 29716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output293
timestamp 1649977179
transform 1 0 27784 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output294
timestamp 1649977179
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output295
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output296
timestamp 1649977179
transform 1 0 86848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output297
timestamp 1649977179
transform 1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output298
timestamp 1649977179
transform 1 0 76820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output299
timestamp 1649977179
transform 1 0 86296 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output300
timestamp 1649977179
transform 1 0 40664 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output301
timestamp 1649977179
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output302
timestamp 1649977179
transform 1 0 3128 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output303
timestamp 1649977179
transform 1 0 87492 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output304
timestamp 1649977179
transform 1 0 13616 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output305
timestamp 1649977179
transform 1 0 88044 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output306
timestamp 1649977179
transform 1 0 75900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output307
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output308
timestamp 1649977179
transform 1 0 27324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output309
timestamp 1649977179
transform 1 0 88044 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output310
timestamp 1649977179
transform 1 0 71300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output311
timestamp 1649977179
transform 1 0 69644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output312
timestamp 1649977179
transform 1 0 27140 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output313
timestamp 1649977179
transform 1 0 37444 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output314
timestamp 1649977179
transform 1 0 42596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output315
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output316
timestamp 1649977179
transform 1 0 20608 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output317
timestamp 1649977179
transform 1 0 87492 0 -1 4352
box -38 -48 314 592
<< labels >>
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 5170 29200 5226 30000 0 FreeSans 224 90 0 0 data_chip_en
port 1 nsew signal tristate
flabel metal3 s 89200 7488 90000 7608 0 FreeSans 480 0 0 0 data_in[0]
port 2 nsew signal tristate
flabel metal2 s 35438 29200 35494 30000 0 FreeSans 224 90 0 0 data_in[10]
port 3 nsew signal tristate
flabel metal3 s 89200 11568 90000 11688 0 FreeSans 480 0 0 0 data_in[11]
port 4 nsew signal tristate
flabel metal2 s 14830 29200 14886 30000 0 FreeSans 224 90 0 0 data_in[12]
port 5 nsew signal tristate
flabel metal2 s 72146 29200 72202 30000 0 FreeSans 224 90 0 0 data_in[13]
port 6 nsew signal tristate
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 data_in[14]
port 7 nsew signal tristate
flabel metal2 s 42522 29200 42578 30000 0 FreeSans 224 90 0 0 data_in[15]
port 8 nsew signal tristate
flabel metal2 s 34794 29200 34850 30000 0 FreeSans 224 90 0 0 data_in[16]
port 9 nsew signal tristate
flabel metal2 s 10322 29200 10378 30000 0 FreeSans 224 90 0 0 data_in[17]
port 10 nsew signal tristate
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 data_in[18]
port 11 nsew signal tristate
flabel metal2 s 52182 29200 52238 30000 0 FreeSans 224 90 0 0 data_in[19]
port 12 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 data_in[1]
port 13 nsew signal tristate
flabel metal2 s 662 29200 718 30000 0 FreeSans 224 90 0 0 data_in[20]
port 14 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 data_in[21]
port 15 nsew signal tristate
flabel metal2 s 18 29200 74 30000 0 FreeSans 224 90 0 0 data_in[22]
port 16 nsew signal tristate
flabel metal2 s 61842 29200 61898 30000 0 FreeSans 224 90 0 0 data_in[23]
port 17 nsew signal tristate
flabel metal2 s 45742 29200 45798 30000 0 FreeSans 224 90 0 0 data_in[24]
port 18 nsew signal tristate
flabel metal2 s 69570 0 69626 800 0 FreeSans 224 90 0 0 data_in[25]
port 19 nsew signal tristate
flabel metal2 s 87602 0 87658 800 0 FreeSans 224 90 0 0 data_in[26]
port 20 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 data_in[27]
port 21 nsew signal tristate
flabel metal2 s 71502 29200 71558 30000 0 FreeSans 224 90 0 0 data_in[28]
port 22 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 data_in[29]
port 23 nsew signal tristate
flabel metal2 s 33506 29200 33562 30000 0 FreeSans 224 90 0 0 data_in[2]
port 24 nsew signal tristate
flabel metal2 s 19982 29200 20038 30000 0 FreeSans 224 90 0 0 data_in[30]
port 25 nsew signal tristate
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 data_in[31]
port 26 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 data_in[3]
port 27 nsew signal tristate
flabel metal2 s 65062 29200 65118 30000 0 FreeSans 224 90 0 0 data_in[4]
port 28 nsew signal tristate
flabel metal2 s 7102 29200 7158 30000 0 FreeSans 224 90 0 0 data_in[5]
port 29 nsew signal tristate
flabel metal2 s 38658 29200 38714 30000 0 FreeSans 224 90 0 0 data_in[6]
port 30 nsew signal tristate
flabel metal2 s 39302 29200 39358 30000 0 FreeSans 224 90 0 0 data_in[7]
port 31 nsew signal tristate
flabel metal2 s 77298 29200 77354 30000 0 FreeSans 224 90 0 0 data_in[8]
port 32 nsew signal tristate
flabel metal2 s 89534 0 89590 800 0 FreeSans 224 90 0 0 data_in[9]
port 33 nsew signal tristate
flabel metal2 s 36082 29200 36138 30000 0 FreeSans 224 90 0 0 data_index[0]
port 34 nsew signal tristate
flabel metal3 s 89200 21088 90000 21208 0 FreeSans 480 0 0 0 data_index[1]
port 35 nsew signal tristate
flabel metal2 s 81806 29200 81862 30000 0 FreeSans 224 90 0 0 data_index[2]
port 36 nsew signal tristate
flabel metal3 s 89200 28568 90000 28688 0 FreeSans 480 0 0 0 data_index[3]
port 37 nsew signal tristate
flabel metal2 s 83094 0 83150 800 0 FreeSans 224 90 0 0 data_index[4]
port 38 nsew signal tristate
flabel metal2 s 15474 29200 15530 30000 0 FreeSans 224 90 0 0 data_index[5]
port 39 nsew signal tristate
flabel metal2 s 74078 29200 74134 30000 0 FreeSans 224 90 0 0 data_index[6]
port 40 nsew signal tristate
flabel metal2 s 72790 0 72846 800 0 FreeSans 224 90 0 0 data_index[7]
port 41 nsew signal tristate
flabel metal2 s 16118 29200 16174 30000 0 FreeSans 224 90 0 0 data_out[0]
port 42 nsew signal input
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 data_out[10]
port 43 nsew signal input
flabel metal3 s 89200 26528 90000 26648 0 FreeSans 480 0 0 0 data_out[11]
port 44 nsew signal input
flabel metal2 s 12898 29200 12954 30000 0 FreeSans 224 90 0 0 data_out[12]
port 45 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 data_out[13]
port 46 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 data_out[14]
port 47 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 data_out[15]
port 48 nsew signal input
flabel metal2 s 41878 29200 41934 30000 0 FreeSans 224 90 0 0 data_out[16]
port 49 nsew signal input
flabel metal3 s 89200 8848 90000 8968 0 FreeSans 480 0 0 0 data_out[17]
port 50 nsew signal input
flabel metal2 s 68926 0 68982 800 0 FreeSans 224 90 0 0 data_out[18]
port 51 nsew signal input
flabel metal2 s 6458 29200 6514 30000 0 FreeSans 224 90 0 0 data_out[19]
port 52 nsew signal input
flabel metal2 s 59910 0 59966 800 0 FreeSans 224 90 0 0 data_out[1]
port 53 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 data_out[20]
port 54 nsew signal input
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 data_out[21]
port 55 nsew signal input
flabel metal2 s 11610 29200 11666 30000 0 FreeSans 224 90 0 0 data_out[22]
port 56 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 data_out[23]
port 57 nsew signal input
flabel metal2 s 87602 29200 87658 30000 0 FreeSans 224 90 0 0 data_out[24]
port 58 nsew signal input
flabel metal3 s 89200 8168 90000 8288 0 FreeSans 480 0 0 0 data_out[25]
port 59 nsew signal input
flabel metal2 s 83738 29200 83794 30000 0 FreeSans 224 90 0 0 data_out[26]
port 60 nsew signal input
flabel metal2 s 23846 29200 23902 30000 0 FreeSans 224 90 0 0 data_out[27]
port 61 nsew signal input
flabel metal2 s 21270 29200 21326 30000 0 FreeSans 224 90 0 0 data_out[28]
port 62 nsew signal input
flabel metal2 s 85026 29200 85082 30000 0 FreeSans 224 90 0 0 data_out[29]
port 63 nsew signal input
flabel metal2 s 4526 29200 4582 30000 0 FreeSans 224 90 0 0 data_out[2]
port 64 nsew signal input
flabel metal3 s 89200 6808 90000 6928 0 FreeSans 480 0 0 0 data_out[30]
port 65 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 data_out[31]
port 66 nsew signal input
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 data_out[3]
port 67 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 data_out[4]
port 68 nsew signal input
flabel metal2 s 51538 29200 51594 30000 0 FreeSans 224 90 0 0 data_out[5]
port 69 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 data_out[6]
port 70 nsew signal input
flabel metal3 s 89200 10888 90000 11008 0 FreeSans 480 0 0 0 data_out[7]
port 71 nsew signal input
flabel metal2 s 30930 29200 30986 30000 0 FreeSans 224 90 0 0 data_out[8]
port 72 nsew signal input
flabel metal2 s 54114 29200 54170 30000 0 FreeSans 224 90 0 0 data_out[9]
port 73 nsew signal input
flabel metal2 s 88246 29200 88302 30000 0 FreeSans 224 90 0 0 data_write_en
port 74 nsew signal tristate
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 ld_data_o[0]
port 75 nsew signal tristate
flabel metal2 s 74722 29200 74778 30000 0 FreeSans 224 90 0 0 ld_data_o[10]
port 76 nsew signal tristate
flabel metal3 s 89200 2728 90000 2848 0 FreeSans 480 0 0 0 ld_data_o[11]
port 77 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 ld_data_o[12]
port 78 nsew signal tristate
flabel metal2 s 43810 29200 43866 30000 0 FreeSans 224 90 0 0 ld_data_o[13]
port 79 nsew signal tristate
flabel metal2 s 65706 0 65762 800 0 FreeSans 224 90 0 0 ld_data_o[14]
port 80 nsew signal tristate
flabel metal3 s 89200 19048 90000 19168 0 FreeSans 480 0 0 0 ld_data_o[15]
port 81 nsew signal tristate
flabel metal2 s 45098 29200 45154 30000 0 FreeSans 224 90 0 0 ld_data_o[16]
port 82 nsew signal tristate
flabel metal2 s 85670 0 85726 800 0 FreeSans 224 90 0 0 ld_data_o[17]
port 83 nsew signal tristate
flabel metal2 s 9034 29200 9090 30000 0 FreeSans 224 90 0 0 ld_data_o[18]
port 84 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 ld_data_o[19]
port 85 nsew signal tristate
flabel metal3 s 89200 13608 90000 13728 0 FreeSans 480 0 0 0 ld_data_o[1]
port 86 nsew signal tristate
flabel metal2 s 72790 29200 72846 30000 0 FreeSans 224 90 0 0 ld_data_o[20]
port 87 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 ld_data_o[21]
port 88 nsew signal tristate
flabel metal3 s 89200 4768 90000 4888 0 FreeSans 480 0 0 0 ld_data_o[22]
port 89 nsew signal tristate
flabel metal2 s 88890 29200 88946 30000 0 FreeSans 224 90 0 0 ld_data_o[23]
port 90 nsew signal tristate
flabel metal2 s 69570 29200 69626 30000 0 FreeSans 224 90 0 0 ld_data_o[24]
port 91 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 ld_data_o[25]
port 92 nsew signal tristate
flabel metal2 s 59266 29200 59322 30000 0 FreeSans 224 90 0 0 ld_data_o[26]
port 93 nsew signal tristate
flabel metal3 s 89200 4088 90000 4208 0 FreeSans 480 0 0 0 ld_data_o[27]
port 94 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 ld_data_o[28]
port 95 nsew signal tristate
flabel metal2 s 86958 29200 87014 30000 0 FreeSans 224 90 0 0 ld_data_o[29]
port 96 nsew signal tristate
flabel metal2 s 62486 29200 62542 30000 0 FreeSans 224 90 0 0 ld_data_o[2]
port 97 nsew signal tristate
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 ld_data_o[30]
port 98 nsew signal tristate
flabel metal2 s 61842 0 61898 800 0 FreeSans 224 90 0 0 ld_data_o[31]
port 99 nsew signal tristate
flabel metal3 s 89200 8 90000 128 0 FreeSans 480 0 0 0 ld_data_o[3]
port 100 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 ld_data_o[4]
port 101 nsew signal tristate
flabel metal2 s 50894 29200 50950 30000 0 FreeSans 224 90 0 0 ld_data_o[5]
port 102 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 ld_data_o[6]
port 103 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 ld_data_o[7]
port 104 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 ld_data_o[8]
port 105 nsew signal tristate
flabel metal2 s 65062 0 65118 800 0 FreeSans 224 90 0 0 ld_data_o[9]
port 106 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 req_addr_i[0]
port 107 nsew signal input
flabel metal2 s 79874 29200 79930 30000 0 FreeSans 224 90 0 0 req_addr_i[10]
port 108 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 req_addr_i[11]
port 109 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 req_addr_i[12]
port 110 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 req_addr_i[13]
port 111 nsew signal input
flabel metal2 s 44454 29200 44510 30000 0 FreeSans 224 90 0 0 req_addr_i[14]
port 112 nsew signal input
flabel metal2 s 70214 0 70270 800 0 FreeSans 224 90 0 0 req_addr_i[15]
port 113 nsew signal input
flabel metal2 s 28998 29200 29054 30000 0 FreeSans 224 90 0 0 req_addr_i[16]
port 114 nsew signal input
flabel metal2 s 22558 29200 22614 30000 0 FreeSans 224 90 0 0 req_addr_i[17]
port 115 nsew signal input
flabel metal2 s 66994 29200 67050 30000 0 FreeSans 224 90 0 0 req_addr_i[18]
port 116 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 req_addr_i[19]
port 117 nsew signal input
flabel metal2 s 53470 29200 53526 30000 0 FreeSans 224 90 0 0 req_addr_i[1]
port 118 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 req_addr_i[20]
port 119 nsew signal input
flabel metal3 s 89200 6128 90000 6248 0 FreeSans 480 0 0 0 req_addr_i[21]
port 120 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 req_addr_i[22]
port 121 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 req_addr_i[23]
port 122 nsew signal input
flabel metal3 s 89200 18368 90000 18488 0 FreeSans 480 0 0 0 req_addr_i[24]
port 123 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 req_addr_i[25]
port 124 nsew signal input
flabel metal2 s 36726 29200 36782 30000 0 FreeSans 224 90 0 0 req_addr_i[26]
port 125 nsew signal input
flabel metal2 s 28354 29200 28410 30000 0 FreeSans 224 90 0 0 req_addr_i[27]
port 126 nsew signal input
flabel metal2 s 16762 29200 16818 30000 0 FreeSans 224 90 0 0 req_addr_i[28]
port 127 nsew signal input
flabel metal2 s 82450 29200 82506 30000 0 FreeSans 224 90 0 0 req_addr_i[29]
port 128 nsew signal input
flabel metal2 s 63130 0 63186 800 0 FreeSans 224 90 0 0 req_addr_i[2]
port 129 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 req_addr_i[30]
port 130 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 req_addr_i[31]
port 131 nsew signal input
flabel metal2 s 1306 29200 1362 30000 0 FreeSans 224 90 0 0 req_addr_i[3]
port 132 nsew signal input
flabel metal2 s 89534 29200 89590 30000 0 FreeSans 224 90 0 0 req_addr_i[4]
port 133 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 req_addr_i[5]
port 134 nsew signal input
flabel metal2 s 85026 0 85082 800 0 FreeSans 224 90 0 0 req_addr_i[6]
port 135 nsew signal input
flabel metal2 s 23202 29200 23258 30000 0 FreeSans 224 90 0 0 req_addr_i[7]
port 136 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 req_addr_i[8]
port 137 nsew signal input
flabel metal2 s 67638 29200 67694 30000 0 FreeSans 224 90 0 0 req_addr_i[9]
port 138 nsew signal input
flabel metal3 s 89200 23128 90000 23248 0 FreeSans 480 0 0 0 req_ready_o
port 139 nsew signal tristate
flabel metal2 s 68282 29200 68338 30000 0 FreeSans 224 90 0 0 req_valid_i
port 140 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 resp_addr_o[0]
port 141 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 resp_addr_o[10]
port 142 nsew signal tristate
flabel metal2 s 21914 29200 21970 30000 0 FreeSans 224 90 0 0 resp_addr_o[11]
port 143 nsew signal tristate
flabel metal3 s 89200 21768 90000 21888 0 FreeSans 480 0 0 0 resp_addr_o[12]
port 144 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 resp_addr_o[13]
port 145 nsew signal tristate
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 resp_addr_o[14]
port 146 nsew signal tristate
flabel metal2 s 75366 29200 75422 30000 0 FreeSans 224 90 0 0 resp_addr_o[15]
port 147 nsew signal tristate
flabel metal2 s 79874 0 79930 800 0 FreeSans 224 90 0 0 resp_addr_o[16]
port 148 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 resp_addr_o[17]
port 149 nsew signal tristate
flabel metal2 s 56690 29200 56746 30000 0 FreeSans 224 90 0 0 resp_addr_o[18]
port 150 nsew signal tristate
flabel metal2 s 85670 29200 85726 30000 0 FreeSans 224 90 0 0 resp_addr_o[19]
port 151 nsew signal tristate
flabel metal2 s 81162 0 81218 800 0 FreeSans 224 90 0 0 resp_addr_o[1]
port 152 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 resp_addr_o[20]
port 153 nsew signal tristate
flabel metal2 s 48962 29200 49018 30000 0 FreeSans 224 90 0 0 resp_addr_o[21]
port 154 nsew signal tristate
flabel metal3 s 89200 16328 90000 16448 0 FreeSans 480 0 0 0 resp_addr_o[22]
port 155 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 resp_addr_o[23]
port 156 nsew signal tristate
flabel metal2 s 65706 29200 65762 30000 0 FreeSans 224 90 0 0 resp_addr_o[24]
port 157 nsew signal tristate
flabel metal2 s 60554 29200 60610 30000 0 FreeSans 224 90 0 0 resp_addr_o[25]
port 158 nsew signal tristate
flabel metal2 s 62486 0 62542 800 0 FreeSans 224 90 0 0 resp_addr_o[26]
port 159 nsew signal tristate
flabel metal2 s 56046 29200 56102 30000 0 FreeSans 224 90 0 0 resp_addr_o[27]
port 160 nsew signal tristate
flabel metal2 s 41234 29200 41290 30000 0 FreeSans 224 90 0 0 resp_addr_o[28]
port 161 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 resp_addr_o[29]
port 162 nsew signal tristate
flabel metal2 s 66994 0 67050 800 0 FreeSans 224 90 0 0 resp_addr_o[2]
port 163 nsew signal tristate
flabel metal2 s 84382 0 84438 800 0 FreeSans 224 90 0 0 resp_addr_o[30]
port 164 nsew signal tristate
flabel metal2 s 77298 0 77354 800 0 FreeSans 224 90 0 0 resp_addr_o[31]
port 165 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 resp_addr_o[3]
port 166 nsew signal tristate
flabel metal2 s 46386 29200 46442 30000 0 FreeSans 224 90 0 0 resp_addr_o[4]
port 167 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 resp_addr_o[5]
port 168 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 resp_addr_o[6]
port 169 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 resp_addr_o[7]
port 170 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 resp_addr_o[8]
port 171 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 resp_addr_o[9]
port 172 nsew signal tristate
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 resp_ready_i
port 173 nsew signal input
flabel metal2 s 76654 0 76710 800 0 FreeSans 224 90 0 0 resp_valid_o
port 174 nsew signal tristate
flabel metal3 s 89200 14968 90000 15088 0 FreeSans 480 0 0 0 rstn
port 175 nsew signal input
flabel metal2 s 43166 29200 43222 30000 0 FreeSans 224 90 0 0 tag_chip_en
port 176 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 tag_data_in[0]
port 177 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 tag_data_in[10]
port 178 nsew signal tristate
flabel metal2 s 81806 0 81862 800 0 FreeSans 224 90 0 0 tag_data_in[11]
port 179 nsew signal tristate
flabel metal2 s 34150 29200 34206 30000 0 FreeSans 224 90 0 0 tag_data_in[12]
port 180 nsew signal tristate
flabel metal2 s 14186 29200 14242 30000 0 FreeSans 224 90 0 0 tag_data_in[13]
port 181 nsew signal tristate
flabel metal2 s 2594 29200 2650 30000 0 FreeSans 224 90 0 0 tag_data_in[14]
port 182 nsew signal tristate
flabel metal2 s 77942 0 77998 800 0 FreeSans 224 90 0 0 tag_data_in[15]
port 183 nsew signal tristate
flabel metal3 s 89200 10208 90000 10328 0 FreeSans 480 0 0 0 tag_data_in[16]
port 184 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 tag_data_in[17]
port 185 nsew signal tristate
flabel metal2 s 32862 29200 32918 30000 0 FreeSans 224 90 0 0 tag_data_in[18]
port 186 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 tag_data_in[19]
port 187 nsew signal tristate
flabel metal3 s 89200 3408 90000 3528 0 FreeSans 480 0 0 0 tag_data_in[1]
port 188 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 tag_data_in[20]
port 189 nsew signal tristate
flabel metal3 s 89200 19728 90000 19848 0 FreeSans 480 0 0 0 tag_data_in[21]
port 190 nsew signal tristate
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 tag_data_in[22]
port 191 nsew signal tristate
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 tag_data_in[23]
port 192 nsew signal tristate
flabel metal2 s 64418 29200 64474 30000 0 FreeSans 224 90 0 0 tag_data_in[24]
port 193 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 tag_data_in[25]
port 194 nsew signal tristate
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 tag_data_in[26]
port 195 nsew signal tristate
flabel metal3 s 89200 17008 90000 17128 0 FreeSans 480 0 0 0 tag_data_in[27]
port 196 nsew signal tristate
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 tag_data_in[28]
port 197 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 tag_data_in[29]
port 198 nsew signal tristate
flabel metal2 s 18050 29200 18106 30000 0 FreeSans 224 90 0 0 tag_data_in[2]
port 199 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 tag_data_in[30]
port 200 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 tag_data_in[31]
port 201 nsew signal tristate
flabel metal3 s 89200 24488 90000 24608 0 FreeSans 480 0 0 0 tag_data_in[3]
port 202 nsew signal tristate
flabel metal2 s 24490 29200 24546 30000 0 FreeSans 224 90 0 0 tag_data_in[4]
port 203 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 tag_data_in[5]
port 204 nsew signal tristate
flabel metal2 s 3882 29200 3938 30000 0 FreeSans 224 90 0 0 tag_data_in[6]
port 205 nsew signal tristate
flabel metal2 s 78586 0 78642 800 0 FreeSans 224 90 0 0 tag_data_in[7]
port 206 nsew signal tristate
flabel metal2 s 38014 29200 38070 30000 0 FreeSans 224 90 0 0 tag_data_in[8]
port 207 nsew signal tristate
flabel metal2 s 57978 29200 58034 30000 0 FreeSans 224 90 0 0 tag_data_in[9]
port 208 nsew signal tristate
flabel metal2 s 66350 29200 66406 30000 0 FreeSans 224 90 0 0 tag_index[0]
port 209 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 tag_index[1]
port 210 nsew signal tristate
flabel metal2 s 86958 0 87014 800 0 FreeSans 224 90 0 0 tag_index[2]
port 211 nsew signal tristate
flabel metal2 s 18694 29200 18750 30000 0 FreeSans 224 90 0 0 tag_index[3]
port 212 nsew signal tristate
flabel metal2 s 52826 29200 52882 30000 0 FreeSans 224 90 0 0 tag_index[4]
port 213 nsew signal tristate
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 tag_index[5]
port 214 nsew signal tristate
flabel metal3 s 89200 23808 90000 23928 0 FreeSans 480 0 0 0 tag_index[6]
port 215 nsew signal tristate
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 tag_index[7]
port 216 nsew signal tristate
flabel metal2 s 79230 29200 79286 30000 0 FreeSans 224 90 0 0 tag_out[0]
port 217 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 tag_out[10]
port 218 nsew signal input
flabel metal2 s 30286 29200 30342 30000 0 FreeSans 224 90 0 0 tag_out[11]
port 219 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 tag_out[12]
port 220 nsew signal input
flabel metal2 s 80518 0 80574 800 0 FreeSans 224 90 0 0 tag_out[13]
port 221 nsew signal input
flabel metal2 s 31574 29200 31630 30000 0 FreeSans 224 90 0 0 tag_out[14]
port 222 nsew signal input
flabel metal2 s 88890 0 88946 800 0 FreeSans 224 90 0 0 tag_out[15]
port 223 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 tag_out[16]
port 224 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 tag_out[17]
port 225 nsew signal input
flabel metal2 s 61198 29200 61254 30000 0 FreeSans 224 90 0 0 tag_out[18]
port 226 nsew signal input
flabel metal3 s 89200 27208 90000 27328 0 FreeSans 480 0 0 0 tag_out[19]
port 227 nsew signal input
flabel metal2 s 10966 29200 11022 30000 0 FreeSans 224 90 0 0 tag_out[1]
port 228 nsew signal input
flabel metal2 s 58622 29200 58678 30000 0 FreeSans 224 90 0 0 tag_out[20]
port 229 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 tag_out[21]
port 230 nsew signal input
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 tag_out[22]
port 231 nsew signal input
flabel metal2 s 54758 29200 54814 30000 0 FreeSans 224 90 0 0 tag_out[23]
port 232 nsew signal input
flabel metal2 s 73434 0 73490 800 0 FreeSans 224 90 0 0 tag_out[24]
port 233 nsew signal input
flabel metal2 s 80518 29200 80574 30000 0 FreeSans 224 90 0 0 tag_out[25]
port 234 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 tag_out[26]
port 235 nsew signal input
flabel metal2 s 47030 29200 47086 30000 0 FreeSans 224 90 0 0 tag_out[27]
port 236 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 tag_out[28]
port 237 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 tag_out[29]
port 238 nsew signal input
flabel metal3 s 89200 5448 90000 5568 0 FreeSans 480 0 0 0 tag_out[2]
port 239 nsew signal input
flabel metal2 s 5814 29200 5870 30000 0 FreeSans 224 90 0 0 tag_out[30]
port 240 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 tag_out[31]
port 241 nsew signal input
flabel metal2 s 19338 29200 19394 30000 0 FreeSans 224 90 0 0 tag_out[3]
port 242 nsew signal input
flabel metal2 s 72146 0 72202 800 0 FreeSans 224 90 0 0 tag_out[4]
port 243 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 tag_out[5]
port 244 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 tag_out[6]
port 245 nsew signal input
flabel metal3 s 89200 25168 90000 25288 0 FreeSans 480 0 0 0 tag_out[7]
port 246 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 tag_out[8]
port 247 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 tag_out[9]
port 248 nsew signal input
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 tag_write_en
port 249 nsew signal tristate
flabel metal4 s 11918 2128 12238 27792 0 FreeSans 1920 90 0 0 vccd1
port 250 nsew power bidirectional
flabel metal4 s 33866 2128 34186 27792 0 FreeSans 1920 90 0 0 vccd1
port 250 nsew power bidirectional
flabel metal4 s 55814 2128 56134 27792 0 FreeSans 1920 90 0 0 vccd1
port 250 nsew power bidirectional
flabel metal4 s 77762 2128 78082 27792 0 FreeSans 1920 90 0 0 vccd1
port 250 nsew power bidirectional
flabel metal4 s 22892 2128 23212 27792 0 FreeSans 1920 90 0 0 vssd1
port 251 nsew ground bidirectional
flabel metal4 s 44840 2128 45160 27792 0 FreeSans 1920 90 0 0 vssd1
port 251 nsew ground bidirectional
flabel metal4 s 66788 2128 67108 27792 0 FreeSans 1920 90 0 0 vssd1
port 251 nsew ground bidirectional
flabel metal2 s 48318 29200 48374 30000 0 FreeSans 224 90 0 0 wb_ack_i
port 252 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 wb_adr_o[0]
port 253 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 wb_adr_o[10]
port 254 nsew signal tristate
flabel metal2 s 59910 29200 59966 30000 0 FreeSans 224 90 0 0 wb_adr_o[11]
port 255 nsew signal tristate
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 wb_adr_o[12]
port 256 nsew signal tristate
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 wb_adr_o[13]
port 257 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 wb_adr_o[14]
port 258 nsew signal tristate
flabel metal2 s 7746 29200 7802 30000 0 FreeSans 224 90 0 0 wb_adr_o[15]
port 259 nsew signal tristate
flabel metal2 s 79230 0 79286 800 0 FreeSans 224 90 0 0 wb_adr_o[16]
port 260 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 wb_adr_o[17]
port 261 nsew signal tristate
flabel metal2 s 83094 29200 83150 30000 0 FreeSans 224 90 0 0 wb_adr_o[18]
port 262 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 wb_adr_o[19]
port 263 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 wb_adr_o[1]
port 264 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wb_adr_o[20]
port 265 nsew signal tristate
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 wb_adr_o[21]
port 266 nsew signal tristate
flabel metal2 s 71502 0 71558 800 0 FreeSans 224 90 0 0 wb_adr_o[22]
port 267 nsew signal tristate
flabel metal2 s 57334 29200 57390 30000 0 FreeSans 224 90 0 0 wb_adr_o[23]
port 268 nsew signal tristate
flabel metal3 s 89200 15648 90000 15768 0 FreeSans 480 0 0 0 wb_adr_o[24]
port 269 nsew signal tristate
flabel metal2 s 26422 29200 26478 30000 0 FreeSans 224 90 0 0 wb_adr_o[25]
port 270 nsew signal tristate
flabel metal2 s 29642 29200 29698 30000 0 FreeSans 224 90 0 0 wb_adr_o[26]
port 271 nsew signal tristate
flabel metal2 s 27710 29200 27766 30000 0 FreeSans 224 90 0 0 wb_adr_o[27]
port 272 nsew signal tristate
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 wb_adr_o[28]
port 273 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 wb_adr_o[29]
port 274 nsew signal tristate
flabel metal2 s 86314 0 86370 800 0 FreeSans 224 90 0 0 wb_adr_o[2]
port 275 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 wb_adr_o[30]
port 276 nsew signal tristate
flabel metal2 s 76654 29200 76710 30000 0 FreeSans 224 90 0 0 wb_adr_o[31]
port 277 nsew signal tristate
flabel metal3 s 89200 29248 90000 29368 0 FreeSans 480 0 0 0 wb_adr_o[3]
port 278 nsew signal tristate
flabel metal2 s 40590 29200 40646 30000 0 FreeSans 224 90 0 0 wb_adr_o[4]
port 279 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wb_adr_o[5]
port 280 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 wb_adr_o[6]
port 281 nsew signal tristate
flabel metal3 s 89200 27888 90000 28008 0 FreeSans 480 0 0 0 wb_adr_o[7]
port 282 nsew signal tristate
flabel metal2 s 13542 29200 13598 30000 0 FreeSans 224 90 0 0 wb_adr_o[8]
port 283 nsew signal tristate
flabel metal3 s 89200 12248 90000 12368 0 FreeSans 480 0 0 0 wb_adr_o[9]
port 284 nsew signal tristate
flabel metal2 s 75366 0 75422 800 0 FreeSans 224 90 0 0 wb_bl_o[0]
port 285 nsew signal tristate
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 wb_bl_o[1]
port 286 nsew signal tristate
flabel metal2 s 84382 29200 84438 30000 0 FreeSans 224 90 0 0 wb_bl_o[2]
port 287 nsew signal tristate
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 wb_bl_o[3]
port 288 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wb_bl_o[4]
port 289 nsew signal tristate
flabel metal3 s 89200 2048 90000 2168 0 FreeSans 480 0 0 0 wb_bl_o[5]
port 290 nsew signal tristate
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 wb_bl_o[6]
port 291 nsew signal tristate
flabel metal2 s 74078 0 74134 800 0 FreeSans 224 90 0 0 wb_bl_o[7]
port 292 nsew signal tristate
flabel metal2 s 8390 29200 8446 30000 0 FreeSans 224 90 0 0 wb_bl_o[8]
port 293 nsew signal tristate
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 wb_bl_o[9]
port 294 nsew signal tristate
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wb_bry_o
port 295 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 wb_cyc_o
port 296 nsew signal tristate
flabel metal2 s 82450 0 82506 800 0 FreeSans 224 90 0 0 wb_dat_i[0]
port 297 nsew signal input
flabel metal2 s 81162 29200 81218 30000 0 FreeSans 224 90 0 0 wb_dat_i[10]
port 298 nsew signal input
flabel metal3 s 89200 20408 90000 20528 0 FreeSans 480 0 0 0 wb_dat_i[11]
port 299 nsew signal input
flabel metal2 s 61198 0 61254 800 0 FreeSans 224 90 0 0 wb_dat_i[12]
port 300 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 wb_dat_i[13]
port 301 nsew signal input
flabel metal3 s 89200 688 90000 808 0 FreeSans 480 0 0 0 wb_dat_i[14]
port 302 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 wb_dat_i[15]
port 303 nsew signal input
flabel metal3 s 89200 22448 90000 22568 0 FreeSans 480 0 0 0 wb_dat_i[16]
port 304 nsew signal input
flabel metal2 s 77942 29200 77998 30000 0 FreeSans 224 90 0 0 wb_dat_i[17]
port 305 nsew signal input
flabel metal2 s 64418 0 64474 800 0 FreeSans 224 90 0 0 wb_dat_i[18]
port 306 nsew signal input
flabel metal2 s 76010 29200 76066 30000 0 FreeSans 224 90 0 0 wb_dat_i[19]
port 307 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 wb_dat_i[1]
port 308 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 wb_dat_i[20]
port 309 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 wb_dat_i[21]
port 310 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 wb_dat_i[22]
port 311 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 wb_dat_i[23]
port 312 nsew signal input
flabel metal2 s 3238 29200 3294 30000 0 FreeSans 224 90 0 0 wb_dat_i[24]
port 313 nsew signal input
flabel metal2 s 25778 29200 25834 30000 0 FreeSans 224 90 0 0 wb_dat_i[25]
port 314 nsew signal input
flabel metal2 s 49606 29200 49662 30000 0 FreeSans 224 90 0 0 wb_dat_i[26]
port 315 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 wb_dat_i[27]
port 316 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wb_dat_i[28]
port 317 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 wb_dat_i[29]
port 318 nsew signal input
flabel metal2 s 63774 29200 63830 30000 0 FreeSans 224 90 0 0 wb_dat_i[2]
port 319 nsew signal input
flabel metal2 s 50250 29200 50306 30000 0 FreeSans 224 90 0 0 wb_dat_i[30]
port 320 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 wb_dat_i[31]
port 321 nsew signal input
flabel metal2 s 73434 29200 73490 30000 0 FreeSans 224 90 0 0 wb_dat_i[3]
port 322 nsew signal input
flabel metal2 s 74722 0 74778 800 0 FreeSans 224 90 0 0 wb_dat_i[4]
port 323 nsew signal input
flabel metal2 s 12254 29200 12310 30000 0 FreeSans 224 90 0 0 wb_dat_i[5]
port 324 nsew signal input
flabel metal3 s 89200 14288 90000 14408 0 FreeSans 480 0 0 0 wb_dat_i[6]
port 325 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wb_dat_i[7]
port 326 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wb_dat_i[8]
port 327 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 wb_dat_i[9]
port 328 nsew signal input
flabel metal3 s 89200 12928 90000 13048 0 FreeSans 480 0 0 0 wb_stb_o
port 329 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 wb_we_o
port 330 nsew signal tristate
flabel metal2 s 70214 29200 70270 30000 0 FreeSans 224 90 0 0 write_data_mask[0]
port 331 nsew signal tristate
flabel metal2 s 68926 29200 68982 30000 0 FreeSans 224 90 0 0 write_data_mask[1]
port 332 nsew signal tristate
flabel metal2 s 27066 29200 27122 30000 0 FreeSans 224 90 0 0 write_data_mask[2]
port 333 nsew signal tristate
flabel metal2 s 37370 29200 37426 30000 0 FreeSans 224 90 0 0 write_data_mask[3]
port 334 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 write_tag_mask[0]
port 335 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 write_tag_mask[1]
port 336 nsew signal tristate
flabel metal2 s 20626 29200 20682 30000 0 FreeSans 224 90 0 0 write_tag_mask[2]
port 337 nsew signal tristate
flabel metal2 s 88246 0 88302 800 0 FreeSans 224 90 0 0 write_tag_mask[3]
port 338 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 90000 30000
<< end >>
