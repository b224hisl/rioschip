VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bus_arbiter
  CLASS BLOCK ;
  FOREIGN bus_arbiter ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 150.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 44.240 600.000 44.840 ;
    END
  END clk
  PIN m2_dcache_wbd_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 146.000 93.750 150.000 ;
    END
  END m2_dcache_wbd_ack_o
  PIN m2_dcache_wbd_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 146.000 373.890 150.000 ;
    END
  END m2_dcache_wbd_adr_i[0]
  PIN m2_dcache_wbd_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 146.000 32.570 150.000 ;
    END
  END m2_dcache_wbd_adr_i[10]
  PIN m2_dcache_wbd_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END m2_dcache_wbd_adr_i[11]
  PIN m2_dcache_wbd_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 146.000 196.790 150.000 ;
    END
  END m2_dcache_wbd_adr_i[12]
  PIN m2_dcache_wbd_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 146.000 219.330 150.000 ;
    END
  END m2_dcache_wbd_adr_i[13]
  PIN m2_dcache_wbd_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 146.000 55.110 150.000 ;
    END
  END m2_dcache_wbd_adr_i[14]
  PIN m2_dcache_wbd_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 146.000 142.050 150.000 ;
    END
  END m2_dcache_wbd_adr_i[15]
  PIN m2_dcache_wbd_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 146.000 167.810 150.000 ;
    END
  END m2_dcache_wbd_adr_i[16]
  PIN m2_dcache_wbd_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 81.640 600.000 82.240 ;
    END
  END m2_dcache_wbd_adr_i[17]
  PIN m2_dcache_wbd_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END m2_dcache_wbd_adr_i[18]
  PIN m2_dcache_wbd_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 146.000 332.030 150.000 ;
    END
  END m2_dcache_wbd_adr_i[19]
  PIN m2_dcache_wbd_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END m2_dcache_wbd_adr_i[1]
  PIN m2_dcache_wbd_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END m2_dcache_wbd_adr_i[20]
  PIN m2_dcache_wbd_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 115.640 600.000 116.240 ;
    END
  END m2_dcache_wbd_adr_i[21]
  PIN m2_dcache_wbd_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END m2_dcache_wbd_adr_i[22]
  PIN m2_dcache_wbd_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END m2_dcache_wbd_adr_i[23]
  PIN m2_dcache_wbd_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END m2_dcache_wbd_adr_i[24]
  PIN m2_dcache_wbd_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 146.000 512.350 150.000 ;
    END
  END m2_dcache_wbd_adr_i[25]
  PIN m2_dcache_wbd_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 146.000 296.610 150.000 ;
    END
  END m2_dcache_wbd_adr_i[26]
  PIN m2_dcache_wbd_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END m2_dcache_wbd_adr_i[27]
  PIN m2_dcache_wbd_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END m2_dcache_wbd_adr_i[28]
  PIN m2_dcache_wbd_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END m2_dcache_wbd_adr_i[29]
  PIN m2_dcache_wbd_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 146.000 579.970 150.000 ;
    END
  END m2_dcache_wbd_adr_i[2]
  PIN m2_dcache_wbd_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END m2_dcache_wbd_adr_i[30]
  PIN m2_dcache_wbd_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END m2_dcache_wbd_adr_i[31]
  PIN m2_dcache_wbd_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END m2_dcache_wbd_adr_i[3]
  PIN m2_dcache_wbd_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 10.240 600.000 10.840 ;
    END
  END m2_dcache_wbd_adr_i[4]
  PIN m2_dcache_wbd_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 146.000 174.250 150.000 ;
    END
  END m2_dcache_wbd_adr_i[5]
  PIN m2_dcache_wbd_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 146.000 119.510 150.000 ;
    END
  END m2_dcache_wbd_adr_i[6]
  PIN m2_dcache_wbd_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 20.440 600.000 21.040 ;
    END
  END m2_dcache_wbd_adr_i[7]
  PIN m2_dcache_wbd_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END m2_dcache_wbd_adr_i[8]
  PIN m2_dcache_wbd_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 146.000 13.250 150.000 ;
    END
  END m2_dcache_wbd_adr_i[9]
  PIN m2_dcache_wbd_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END m2_dcache_wbd_cyc_i
  PIN m2_dcache_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 105.440 600.000 106.040 ;
    END
  END m2_dcache_wbd_dat_i[0]
  PIN m2_dcache_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 146.000 364.230 150.000 ;
    END
  END m2_dcache_wbd_dat_i[10]
  PIN m2_dcache_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 146.000 328.810 150.000 ;
    END
  END m2_dcache_wbd_dat_i[11]
  PIN m2_dcache_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 146.000 341.690 150.000 ;
    END
  END m2_dcache_wbd_dat_i[12]
  PIN m2_dcache_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 146.000 187.130 150.000 ;
    END
  END m2_dcache_wbd_dat_i[13]
  PIN m2_dcache_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END m2_dcache_wbd_dat_i[14]
  PIN m2_dcache_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END m2_dcache_wbd_dat_i[15]
  PIN m2_dcache_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 146.000 145.270 150.000 ;
    END
  END m2_dcache_wbd_dat_i[16]
  PIN m2_dcache_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END m2_dcache_wbd_dat_i[17]
  PIN m2_dcache_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 146.000 267.630 150.000 ;
    END
  END m2_dcache_wbd_dat_i[18]
  PIN m2_dcache_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 146.000 45.450 150.000 ;
    END
  END m2_dcache_wbd_dat_i[19]
  PIN m2_dcache_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END m2_dcache_wbd_dat_i[1]
  PIN m2_dcache_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 146.000 26.130 150.000 ;
    END
  END m2_dcache_wbd_dat_i[20]
  PIN m2_dcache_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 146.000 67.990 150.000 ;
    END
  END m2_dcache_wbd_dat_i[21]
  PIN m2_dcache_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END m2_dcache_wbd_dat_i[22]
  PIN m2_dcache_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END m2_dcache_wbd_dat_i[23]
  PIN m2_dcache_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END m2_dcache_wbd_dat_i[24]
  PIN m2_dcache_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 146.000 77.650 150.000 ;
    END
  END m2_dcache_wbd_dat_i[25]
  PIN m2_dcache_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END m2_dcache_wbd_dat_i[26]
  PIN m2_dcache_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END m2_dcache_wbd_dat_i[27]
  PIN m2_dcache_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 146.000 393.210 150.000 ;
    END
  END m2_dcache_wbd_dat_i[28]
  PIN m2_dcache_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 146.000 135.610 150.000 ;
    END
  END m2_dcache_wbd_dat_i[29]
  PIN m2_dcache_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 146.000 354.570 150.000 ;
    END
  END m2_dcache_wbd_dat_i[2]
  PIN m2_dcache_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 146.000 428.630 150.000 ;
    END
  END m2_dcache_wbd_dat_i[30]
  PIN m2_dcache_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END m2_dcache_wbd_dat_i[31]
  PIN m2_dcache_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 146.000 315.930 150.000 ;
    END
  END m2_dcache_wbd_dat_i[3]
  PIN m2_dcache_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END m2_dcache_wbd_dat_i[4]
  PIN m2_dcache_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 146.000 80.870 150.000 ;
    END
  END m2_dcache_wbd_dat_i[5]
  PIN m2_dcache_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END m2_dcache_wbd_dat_i[6]
  PIN m2_dcache_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END m2_dcache_wbd_dat_i[7]
  PIN m2_dcache_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 146.000 534.890 150.000 ;
    END
  END m2_dcache_wbd_dat_i[8]
  PIN m2_dcache_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 13.640 600.000 14.240 ;
    END
  END m2_dcache_wbd_dat_i[9]
  PIN m2_dcache_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END m2_dcache_wbd_dat_o[0]
  PIN m2_dcache_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END m2_dcache_wbd_dat_o[10]
  PIN m2_dcache_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END m2_dcache_wbd_dat_o[11]
  PIN m2_dcache_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 146.000 39.010 150.000 ;
    END
  END m2_dcache_wbd_dat_o[12]
  PIN m2_dcache_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 146.000 286.950 150.000 ;
    END
  END m2_dcache_wbd_dat_o[13]
  PIN m2_dcache_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 146.000 212.890 150.000 ;
    END
  END m2_dcache_wbd_dat_o[14]
  PIN m2_dcache_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 146.000 522.010 150.000 ;
    END
  END m2_dcache_wbd_dat_o[15]
  PIN m2_dcache_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 146.000 406.090 150.000 ;
    END
  END m2_dcache_wbd_dat_o[16]
  PIN m2_dcache_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END m2_dcache_wbd_dat_o[17]
  PIN m2_dcache_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 146.000 177.470 150.000 ;
    END
  END m2_dcache_wbd_dat_o[18]
  PIN m2_dcache_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END m2_dcache_wbd_dat_o[19]
  PIN m2_dcache_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END m2_dcache_wbd_dat_o[1]
  PIN m2_dcache_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END m2_dcache_wbd_dat_o[20]
  PIN m2_dcache_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 146.000 544.550 150.000 ;
    END
  END m2_dcache_wbd_dat_o[21]
  PIN m2_dcache_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 146.000 228.990 150.000 ;
    END
  END m2_dcache_wbd_dat_o[22]
  PIN m2_dcache_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END m2_dcache_wbd_dat_o[23]
  PIN m2_dcache_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END m2_dcache_wbd_dat_o[24]
  PIN m2_dcache_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 146.000 48.670 150.000 ;
    END
  END m2_dcache_wbd_dat_o[25]
  PIN m2_dcache_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 146.000 467.270 150.000 ;
    END
  END m2_dcache_wbd_dat_o[26]
  PIN m2_dcache_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END m2_dcache_wbd_dat_o[27]
  PIN m2_dcache_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 146.000 190.350 150.000 ;
    END
  END m2_dcache_wbd_dat_o[28]
  PIN m2_dcache_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 146.000 412.530 150.000 ;
    END
  END m2_dcache_wbd_dat_o[29]
  PIN m2_dcache_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END m2_dcache_wbd_dat_o[2]
  PIN m2_dcache_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END m2_dcache_wbd_dat_o[30]
  PIN m2_dcache_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END m2_dcache_wbd_dat_o[31]
  PIN m2_dcache_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END m2_dcache_wbd_dat_o[3]
  PIN m2_dcache_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END m2_dcache_wbd_dat_o[4]
  PIN m2_dcache_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 146.000 338.470 150.000 ;
    END
  END m2_dcache_wbd_dat_o[5]
  PIN m2_dcache_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 125.840 600.000 126.440 ;
    END
  END m2_dcache_wbd_dat_o[6]
  PIN m2_dcache_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 146.000 264.410 150.000 ;
    END
  END m2_dcache_wbd_dat_o[7]
  PIN m2_dcache_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END m2_dcache_wbd_dat_o[8]
  PIN m2_dcache_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END m2_dcache_wbd_dat_o[9]
  PIN m2_dcache_wbd_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END m2_dcache_wbd_sel_i[0]
  PIN m2_dcache_wbd_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END m2_dcache_wbd_sel_i[1]
  PIN m2_dcache_wbd_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 146.000 589.630 150.000 ;
    END
  END m2_dcache_wbd_sel_i[2]
  PIN m2_dcache_wbd_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END m2_dcache_wbd_sel_i[3]
  PIN m2_dcache_wbd_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 139.440 600.000 140.040 ;
    END
  END m2_dcache_wbd_stb_i
  PIN m2_dcache_wbd_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END m2_dcache_wbd_we_i
  PIN m2_others_wbd_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END m2_others_wbd_ack_o
  PIN m2_others_wbd_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 146.000 245.090 150.000 ;
    END
  END m2_others_wbd_adr_i[0]
  PIN m2_others_wbd_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END m2_others_wbd_adr_i[10]
  PIN m2_others_wbd_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END m2_others_wbd_adr_i[11]
  PIN m2_others_wbd_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END m2_others_wbd_adr_i[12]
  PIN m2_others_wbd_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 71.440 600.000 72.040 ;
    END
  END m2_others_wbd_adr_i[13]
  PIN m2_others_wbd_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 146.000 319.150 150.000 ;
    END
  END m2_others_wbd_adr_i[14]
  PIN m2_others_wbd_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END m2_others_wbd_adr_i[15]
  PIN m2_others_wbd_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END m2_others_wbd_adr_i[16]
  PIN m2_others_wbd_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END m2_others_wbd_adr_i[17]
  PIN m2_others_wbd_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 146.000 154.930 150.000 ;
    END
  END m2_others_wbd_adr_i[18]
  PIN m2_others_wbd_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END m2_others_wbd_adr_i[19]
  PIN m2_others_wbd_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 146.000 61.550 150.000 ;
    END
  END m2_others_wbd_adr_i[1]
  PIN m2_others_wbd_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END m2_others_wbd_adr_i[20]
  PIN m2_others_wbd_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 146.000 180.690 150.000 ;
    END
  END m2_others_wbd_adr_i[21]
  PIN m2_others_wbd_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END m2_others_wbd_adr_i[22]
  PIN m2_others_wbd_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END m2_others_wbd_adr_i[23]
  PIN m2_others_wbd_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 30.640 600.000 31.240 ;
    END
  END m2_others_wbd_adr_i[24]
  PIN m2_others_wbd_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 146.000 415.750 150.000 ;
    END
  END m2_others_wbd_adr_i[25]
  PIN m2_others_wbd_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END m2_others_wbd_adr_i[26]
  PIN m2_others_wbd_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 146.000 87.310 150.000 ;
    END
  END m2_others_wbd_adr_i[27]
  PIN m2_others_wbd_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END m2_others_wbd_adr_i[28]
  PIN m2_others_wbd_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END m2_others_wbd_adr_i[29]
  PIN m2_others_wbd_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 146.000 158.150 150.000 ;
    END
  END m2_others_wbd_adr_i[2]
  PIN m2_others_wbd_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 146.000 322.370 150.000 ;
    END
  END m2_others_wbd_adr_i[30]
  PIN m2_others_wbd_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 146.000 441.510 150.000 ;
    END
  END m2_others_wbd_adr_i[31]
  PIN m2_others_wbd_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 146.000 261.190 150.000 ;
    END
  END m2_others_wbd_adr_i[3]
  PIN m2_others_wbd_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 68.040 600.000 68.640 ;
    END
  END m2_others_wbd_adr_i[4]
  PIN m2_others_wbd_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END m2_others_wbd_adr_i[5]
  PIN m2_others_wbd_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END m2_others_wbd_adr_i[6]
  PIN m2_others_wbd_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END m2_others_wbd_adr_i[7]
  PIN m2_others_wbd_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 146.000 457.610 150.000 ;
    END
  END m2_others_wbd_adr_i[8]
  PIN m2_others_wbd_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END m2_others_wbd_adr_i[9]
  PIN m2_others_wbd_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END m2_others_wbd_cyc_i
  PIN m2_others_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 146.000 592.850 150.000 ;
    END
  END m2_others_wbd_dat_i[0]
  PIN m2_others_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END m2_others_wbd_dat_i[10]
  PIN m2_others_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 146.000 380.330 150.000 ;
    END
  END m2_others_wbd_dat_i[11]
  PIN m2_others_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 146.240 600.000 146.840 ;
    END
  END m2_others_wbd_dat_i[12]
  PIN m2_others_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 146.000 599.290 150.000 ;
    END
  END m2_others_wbd_dat_i[13]
  PIN m2_others_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END m2_others_wbd_dat_i[14]
  PIN m2_others_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 146.000 447.950 150.000 ;
    END
  END m2_others_wbd_dat_i[15]
  PIN m2_others_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 146.000 370.670 150.000 ;
    END
  END m2_others_wbd_dat_i[16]
  PIN m2_others_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 146.000 35.790 150.000 ;
    END
  END m2_others_wbd_dat_i[17]
  PIN m2_others_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 0.040 600.000 0.640 ;
    END
  END m2_others_wbd_dat_i[18]
  PIN m2_others_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 146.000 383.550 150.000 ;
    END
  END m2_others_wbd_dat_i[19]
  PIN m2_others_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END m2_others_wbd_dat_i[1]
  PIN m2_others_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 146.000 6.810 150.000 ;
    END
  END m2_others_wbd_dat_i[20]
  PIN m2_others_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END m2_others_wbd_dat_i[21]
  PIN m2_others_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 146.000 71.210 150.000 ;
    END
  END m2_others_wbd_dat_i[22]
  PIN m2_others_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END m2_others_wbd_dat_i[23]
  PIN m2_others_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 146.000 560.650 150.000 ;
    END
  END m2_others_wbd_dat_i[24]
  PIN m2_others_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END m2_others_wbd_dat_i[25]
  PIN m2_others_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END m2_others_wbd_dat_i[26]
  PIN m2_others_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END m2_others_wbd_dat_i[27]
  PIN m2_others_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END m2_others_wbd_dat_i[28]
  PIN m2_others_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END m2_others_wbd_dat_i[29]
  PIN m2_others_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 146.000 505.910 150.000 ;
    END
  END m2_others_wbd_dat_i[2]
  PIN m2_others_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END m2_others_wbd_dat_i[30]
  PIN m2_others_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 146.000 109.850 150.000 ;
    END
  END m2_others_wbd_dat_i[31]
  PIN m2_others_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 146.000 493.030 150.000 ;
    END
  END m2_others_wbd_dat_i[3]
  PIN m2_others_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 91.840 600.000 92.440 ;
    END
  END m2_others_wbd_dat_i[4]
  PIN m2_others_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END m2_others_wbd_dat_i[5]
  PIN m2_others_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 146.000 241.870 150.000 ;
    END
  END m2_others_wbd_dat_i[6]
  PIN m2_others_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END m2_others_wbd_dat_i[7]
  PIN m2_others_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 146.000 90.530 150.000 ;
    END
  END m2_others_wbd_dat_i[8]
  PIN m2_others_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 146.000 125.950 150.000 ;
    END
  END m2_others_wbd_dat_i[9]
  PIN m2_others_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 146.000 103.410 150.000 ;
    END
  END m2_others_wbd_dat_o[0]
  PIN m2_others_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 6.840 600.000 7.440 ;
    END
  END m2_others_wbd_dat_o[10]
  PIN m2_others_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 23.840 600.000 24.440 ;
    END
  END m2_others_wbd_dat_o[11]
  PIN m2_others_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END m2_others_wbd_dat_o[12]
  PIN m2_others_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 146.000 277.290 150.000 ;
    END
  END m2_others_wbd_dat_o[13]
  PIN m2_others_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END m2_others_wbd_dat_o[14]
  PIN m2_others_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END m2_others_wbd_dat_o[15]
  PIN m2_others_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 64.640 600.000 65.240 ;
    END
  END m2_others_wbd_dat_o[16]
  PIN m2_others_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 146.000 489.810 150.000 ;
    END
  END m2_others_wbd_dat_o[17]
  PIN m2_others_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END m2_others_wbd_dat_o[18]
  PIN m2_others_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 146.000 460.830 150.000 ;
    END
  END m2_others_wbd_dat_o[19]
  PIN m2_others_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END m2_others_wbd_dat_o[1]
  PIN m2_others_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 146.000 283.730 150.000 ;
    END
  END m2_others_wbd_dat_o[20]
  PIN m2_others_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 47.640 600.000 48.240 ;
    END
  END m2_others_wbd_dat_o[21]
  PIN m2_others_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END m2_others_wbd_dat_o[22]
  PIN m2_others_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 146.000 502.690 150.000 ;
    END
  END m2_others_wbd_dat_o[23]
  PIN m2_others_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 146.000 22.910 150.000 ;
    END
  END m2_others_wbd_dat_o[24]
  PIN m2_others_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END m2_others_wbd_dat_o[25]
  PIN m2_others_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END m2_others_wbd_dat_o[26]
  PIN m2_others_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 102.040 600.000 102.640 ;
    END
  END m2_others_wbd_dat_o[27]
  PIN m2_others_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END m2_others_wbd_dat_o[28]
  PIN m2_others_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END m2_others_wbd_dat_o[29]
  PIN m2_others_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END m2_others_wbd_dat_o[2]
  PIN m2_others_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END m2_others_wbd_dat_o[30]
  PIN m2_others_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 146.000 148.490 150.000 ;
    END
  END m2_others_wbd_dat_o[31]
  PIN m2_others_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 146.000 254.750 150.000 ;
    END
  END m2_others_wbd_dat_o[3]
  PIN m2_others_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 146.000 470.490 150.000 ;
    END
  END m2_others_wbd_dat_o[4]
  PIN m2_others_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END m2_others_wbd_dat_o[5]
  PIN m2_others_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END m2_others_wbd_dat_o[6]
  PIN m2_others_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 146.000 586.410 150.000 ;
    END
  END m2_others_wbd_dat_o[7]
  PIN m2_others_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 146.000 386.770 150.000 ;
    END
  END m2_others_wbd_dat_o[8]
  PIN m2_others_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END m2_others_wbd_dat_o[9]
  PIN m2_others_wbd_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 146.000 16.470 150.000 ;
    END
  END m2_others_wbd_sel_i[0]
  PIN m2_others_wbd_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END m2_others_wbd_sel_i[1]
  PIN m2_others_wbd_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 146.000 554.210 150.000 ;
    END
  END m2_others_wbd_sel_i[2]
  PIN m2_others_wbd_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END m2_others_wbd_sel_i[3]
  PIN m2_others_wbd_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END m2_others_wbd_stb_i
  PIN m2_others_wbd_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END m2_others_wbd_we_i
  PIN m2_wbd_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END m2_wbd_ack_i
  PIN m2_wbd_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 146.000 309.490 150.000 ;
    END
  END m2_wbd_adr_o[0]
  PIN m2_wbd_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 146.000 293.390 150.000 ;
    END
  END m2_wbd_adr_o[10]
  PIN m2_wbd_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END m2_wbd_adr_o[11]
  PIN m2_wbd_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END m2_wbd_adr_o[12]
  PIN m2_wbd_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 146.000 438.290 150.000 ;
    END
  END m2_wbd_adr_o[13]
  PIN m2_wbd_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 122.440 600.000 123.040 ;
    END
  END m2_wbd_adr_o[14]
  PIN m2_wbd_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 146.000 306.270 150.000 ;
    END
  END m2_wbd_adr_o[15]
  PIN m2_wbd_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 146.000 418.970 150.000 ;
    END
  END m2_wbd_adr_o[16]
  PIN m2_wbd_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 146.000 451.170 150.000 ;
    END
  END m2_wbd_adr_o[17]
  PIN m2_wbd_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END m2_wbd_adr_o[18]
  PIN m2_wbd_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 146.000 396.430 150.000 ;
    END
  END m2_wbd_adr_o[19]
  PIN m2_wbd_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END m2_wbd_adr_o[1]
  PIN m2_wbd_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 146.000 557.430 150.000 ;
    END
  END m2_wbd_adr_o[20]
  PIN m2_wbd_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 146.000 483.370 150.000 ;
    END
  END m2_wbd_adr_o[21]
  PIN m2_wbd_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END m2_wbd_adr_o[22]
  PIN m2_wbd_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END m2_wbd_adr_o[23]
  PIN m2_wbd_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 146.000 251.530 150.000 ;
    END
  END m2_wbd_adr_o[24]
  PIN m2_wbd_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END m2_wbd_adr_o[25]
  PIN m2_wbd_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 146.000 122.730 150.000 ;
    END
  END m2_wbd_adr_o[26]
  PIN m2_wbd_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END m2_wbd_adr_o[27]
  PIN m2_wbd_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 146.000 235.430 150.000 ;
    END
  END m2_wbd_adr_o[28]
  PIN m2_wbd_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END m2_wbd_adr_o[29]
  PIN m2_wbd_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END m2_wbd_adr_o[2]
  PIN m2_wbd_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 146.000 538.110 150.000 ;
    END
  END m2_wbd_adr_o[30]
  PIN m2_wbd_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 112.240 600.000 112.840 ;
    END
  END m2_wbd_adr_o[31]
  PIN m2_wbd_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END m2_wbd_adr_o[3]
  PIN m2_wbd_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END m2_wbd_adr_o[4]
  PIN m2_wbd_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END m2_wbd_adr_o[5]
  PIN m2_wbd_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END m2_wbd_adr_o[6]
  PIN m2_wbd_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END m2_wbd_adr_o[7]
  PIN m2_wbd_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END m2_wbd_adr_o[8]
  PIN m2_wbd_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 146.000 425.410 150.000 ;
    END
  END m2_wbd_adr_o[9]
  PIN m2_wbd_bl_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END m2_wbd_bl_o[0]
  PIN m2_wbd_bl_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 78.240 600.000 78.840 ;
    END
  END m2_wbd_bl_o[1]
  PIN m2_wbd_bl_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END m2_wbd_bl_o[2]
  PIN m2_wbd_bl_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 146.000 576.750 150.000 ;
    END
  END m2_wbd_bl_o[3]
  PIN m2_wbd_bl_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END m2_wbd_bl_o[4]
  PIN m2_wbd_bl_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END m2_wbd_bl_o[5]
  PIN m2_wbd_bl_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 146.000 567.090 150.000 ;
    END
  END m2_wbd_bl_o[6]
  PIN m2_wbd_bl_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END m2_wbd_bl_o[7]
  PIN m2_wbd_bl_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END m2_wbd_bl_o[8]
  PIN m2_wbd_bl_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END m2_wbd_bl_o[9]
  PIN m2_wbd_bry_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END m2_wbd_bry_o
  PIN m2_wbd_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END m2_wbd_cyc_o
  PIN m2_wbd_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 146.000 402.870 150.000 ;
    END
  END m2_wbd_dat_i[0]
  PIN m2_wbd_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 57.840 600.000 58.440 ;
    END
  END m2_wbd_dat_i[10]
  PIN m2_wbd_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 146.000 209.670 150.000 ;
    END
  END m2_wbd_dat_i[11]
  PIN m2_wbd_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 146.000 232.210 150.000 ;
    END
  END m2_wbd_dat_i[12]
  PIN m2_wbd_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 146.000 222.550 150.000 ;
    END
  END m2_wbd_dat_i[13]
  PIN m2_wbd_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END m2_wbd_dat_i[14]
  PIN m2_wbd_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END m2_wbd_dat_i[15]
  PIN m2_wbd_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END m2_wbd_dat_i[16]
  PIN m2_wbd_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END m2_wbd_dat_i[17]
  PIN m2_wbd_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 146.000 525.230 150.000 ;
    END
  END m2_wbd_dat_i[18]
  PIN m2_wbd_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 136.040 600.000 136.640 ;
    END
  END m2_wbd_dat_i[19]
  PIN m2_wbd_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 146.000 299.830 150.000 ;
    END
  END m2_wbd_dat_i[1]
  PIN m2_wbd_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END m2_wbd_dat_i[20]
  PIN m2_wbd_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END m2_wbd_dat_i[21]
  PIN m2_wbd_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 132.640 600.000 133.240 ;
    END
  END m2_wbd_dat_i[22]
  PIN m2_wbd_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 146.000 132.390 150.000 ;
    END
  END m2_wbd_dat_i[23]
  PIN m2_wbd_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 34.040 600.000 34.640 ;
    END
  END m2_wbd_dat_i[24]
  PIN m2_wbd_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END m2_wbd_dat_i[25]
  PIN m2_wbd_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 146.000 0.370 150.000 ;
    END
  END m2_wbd_dat_i[26]
  PIN m2_wbd_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 146.000 570.310 150.000 ;
    END
  END m2_wbd_dat_i[27]
  PIN m2_wbd_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 146.000 361.010 150.000 ;
    END
  END m2_wbd_dat_i[28]
  PIN m2_wbd_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END m2_wbd_dat_i[29]
  PIN m2_wbd_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END m2_wbd_dat_i[2]
  PIN m2_wbd_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END m2_wbd_dat_i[30]
  PIN m2_wbd_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END m2_wbd_dat_i[31]
  PIN m2_wbd_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 146.000 100.190 150.000 ;
    END
  END m2_wbd_dat_i[3]
  PIN m2_wbd_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END m2_wbd_dat_i[4]
  PIN m2_wbd_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END m2_wbd_dat_i[5]
  PIN m2_wbd_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END m2_wbd_dat_i[6]
  PIN m2_wbd_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END m2_wbd_dat_i[7]
  PIN m2_wbd_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 146.000 547.770 150.000 ;
    END
  END m2_wbd_dat_i[8]
  PIN m2_wbd_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 88.440 600.000 89.040 ;
    END
  END m2_wbd_dat_i[9]
  PIN m2_wbd_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END m2_wbd_dat_o[0]
  PIN m2_wbd_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END m2_wbd_dat_o[10]
  PIN m2_wbd_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END m2_wbd_dat_o[11]
  PIN m2_wbd_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END m2_wbd_dat_o[12]
  PIN m2_wbd_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 98.640 600.000 99.240 ;
    END
  END m2_wbd_dat_o[13]
  PIN m2_wbd_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 146.000 528.450 150.000 ;
    END
  END m2_wbd_dat_o[14]
  PIN m2_wbd_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END m2_wbd_dat_o[15]
  PIN m2_wbd_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 146.000 515.570 150.000 ;
    END
  END m2_wbd_dat_o[16]
  PIN m2_wbd_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END m2_wbd_dat_o[17]
  PIN m2_wbd_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END m2_wbd_dat_o[18]
  PIN m2_wbd_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END m2_wbd_dat_o[19]
  PIN m2_wbd_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END m2_wbd_dat_o[1]
  PIN m2_wbd_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END m2_wbd_dat_o[20]
  PIN m2_wbd_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 146.000 58.330 150.000 ;
    END
  END m2_wbd_dat_o[21]
  PIN m2_wbd_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 146.000 200.010 150.000 ;
    END
  END m2_wbd_dat_o[22]
  PIN m2_wbd_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 146.000 348.130 150.000 ;
    END
  END m2_wbd_dat_o[23]
  PIN m2_wbd_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 146.000 3.590 150.000 ;
    END
  END m2_wbd_dat_o[24]
  PIN m2_wbd_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END m2_wbd_dat_o[25]
  PIN m2_wbd_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END m2_wbd_dat_o[26]
  PIN m2_wbd_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 146.000 435.070 150.000 ;
    END
  END m2_wbd_dat_o[27]
  PIN m2_wbd_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 146.000 351.350 150.000 ;
    END
  END m2_wbd_dat_o[28]
  PIN m2_wbd_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END m2_wbd_dat_o[29]
  PIN m2_wbd_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 146.000 499.470 150.000 ;
    END
  END m2_wbd_dat_o[2]
  PIN m2_wbd_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END m2_wbd_dat_o[30]
  PIN m2_wbd_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 146.000 113.070 150.000 ;
    END
  END m2_wbd_dat_o[31]
  PIN m2_wbd_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 54.440 600.000 55.040 ;
    END
  END m2_wbd_dat_o[3]
  PIN m2_wbd_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END m2_wbd_dat_o[4]
  PIN m2_wbd_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END m2_wbd_dat_o[5]
  PIN m2_wbd_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END m2_wbd_dat_o[6]
  PIN m2_wbd_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 40.840 600.000 41.440 ;
    END
  END m2_wbd_dat_o[7]
  PIN m2_wbd_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END m2_wbd_dat_o[8]
  PIN m2_wbd_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 146.000 480.150 150.000 ;
    END
  END m2_wbd_dat_o[9]
  PIN m2_wbd_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 146.000 473.710 150.000 ;
    END
  END m2_wbd_sel_o[0]
  PIN m2_wbd_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 146.000 206.450 150.000 ;
    END
  END m2_wbd_sel_o[1]
  PIN m2_wbd_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 146.000 274.070 150.000 ;
    END
  END m2_wbd_sel_o[2]
  PIN m2_wbd_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END m2_wbd_sel_o[3]
  PIN m2_wbd_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END m2_wbd_stb_o
  PIN m2_wbd_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 146.000 164.590 150.000 ;
    END
  END m2_wbd_we_o
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 78.340 10.640 79.940 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.580 10.640 227.180 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 372.820 10.640 374.420 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 520.060 10.640 521.660 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 151.960 10.640 153.560 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 299.200 10.640 300.800 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.440 10.640 448.040 138.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 138.805 ;
      LAYER met1 ;
        RECT 0.070 5.480 599.310 140.720 ;
      LAYER met2 ;
        RECT 0.650 145.720 3.030 146.610 ;
        RECT 3.870 145.720 6.250 146.610 ;
        RECT 7.090 145.720 12.690 146.610 ;
        RECT 13.530 145.720 15.910 146.610 ;
        RECT 16.750 145.720 22.350 146.610 ;
        RECT 23.190 145.720 25.570 146.610 ;
        RECT 26.410 145.720 32.010 146.610 ;
        RECT 32.850 145.720 35.230 146.610 ;
        RECT 36.070 145.720 38.450 146.610 ;
        RECT 39.290 145.720 44.890 146.610 ;
        RECT 45.730 145.720 48.110 146.610 ;
        RECT 48.950 145.720 54.550 146.610 ;
        RECT 55.390 145.720 57.770 146.610 ;
        RECT 58.610 145.720 60.990 146.610 ;
        RECT 61.830 145.720 67.430 146.610 ;
        RECT 68.270 145.720 70.650 146.610 ;
        RECT 71.490 145.720 77.090 146.610 ;
        RECT 77.930 145.720 80.310 146.610 ;
        RECT 81.150 145.720 86.750 146.610 ;
        RECT 87.590 145.720 89.970 146.610 ;
        RECT 90.810 145.720 93.190 146.610 ;
        RECT 94.030 145.720 99.630 146.610 ;
        RECT 100.470 145.720 102.850 146.610 ;
        RECT 103.690 145.720 109.290 146.610 ;
        RECT 110.130 145.720 112.510 146.610 ;
        RECT 113.350 145.720 118.950 146.610 ;
        RECT 119.790 145.720 122.170 146.610 ;
        RECT 123.010 145.720 125.390 146.610 ;
        RECT 126.230 145.720 131.830 146.610 ;
        RECT 132.670 145.720 135.050 146.610 ;
        RECT 135.890 145.720 141.490 146.610 ;
        RECT 142.330 145.720 144.710 146.610 ;
        RECT 145.550 145.720 147.930 146.610 ;
        RECT 148.770 145.720 154.370 146.610 ;
        RECT 155.210 145.720 157.590 146.610 ;
        RECT 158.430 145.720 164.030 146.610 ;
        RECT 164.870 145.720 167.250 146.610 ;
        RECT 168.090 145.720 173.690 146.610 ;
        RECT 174.530 145.720 176.910 146.610 ;
        RECT 177.750 145.720 180.130 146.610 ;
        RECT 180.970 145.720 186.570 146.610 ;
        RECT 187.410 145.720 189.790 146.610 ;
        RECT 190.630 145.720 196.230 146.610 ;
        RECT 197.070 145.720 199.450 146.610 ;
        RECT 200.290 145.720 205.890 146.610 ;
        RECT 206.730 145.720 209.110 146.610 ;
        RECT 209.950 145.720 212.330 146.610 ;
        RECT 213.170 145.720 218.770 146.610 ;
        RECT 219.610 145.720 221.990 146.610 ;
        RECT 222.830 145.720 228.430 146.610 ;
        RECT 229.270 145.720 231.650 146.610 ;
        RECT 232.490 145.720 234.870 146.610 ;
        RECT 235.710 145.720 241.310 146.610 ;
        RECT 242.150 145.720 244.530 146.610 ;
        RECT 245.370 145.720 250.970 146.610 ;
        RECT 251.810 145.720 254.190 146.610 ;
        RECT 255.030 145.720 260.630 146.610 ;
        RECT 261.470 145.720 263.850 146.610 ;
        RECT 264.690 145.720 267.070 146.610 ;
        RECT 267.910 145.720 273.510 146.610 ;
        RECT 274.350 145.720 276.730 146.610 ;
        RECT 277.570 145.720 283.170 146.610 ;
        RECT 284.010 145.720 286.390 146.610 ;
        RECT 287.230 145.720 292.830 146.610 ;
        RECT 293.670 145.720 296.050 146.610 ;
        RECT 296.890 145.720 299.270 146.610 ;
        RECT 300.110 145.720 305.710 146.610 ;
        RECT 306.550 145.720 308.930 146.610 ;
        RECT 309.770 145.720 315.370 146.610 ;
        RECT 316.210 145.720 318.590 146.610 ;
        RECT 319.430 145.720 321.810 146.610 ;
        RECT 322.650 145.720 328.250 146.610 ;
        RECT 329.090 145.720 331.470 146.610 ;
        RECT 332.310 145.720 337.910 146.610 ;
        RECT 338.750 145.720 341.130 146.610 ;
        RECT 341.970 145.720 347.570 146.610 ;
        RECT 348.410 145.720 350.790 146.610 ;
        RECT 351.630 145.720 354.010 146.610 ;
        RECT 354.850 145.720 360.450 146.610 ;
        RECT 361.290 145.720 363.670 146.610 ;
        RECT 364.510 145.720 370.110 146.610 ;
        RECT 370.950 145.720 373.330 146.610 ;
        RECT 374.170 145.720 379.770 146.610 ;
        RECT 380.610 145.720 382.990 146.610 ;
        RECT 383.830 145.720 386.210 146.610 ;
        RECT 387.050 145.720 392.650 146.610 ;
        RECT 393.490 145.720 395.870 146.610 ;
        RECT 396.710 145.720 402.310 146.610 ;
        RECT 403.150 145.720 405.530 146.610 ;
        RECT 406.370 145.720 411.970 146.610 ;
        RECT 412.810 145.720 415.190 146.610 ;
        RECT 416.030 145.720 418.410 146.610 ;
        RECT 419.250 145.720 424.850 146.610 ;
        RECT 425.690 145.720 428.070 146.610 ;
        RECT 428.910 145.720 434.510 146.610 ;
        RECT 435.350 145.720 437.730 146.610 ;
        RECT 438.570 145.720 440.950 146.610 ;
        RECT 441.790 145.720 447.390 146.610 ;
        RECT 448.230 145.720 450.610 146.610 ;
        RECT 451.450 145.720 457.050 146.610 ;
        RECT 457.890 145.720 460.270 146.610 ;
        RECT 461.110 145.720 466.710 146.610 ;
        RECT 467.550 145.720 469.930 146.610 ;
        RECT 470.770 145.720 473.150 146.610 ;
        RECT 473.990 145.720 479.590 146.610 ;
        RECT 480.430 145.720 482.810 146.610 ;
        RECT 483.650 145.720 489.250 146.610 ;
        RECT 490.090 145.720 492.470 146.610 ;
        RECT 493.310 145.720 498.910 146.610 ;
        RECT 499.750 145.720 502.130 146.610 ;
        RECT 502.970 145.720 505.350 146.610 ;
        RECT 506.190 145.720 511.790 146.610 ;
        RECT 512.630 145.720 515.010 146.610 ;
        RECT 515.850 145.720 521.450 146.610 ;
        RECT 522.290 145.720 524.670 146.610 ;
        RECT 525.510 145.720 527.890 146.610 ;
        RECT 528.730 145.720 534.330 146.610 ;
        RECT 535.170 145.720 537.550 146.610 ;
        RECT 538.390 145.720 543.990 146.610 ;
        RECT 544.830 145.720 547.210 146.610 ;
        RECT 548.050 145.720 553.650 146.610 ;
        RECT 554.490 145.720 556.870 146.610 ;
        RECT 557.710 145.720 560.090 146.610 ;
        RECT 560.930 145.720 566.530 146.610 ;
        RECT 567.370 145.720 569.750 146.610 ;
        RECT 570.590 145.720 576.190 146.610 ;
        RECT 577.030 145.720 579.410 146.610 ;
        RECT 580.250 145.720 585.850 146.610 ;
        RECT 586.690 145.720 589.070 146.610 ;
        RECT 589.910 145.720 592.290 146.610 ;
        RECT 593.130 145.720 598.730 146.610 ;
        RECT 0.100 4.280 599.280 145.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 99.630 4.280 ;
        RECT 100.470 0.155 102.850 4.280 ;
        RECT 103.690 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 141.490 4.280 ;
        RECT 142.330 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.930 4.280 ;
        RECT 148.770 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 164.030 4.280 ;
        RECT 164.870 0.155 167.250 4.280 ;
        RECT 168.090 0.155 173.690 4.280 ;
        RECT 174.530 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 186.570 4.280 ;
        RECT 187.410 0.155 189.790 4.280 ;
        RECT 190.630 0.155 196.230 4.280 ;
        RECT 197.070 0.155 199.450 4.280 ;
        RECT 200.290 0.155 202.670 4.280 ;
        RECT 203.510 0.155 209.110 4.280 ;
        RECT 209.950 0.155 212.330 4.280 ;
        RECT 213.170 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.990 4.280 ;
        RECT 222.830 0.155 228.430 4.280 ;
        RECT 229.270 0.155 231.650 4.280 ;
        RECT 232.490 0.155 234.870 4.280 ;
        RECT 235.710 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 250.970 4.280 ;
        RECT 251.810 0.155 254.190 4.280 ;
        RECT 255.030 0.155 260.630 4.280 ;
        RECT 261.470 0.155 263.850 4.280 ;
        RECT 264.690 0.155 267.070 4.280 ;
        RECT 267.910 0.155 273.510 4.280 ;
        RECT 274.350 0.155 276.730 4.280 ;
        RECT 277.570 0.155 283.170 4.280 ;
        RECT 284.010 0.155 286.390 4.280 ;
        RECT 287.230 0.155 289.610 4.280 ;
        RECT 290.450 0.155 296.050 4.280 ;
        RECT 296.890 0.155 299.270 4.280 ;
        RECT 300.110 0.155 305.710 4.280 ;
        RECT 306.550 0.155 308.930 4.280 ;
        RECT 309.770 0.155 315.370 4.280 ;
        RECT 316.210 0.155 318.590 4.280 ;
        RECT 319.430 0.155 321.810 4.280 ;
        RECT 322.650 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.470 4.280 ;
        RECT 332.310 0.155 337.910 4.280 ;
        RECT 338.750 0.155 341.130 4.280 ;
        RECT 341.970 0.155 347.570 4.280 ;
        RECT 348.410 0.155 350.790 4.280 ;
        RECT 351.630 0.155 354.010 4.280 ;
        RECT 354.850 0.155 360.450 4.280 ;
        RECT 361.290 0.155 363.670 4.280 ;
        RECT 364.510 0.155 370.110 4.280 ;
        RECT 370.950 0.155 373.330 4.280 ;
        RECT 374.170 0.155 376.550 4.280 ;
        RECT 377.390 0.155 382.990 4.280 ;
        RECT 383.830 0.155 386.210 4.280 ;
        RECT 387.050 0.155 392.650 4.280 ;
        RECT 393.490 0.155 395.870 4.280 ;
        RECT 396.710 0.155 402.310 4.280 ;
        RECT 403.150 0.155 405.530 4.280 ;
        RECT 406.370 0.155 408.750 4.280 ;
        RECT 409.590 0.155 415.190 4.280 ;
        RECT 416.030 0.155 418.410 4.280 ;
        RECT 419.250 0.155 424.850 4.280 ;
        RECT 425.690 0.155 428.070 4.280 ;
        RECT 428.910 0.155 434.510 4.280 ;
        RECT 435.350 0.155 437.730 4.280 ;
        RECT 438.570 0.155 440.950 4.280 ;
        RECT 441.790 0.155 447.390 4.280 ;
        RECT 448.230 0.155 450.610 4.280 ;
        RECT 451.450 0.155 457.050 4.280 ;
        RECT 457.890 0.155 460.270 4.280 ;
        RECT 461.110 0.155 463.490 4.280 ;
        RECT 464.330 0.155 469.930 4.280 ;
        RECT 470.770 0.155 473.150 4.280 ;
        RECT 473.990 0.155 479.590 4.280 ;
        RECT 480.430 0.155 482.810 4.280 ;
        RECT 483.650 0.155 489.250 4.280 ;
        RECT 490.090 0.155 492.470 4.280 ;
        RECT 493.310 0.155 495.690 4.280 ;
        RECT 496.530 0.155 502.130 4.280 ;
        RECT 502.970 0.155 505.350 4.280 ;
        RECT 506.190 0.155 511.790 4.280 ;
        RECT 512.630 0.155 515.010 4.280 ;
        RECT 515.850 0.155 521.450 4.280 ;
        RECT 522.290 0.155 524.670 4.280 ;
        RECT 525.510 0.155 527.890 4.280 ;
        RECT 528.730 0.155 534.330 4.280 ;
        RECT 535.170 0.155 537.550 4.280 ;
        RECT 538.390 0.155 543.990 4.280 ;
        RECT 544.830 0.155 547.210 4.280 ;
        RECT 548.050 0.155 553.650 4.280 ;
        RECT 554.490 0.155 556.870 4.280 ;
        RECT 557.710 0.155 560.090 4.280 ;
        RECT 560.930 0.155 566.530 4.280 ;
        RECT 567.370 0.155 569.750 4.280 ;
        RECT 570.590 0.155 576.190 4.280 ;
        RECT 577.030 0.155 579.410 4.280 ;
        RECT 580.250 0.155 582.630 4.280 ;
        RECT 583.470 0.155 589.070 4.280 ;
        RECT 589.910 0.155 592.290 4.280 ;
        RECT 593.130 0.155 598.730 4.280 ;
      LAYER met3 ;
        RECT 4.000 145.840 595.600 146.690 ;
        RECT 4.000 143.840 596.000 145.840 ;
        RECT 4.400 142.440 596.000 143.840 ;
        RECT 4.000 140.440 596.000 142.440 ;
        RECT 4.400 139.040 595.600 140.440 ;
        RECT 4.000 137.040 596.000 139.040 ;
        RECT 4.000 135.640 595.600 137.040 ;
        RECT 4.000 133.640 596.000 135.640 ;
        RECT 4.400 132.240 595.600 133.640 ;
        RECT 4.000 130.240 596.000 132.240 ;
        RECT 4.400 128.840 596.000 130.240 ;
        RECT 4.000 126.840 596.000 128.840 ;
        RECT 4.000 125.440 595.600 126.840 ;
        RECT 4.000 123.440 596.000 125.440 ;
        RECT 4.400 122.040 595.600 123.440 ;
        RECT 4.000 120.040 596.000 122.040 ;
        RECT 4.400 118.640 596.000 120.040 ;
        RECT 4.000 116.640 596.000 118.640 ;
        RECT 4.400 115.240 595.600 116.640 ;
        RECT 4.000 113.240 596.000 115.240 ;
        RECT 4.000 111.840 595.600 113.240 ;
        RECT 4.000 109.840 596.000 111.840 ;
        RECT 4.400 108.440 596.000 109.840 ;
        RECT 4.000 106.440 596.000 108.440 ;
        RECT 4.400 105.040 595.600 106.440 ;
        RECT 4.000 103.040 596.000 105.040 ;
        RECT 4.000 101.640 595.600 103.040 ;
        RECT 4.000 99.640 596.000 101.640 ;
        RECT 4.400 98.240 595.600 99.640 ;
        RECT 4.000 96.240 596.000 98.240 ;
        RECT 4.400 94.840 596.000 96.240 ;
        RECT 4.000 92.840 596.000 94.840 ;
        RECT 4.400 91.440 595.600 92.840 ;
        RECT 4.000 89.440 596.000 91.440 ;
        RECT 4.000 88.040 595.600 89.440 ;
        RECT 4.000 86.040 596.000 88.040 ;
        RECT 4.400 84.640 596.000 86.040 ;
        RECT 4.000 82.640 596.000 84.640 ;
        RECT 4.400 81.240 595.600 82.640 ;
        RECT 4.000 79.240 596.000 81.240 ;
        RECT 4.000 77.840 595.600 79.240 ;
        RECT 4.000 75.840 596.000 77.840 ;
        RECT 4.400 74.440 596.000 75.840 ;
        RECT 4.000 72.440 596.000 74.440 ;
        RECT 4.400 71.040 595.600 72.440 ;
        RECT 4.000 69.040 596.000 71.040 ;
        RECT 4.000 67.640 595.600 69.040 ;
        RECT 4.000 65.640 596.000 67.640 ;
        RECT 4.400 64.240 595.600 65.640 ;
        RECT 4.000 62.240 596.000 64.240 ;
        RECT 4.400 60.840 596.000 62.240 ;
        RECT 4.000 58.840 596.000 60.840 ;
        RECT 4.400 57.440 595.600 58.840 ;
        RECT 4.000 55.440 596.000 57.440 ;
        RECT 4.000 54.040 595.600 55.440 ;
        RECT 4.000 52.040 596.000 54.040 ;
        RECT 4.400 50.640 596.000 52.040 ;
        RECT 4.000 48.640 596.000 50.640 ;
        RECT 4.400 47.240 595.600 48.640 ;
        RECT 4.000 45.240 596.000 47.240 ;
        RECT 4.000 43.840 595.600 45.240 ;
        RECT 4.000 41.840 596.000 43.840 ;
        RECT 4.400 40.440 595.600 41.840 ;
        RECT 4.000 38.440 596.000 40.440 ;
        RECT 4.400 37.040 596.000 38.440 ;
        RECT 4.000 35.040 596.000 37.040 ;
        RECT 4.000 33.640 595.600 35.040 ;
        RECT 4.000 31.640 596.000 33.640 ;
        RECT 4.400 30.240 595.600 31.640 ;
        RECT 4.000 28.240 596.000 30.240 ;
        RECT 4.400 26.840 596.000 28.240 ;
        RECT 4.000 24.840 596.000 26.840 ;
        RECT 4.400 23.440 595.600 24.840 ;
        RECT 4.000 21.440 596.000 23.440 ;
        RECT 4.000 20.040 595.600 21.440 ;
        RECT 4.000 18.040 596.000 20.040 ;
        RECT 4.400 16.640 596.000 18.040 ;
        RECT 4.000 14.640 596.000 16.640 ;
        RECT 4.400 13.240 595.600 14.640 ;
        RECT 4.000 11.240 596.000 13.240 ;
        RECT 4.000 9.840 595.600 11.240 ;
        RECT 4.000 7.840 596.000 9.840 ;
        RECT 4.400 6.440 595.600 7.840 ;
        RECT 4.000 4.440 596.000 6.440 ;
        RECT 4.400 3.040 596.000 4.440 ;
        RECT 4.000 1.040 596.000 3.040 ;
        RECT 4.000 0.175 595.600 1.040 ;
      LAYER met4 ;
        RECT 351.735 131.415 353.905 134.450 ;
  END
END bus_arbiter
END LIBRARY

