magic
tech sky130B
magscale 1 2
timestamp 1662026868
<< obsli1 >>
rect 0 0 584000 704000
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 63402 702788 63408 702840
rect 63460 702828 63466 702840
rect 218974 702828 218980 702840
rect 63460 702800 218980 702828
rect 63460 702788 63466 702800
rect 218974 702788 218980 702800
rect 219032 702788 219038 702840
rect 412634 702788 412640 702840
rect 412692 702828 412698 702840
rect 413646 702828 413652 702840
rect 412692 702800 413652 702828
rect 412692 702788 412698 702800
rect 413646 702788 413652 702800
rect 413704 702788 413710 702840
rect 72970 702720 72976 702772
rect 73028 702760 73034 702772
rect 245654 702760 245660 702772
rect 73028 702732 245660 702760
rect 73028 702720 73034 702732
rect 245654 702720 245660 702732
rect 245712 702720 245718 702772
rect 53742 702652 53748 702704
rect 53800 702692 53806 702704
rect 202782 702692 202788 702704
rect 53800 702664 202788 702692
rect 53800 702652 53806 702664
rect 202782 702652 202788 702664
rect 202840 702692 202846 702704
rect 416774 702692 416780 702704
rect 202840 702664 416780 702692
rect 202840 702652 202846 702664
rect 416774 702652 416780 702664
rect 416832 702652 416838 702704
rect 40494 702584 40500 702636
rect 40552 702624 40558 702636
rect 217318 702624 217324 702636
rect 40552 702596 217324 702624
rect 40552 702584 40558 702596
rect 217318 702584 217324 702596
rect 217376 702584 217382 702636
rect 300118 702584 300124 702636
rect 300176 702624 300182 702636
rect 538214 702624 538220 702636
rect 300176 702596 538220 702624
rect 300176 702584 300182 702596
rect 538214 702584 538220 702596
rect 538272 702584 538278 702636
rect 8110 702516 8116 702568
rect 8168 702556 8174 702568
rect 210418 702556 210424 702568
rect 8168 702528 210424 702556
rect 8168 702516 8174 702528
rect 210418 702516 210424 702528
rect 210476 702516 210482 702568
rect 251082 702516 251088 702568
rect 251140 702556 251146 702568
rect 527174 702556 527180 702568
rect 251140 702528 527180 702556
rect 251140 702516 251146 702528
rect 527174 702516 527180 702528
rect 527232 702516 527238 702568
rect 130378 702448 130384 702500
rect 130436 702488 130442 702500
rect 412634 702488 412640 702500
rect 130436 702460 412640 702488
rect 130436 702448 130442 702460
rect 412634 702448 412640 702460
rect 412692 702448 412698 702500
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 269114 700380 269120 700392
rect 235224 700352 269120 700380
rect 235224 700340 235230 700352
rect 269114 700340 269120 700352
rect 269172 700340 269178 700392
rect 359458 700340 359464 700392
rect 359516 700380 359522 700392
rect 397454 700380 397460 700392
rect 359516 700352 397460 700380
rect 359516 700340 359522 700352
rect 397454 700340 397460 700352
rect 397512 700340 397518 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 39298 700312 39304 700324
rect 24360 700284 39304 700312
rect 24360 700272 24366 700284
rect 39298 700272 39304 700284
rect 39356 700272 39362 700324
rect 52362 700272 52368 700324
rect 52420 700312 52426 700324
rect 137830 700312 137836 700324
rect 52420 700284 137836 700312
rect 52420 700272 52426 700284
rect 137830 700272 137836 700284
rect 137888 700272 137894 700324
rect 154114 700272 154120 700324
rect 154172 700312 154178 700324
rect 247034 700312 247040 700324
rect 154172 700284 247040 700312
rect 154172 700272 154178 700284
rect 247034 700272 247040 700284
rect 247092 700272 247098 700324
rect 332410 700272 332416 700324
rect 332468 700312 332474 700324
rect 429838 700312 429844 700324
rect 332468 700284 429844 700312
rect 332468 700272 332474 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 494790 700272 494796 700324
rect 494848 700312 494854 700324
rect 518158 700312 518164 700324
rect 494848 700284 518164 700312
rect 494848 700272 494854 700284
rect 518158 700272 518164 700284
rect 518216 700272 518222 700324
rect 102778 699660 102784 699712
rect 102836 699700 102842 699712
rect 105446 699700 105452 699712
rect 102836 699672 105452 699700
rect 102836 699660 102842 699672
rect 105446 699660 105452 699672
rect 105504 699660 105510 699712
rect 261478 699660 261484 699712
rect 261536 699700 261542 699712
rect 300118 699700 300124 699712
rect 261536 699672 300124 699700
rect 261536 699660 261542 699672
rect 300118 699660 300124 699672
rect 300176 699660 300182 699712
rect 348786 699660 348792 699712
rect 348844 699700 348850 699712
rect 351178 699700 351184 699712
rect 348844 699672 351184 699700
rect 348844 699660 348850 699672
rect 351178 699660 351184 699672
rect 351236 699660 351242 699712
rect 540238 699660 540244 699712
rect 540296 699700 540302 699712
rect 543458 699700 543464 699712
rect 540296 699672 543464 699700
rect 540296 699660 540302 699672
rect 543458 699660 543464 699672
rect 543516 699660 543522 699712
rect 552658 699660 552664 699712
rect 552716 699700 552722 699712
rect 559650 699700 559656 699712
rect 552716 699672 559656 699700
rect 552716 699660 552722 699672
rect 559650 699660 559656 699672
rect 559708 699660 559714 699712
rect 265618 698912 265624 698964
rect 265676 698952 265682 698964
rect 348786 698952 348792 698964
rect 265676 698924 348792 698952
rect 265676 698912 265682 698924
rect 348786 698912 348792 698924
rect 348844 698912 348850 698964
rect 570598 696940 570604 696992
rect 570656 696980 570662 696992
rect 580166 696980 580172 696992
rect 570656 696952 580172 696980
rect 570656 696940 570662 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 7558 683176 7564 683188
rect 3476 683148 7564 683176
rect 3476 683136 3482 683148
rect 7558 683136 7564 683148
rect 7616 683136 7622 683188
rect 549898 683136 549904 683188
rect 549956 683176 549962 683188
rect 580166 683176 580172 683188
rect 549956 683148 580172 683176
rect 549956 683136 549962 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 542998 670692 543004 670744
rect 543056 670732 543062 670744
rect 580166 670732 580172 670744
rect 543056 670704 580172 670732
rect 543056 670692 543062 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 18598 656928 18604 656940
rect 3476 656900 18604 656928
rect 3476 656888 3482 656900
rect 18598 656888 18604 656900
rect 18656 656888 18662 656940
rect 338758 643084 338764 643136
rect 338816 643124 338822 643136
rect 580166 643124 580172 643136
rect 338816 643096 580172 643124
rect 338816 643084 338822 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 351178 632680 351184 632732
rect 351236 632720 351242 632732
rect 488534 632720 488540 632732
rect 351236 632692 488540 632720
rect 351236 632680 351242 632692
rect 488534 632680 488540 632692
rect 488592 632680 488598 632732
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 17218 632108 17224 632120
rect 3476 632080 17224 632108
rect 3476 632068 3482 632080
rect 17218 632068 17224 632080
rect 17276 632068 17282 632120
rect 337930 630640 337936 630692
rect 337988 630680 337994 630692
rect 580166 630680 580172 630692
rect 337988 630652 580172 630680
rect 337988 630640 337994 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 39298 620236 39304 620288
rect 39356 620276 39362 620288
rect 51074 620276 51080 620288
rect 39356 620248 51080 620276
rect 39356 620236 39362 620248
rect 51074 620236 51080 620248
rect 51132 620236 51138 620288
rect 220722 620236 220728 620288
rect 220780 620276 220786 620288
rect 282914 620276 282920 620288
rect 220780 620248 282920 620276
rect 220780 620236 220786 620248
rect 282914 620236 282920 620248
rect 282972 620236 282978 620288
rect 51074 619624 51080 619676
rect 51132 619664 51138 619676
rect 52270 619664 52276 619676
rect 51132 619636 52276 619664
rect 51132 619624 51138 619636
rect 52270 619624 52276 619636
rect 52328 619664 52334 619676
rect 185578 619664 185584 619676
rect 52328 619636 185584 619664
rect 52328 619624 52334 619636
rect 185578 619624 185584 619636
rect 185636 619624 185642 619676
rect 88334 618876 88340 618928
rect 88392 618916 88398 618928
rect 236638 618916 236644 618928
rect 88392 618888 236644 618916
rect 88392 618876 88398 618888
rect 236638 618876 236644 618888
rect 236696 618876 236702 618928
rect 412634 618876 412640 618928
rect 412692 618916 412698 618928
rect 534350 618916 534356 618928
rect 412692 618888 534356 618916
rect 412692 618876 412698 618888
rect 534350 618876 534356 618888
rect 534408 618876 534414 618928
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 40678 618304 40684 618316
rect 3200 618276 40684 618304
rect 3200 618264 3206 618276
rect 40678 618264 40684 618276
rect 40736 618264 40742 618316
rect 289722 618264 289728 618316
rect 289780 618304 289786 618316
rect 456794 618304 456800 618316
rect 289780 618276 456800 618304
rect 289780 618264 289786 618276
rect 456794 618264 456800 618276
rect 456852 618264 456858 618316
rect 17218 617516 17224 617568
rect 17276 617556 17282 617568
rect 229094 617556 229100 617568
rect 17276 617528 229100 617556
rect 17276 617516 17282 617528
rect 229094 617516 229100 617528
rect 229152 617516 229158 617568
rect 391014 616836 391020 616888
rect 391072 616876 391078 616888
rect 580166 616876 580172 616888
rect 391072 616848 580172 616876
rect 391072 616836 391078 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 358078 616700 358084 616752
rect 358136 616740 358142 616752
rect 359458 616740 359464 616752
rect 358136 616712 359464 616740
rect 358136 616700 358142 616712
rect 359458 616700 359464 616712
rect 359516 616700 359522 616752
rect 227622 616088 227628 616140
rect 227680 616128 227686 616140
rect 331214 616128 331220 616140
rect 227680 616100 331220 616128
rect 227680 616088 227686 616100
rect 331214 616088 331220 616100
rect 331272 616088 331278 616140
rect 400858 616088 400864 616140
rect 400916 616128 400922 616140
rect 552658 616128 552664 616140
rect 400916 616100 552664 616128
rect 400916 616088 400922 616100
rect 552658 616088 552664 616100
rect 552716 616088 552722 616140
rect 260098 615476 260104 615528
rect 260156 615516 260162 615528
rect 510614 615516 510620 615528
rect 260156 615488 510620 615516
rect 260156 615476 260162 615488
rect 510614 615476 510620 615488
rect 510672 615476 510678 615528
rect 169754 614728 169760 614780
rect 169812 614768 169818 614780
rect 245838 614768 245844 614780
rect 169812 614740 245844 614768
rect 169812 614728 169818 614740
rect 245838 614728 245844 614740
rect 245896 614728 245902 614780
rect 288342 614184 288348 614236
rect 288400 614224 288406 614236
rect 483842 614224 483848 614236
rect 288400 614196 483848 614224
rect 288400 614184 288406 614196
rect 483842 614184 483848 614196
rect 483900 614184 483906 614236
rect 229462 614116 229468 614168
rect 229520 614156 229526 614168
rect 264238 614156 264244 614168
rect 229520 614128 264244 614156
rect 229520 614116 229526 614128
rect 264238 614116 264244 614128
rect 264296 614156 264302 614168
rect 536926 614156 536932 614168
rect 264296 614128 536932 614156
rect 264296 614116 264302 614128
rect 536926 614116 536932 614128
rect 536984 614116 536990 614168
rect 338022 613368 338028 613420
rect 338080 613408 338086 613420
rect 364334 613408 364340 613420
rect 338080 613380 364340 613408
rect 338080 613368 338086 613380
rect 364334 613368 364340 613380
rect 364392 613368 364398 613420
rect 420178 613368 420184 613420
rect 420236 613408 420242 613420
rect 477494 613408 477500 613420
rect 420236 613380 477500 613408
rect 420236 613368 420242 613380
rect 477494 613368 477500 613380
rect 477552 613368 477558 613420
rect 289078 612824 289084 612876
rect 289136 612864 289142 612876
rect 390554 612864 390560 612876
rect 289136 612836 390560 612864
rect 289136 612824 289142 612836
rect 390554 612824 390560 612836
rect 390612 612864 390618 612876
rect 391014 612864 391020 612876
rect 390612 612836 391020 612864
rect 390612 612824 390618 612836
rect 391014 612824 391020 612836
rect 391072 612824 391078 612876
rect 300210 612756 300216 612808
rect 300268 612796 300274 612808
rect 493502 612796 493508 612808
rect 300268 612768 493508 612796
rect 300268 612756 300274 612768
rect 493502 612756 493508 612768
rect 493560 612756 493566 612808
rect 537018 612688 537024 612740
rect 537076 612728 537082 612740
rect 540238 612728 540244 612740
rect 537076 612700 540244 612728
rect 537076 612688 537082 612700
rect 540238 612688 540244 612700
rect 540296 612688 540302 612740
rect 275278 611464 275284 611516
rect 275336 611504 275342 611516
rect 402974 611504 402980 611516
rect 275336 611476 402980 611504
rect 275336 611464 275342 611476
rect 402974 611464 402980 611476
rect 403032 611464 403038 611516
rect 327902 611396 327908 611448
rect 327960 611436 327966 611448
rect 537018 611436 537024 611448
rect 327960 611408 537024 611436
rect 327960 611396 327966 611408
rect 537018 611396 537024 611408
rect 537076 611396 537082 611448
rect 178678 611328 178684 611380
rect 178736 611368 178742 611380
rect 450354 611368 450360 611380
rect 178736 611340 450360 611368
rect 178736 611328 178742 611340
rect 450354 611328 450360 611340
rect 450412 611328 450418 611380
rect 292390 610104 292396 610156
rect 292448 610144 292454 610156
rect 388530 610144 388536 610156
rect 292448 610116 388536 610144
rect 292448 610104 292454 610116
rect 388530 610104 388536 610116
rect 388588 610104 388594 610156
rect 223022 610036 223028 610088
rect 223080 610076 223086 610088
rect 249794 610076 249800 610088
rect 223080 610048 249800 610076
rect 223080 610036 223086 610048
rect 249794 610036 249800 610048
rect 249852 610076 249858 610088
rect 491294 610076 491300 610088
rect 249852 610048 491300 610076
rect 249852 610036 249858 610048
rect 491294 610036 491300 610048
rect 491352 610036 491358 610088
rect 191098 609968 191104 610020
rect 191156 610008 191162 610020
rect 469674 610008 469680 610020
rect 191156 609980 469680 610008
rect 191156 609968 191162 609980
rect 469674 609968 469680 609980
rect 469732 609968 469738 610020
rect 273898 608744 273904 608796
rect 273956 608784 273962 608796
rect 431954 608784 431960 608796
rect 273956 608756 431960 608784
rect 273956 608744 273962 608756
rect 431954 608744 431960 608756
rect 432012 608744 432018 608796
rect 207566 608676 207572 608728
rect 207624 608716 207630 608728
rect 253934 608716 253940 608728
rect 207624 608688 253940 608716
rect 207624 608676 207630 608688
rect 253934 608676 253940 608688
rect 253992 608716 253998 608728
rect 436186 608716 436192 608728
rect 253992 608688 436192 608716
rect 253992 608676 253998 608688
rect 436186 608676 436192 608688
rect 436244 608676 436250 608728
rect 232682 608608 232688 608660
rect 232740 608648 232746 608660
rect 252554 608648 252560 608660
rect 232740 608620 252560 608648
rect 232740 608608 232746 608620
rect 252554 608608 252560 608620
rect 252612 608648 252618 608660
rect 498654 608648 498660 608660
rect 252612 608620 498660 608648
rect 252612 608608 252618 608620
rect 498654 608608 498660 608620
rect 498712 608608 498718 608660
rect 462314 607860 462320 607912
rect 462372 607900 462378 607912
rect 534258 607900 534264 607912
rect 462372 607872 534264 607900
rect 462372 607860 462378 607872
rect 534258 607860 534264 607872
rect 534316 607860 534322 607912
rect 306282 607384 306288 607436
rect 306340 607424 306346 607436
rect 452930 607424 452936 607436
rect 306340 607396 452936 607424
rect 306340 607384 306346 607396
rect 452930 607384 452936 607396
rect 452988 607384 452994 607436
rect 169018 607316 169024 607368
rect 169076 607356 169082 607368
rect 412634 607356 412640 607368
rect 169076 607328 412640 607356
rect 169076 607316 169082 607328
rect 412634 607316 412640 607328
rect 412692 607316 412698 607368
rect 295978 607248 295984 607300
rect 296036 607288 296042 607300
rect 562318 607288 562324 607300
rect 296036 607260 562324 607288
rect 296036 607248 296042 607260
rect 562318 607248 562324 607260
rect 562376 607248 562382 607300
rect 63126 607180 63132 607232
rect 63184 607220 63190 607232
rect 443270 607220 443276 607232
rect 63184 607192 443276 607220
rect 63184 607180 63190 607192
rect 443270 607180 443276 607192
rect 443328 607180 443334 607232
rect 319438 606092 319444 606144
rect 319496 606132 319502 606144
rect 378870 606132 378876 606144
rect 319496 606104 378876 606132
rect 319496 606092 319502 606104
rect 378870 606092 378876 606104
rect 378928 606092 378934 606144
rect 324222 606024 324228 606076
rect 324280 606064 324286 606076
rect 448514 606064 448520 606076
rect 324280 606036 448520 606064
rect 324280 606024 324286 606036
rect 448514 606024 448520 606036
rect 448572 606024 448578 606076
rect 333330 605956 333336 606008
rect 333388 605996 333394 606008
rect 520274 605996 520280 606008
rect 333388 605968 520280 605996
rect 333388 605956 333394 605968
rect 520274 605956 520280 605968
rect 520332 605956 520338 606008
rect 119338 605888 119344 605940
rect 119396 605928 119402 605940
rect 409874 605928 409880 605940
rect 119396 605900 409880 605928
rect 119396 605888 119402 605900
rect 409874 605888 409880 605900
rect 409932 605888 409938 605940
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 46198 605860 46204 605872
rect 3292 605832 46204 605860
rect 3292 605820 3298 605832
rect 46198 605820 46204 605832
rect 46256 605820 46262 605872
rect 63494 605820 63500 605872
rect 63552 605860 63558 605872
rect 459554 605860 459560 605872
rect 63552 605832 459560 605860
rect 63552 605820 63558 605832
rect 459554 605820 459560 605832
rect 459612 605820 459618 605872
rect 357434 605140 357440 605192
rect 357492 605180 357498 605192
rect 358078 605180 358084 605192
rect 357492 605152 358084 605180
rect 357492 605140 357498 605152
rect 358078 605140 358084 605152
rect 358136 605140 358142 605192
rect 332502 604732 332508 604784
rect 332560 604772 332566 604784
rect 400214 604772 400220 604784
rect 332560 604744 400220 604772
rect 332560 604732 332566 604744
rect 400214 604732 400220 604744
rect 400272 604772 400278 604784
rect 400858 604772 400864 604784
rect 400272 604744 400864 604772
rect 400272 604732 400278 604744
rect 400858 604732 400864 604744
rect 400916 604732 400922 604784
rect 287698 604664 287704 604716
rect 287756 604704 287762 604716
rect 357434 604704 357440 604716
rect 287756 604676 357440 604704
rect 287756 604664 287762 604676
rect 357434 604664 357440 604676
rect 357492 604664 357498 604716
rect 308398 604596 308404 604648
rect 308456 604636 308462 604648
rect 386414 604636 386420 604648
rect 308456 604608 386420 604636
rect 308456 604596 308462 604608
rect 386414 604596 386420 604608
rect 386472 604596 386478 604648
rect 166258 604528 166264 604580
rect 166316 604568 166322 604580
rect 312538 604568 312544 604580
rect 166316 604540 312544 604568
rect 166316 604528 166322 604540
rect 312538 604528 312544 604540
rect 312596 604568 312602 604580
rect 396074 604568 396080 604580
rect 312596 604540 396080 604568
rect 312596 604528 312602 604540
rect 396074 604528 396080 604540
rect 396132 604528 396138 604580
rect 86218 604460 86224 604512
rect 86276 604500 86282 604512
rect 524414 604500 524420 604512
rect 86276 604472 524420 604500
rect 86276 604460 86282 604472
rect 524414 604460 524420 604472
rect 524472 604460 524478 604512
rect 321462 603304 321468 603356
rect 321520 603344 321526 603356
rect 423950 603344 423956 603356
rect 321520 603316 423956 603344
rect 321520 603304 321526 603316
rect 423950 603304 423956 603316
rect 424008 603304 424014 603356
rect 251174 603276 251180 603288
rect 238726 603248 251180 603276
rect 204346 603168 204352 603220
rect 204404 603208 204410 603220
rect 238726 603208 238754 603248
rect 251174 603236 251180 603248
rect 251232 603276 251238 603288
rect 414382 603276 414388 603288
rect 251232 603248 414388 603276
rect 251232 603236 251238 603248
rect 414382 603236 414388 603248
rect 414440 603236 414446 603288
rect 204404 603180 238754 603208
rect 204404 603168 204410 603180
rect 252462 603168 252468 603220
rect 252520 603208 252526 603220
rect 486878 603208 486884 603220
rect 252520 603180 486884 603208
rect 252520 603168 252526 603180
rect 486878 603168 486884 603180
rect 486936 603168 486942 603220
rect 63310 603100 63316 603152
rect 63368 603140 63374 603152
rect 381446 603140 381452 603152
rect 63368 603112 381452 603140
rect 63368 603100 63374 603112
rect 381446 603100 381452 603112
rect 381504 603100 381510 603152
rect 283558 602012 283564 602064
rect 283616 602052 283622 602064
rect 376754 602052 376760 602064
rect 283616 602024 376760 602052
rect 283616 602012 283622 602024
rect 376754 602012 376760 602024
rect 376812 602012 376818 602064
rect 298002 601944 298008 601996
rect 298060 601984 298066 601996
rect 398190 601984 398196 601996
rect 298060 601956 398196 601984
rect 298060 601944 298066 601956
rect 398190 601944 398196 601956
rect 398248 601944 398254 601996
rect 339034 601876 339040 601928
rect 339092 601916 339098 601928
rect 496078 601916 496084 601928
rect 339092 601888 496084 601916
rect 339092 601876 339098 601888
rect 496078 601876 496084 601888
rect 496136 601876 496142 601928
rect 317230 601808 317236 601860
rect 317288 601848 317294 601860
rect 536834 601848 536840 601860
rect 317288 601820 536840 601848
rect 317288 601808 317294 601820
rect 536834 601808 536840 601820
rect 536892 601808 536898 601860
rect 305638 601740 305644 601792
rect 305696 601780 305702 601792
rect 549254 601780 549260 601792
rect 305696 601752 549260 601780
rect 305696 601740 305702 601752
rect 549254 601740 549260 601752
rect 549312 601780 549318 601792
rect 549898 601780 549904 601792
rect 549312 601752 549904 601780
rect 549312 601740 549318 601752
rect 549898 601740 549904 601752
rect 549956 601740 549962 601792
rect 112438 601672 112444 601724
rect 112496 601712 112502 601724
rect 440694 601712 440700 601724
rect 112496 601684 440700 601712
rect 112496 601672 112502 601684
rect 440694 601672 440700 601684
rect 440752 601672 440758 601724
rect 307018 600652 307024 600704
rect 307076 600692 307082 600704
rect 393314 600692 393320 600704
rect 307076 600664 393320 600692
rect 307076 600652 307082 600664
rect 393314 600652 393320 600664
rect 393372 600652 393378 600704
rect 336642 600584 336648 600636
rect 336700 600624 336706 600636
rect 474182 600624 474188 600636
rect 336700 600596 474188 600624
rect 336700 600584 336706 600596
rect 474182 600584 474188 600596
rect 474240 600584 474246 600636
rect 334802 600516 334808 600568
rect 334860 600556 334866 600568
rect 500954 600556 500960 600568
rect 334860 600528 500960 600556
rect 334860 600516 334866 600528
rect 500954 600516 500960 600528
rect 501012 600516 501018 600568
rect 253198 600448 253204 600500
rect 253256 600488 253262 600500
rect 438854 600488 438860 600500
rect 253256 600460 438860 600488
rect 253256 600448 253262 600460
rect 438854 600448 438860 600460
rect 438912 600448 438918 600500
rect 134518 600380 134524 600432
rect 134576 600420 134582 600432
rect 349890 600420 349896 600432
rect 134576 600392 349896 600420
rect 134576 600380 134582 600392
rect 349890 600380 349896 600392
rect 349948 600380 349954 600432
rect 17218 600312 17224 600364
rect 17276 600352 17282 600364
rect 373994 600352 374000 600364
rect 17276 600324 374000 600352
rect 17276 600312 17282 600324
rect 373994 600312 374000 600324
rect 374052 600312 374058 600364
rect 376754 600312 376760 600364
rect 376812 600352 376818 600364
rect 544470 600352 544476 600364
rect 376812 600324 544476 600352
rect 376812 600312 376818 600324
rect 544470 600312 544476 600324
rect 544528 600312 544534 600364
rect 331858 599292 331864 599344
rect 331916 599332 331922 599344
rect 347958 599332 347964 599344
rect 331916 599304 347964 599332
rect 331916 599292 331922 599304
rect 347958 599292 347964 599304
rect 348016 599292 348022 599344
rect 311802 599224 311808 599276
rect 311860 599264 311866 599276
rect 371786 599264 371792 599276
rect 311860 599236 371792 599264
rect 311860 599224 311866 599236
rect 371786 599224 371792 599236
rect 371844 599224 371850 599276
rect 327810 599156 327816 599208
rect 327868 599196 327874 599208
rect 415394 599196 415400 599208
rect 327868 599168 415400 599196
rect 327868 599156 327874 599168
rect 415394 599156 415400 599168
rect 415452 599156 415458 599208
rect 327718 599088 327724 599140
rect 327776 599128 327782 599140
rect 422294 599128 422300 599140
rect 327776 599100 422300 599128
rect 327776 599088 327782 599100
rect 422294 599088 422300 599100
rect 422352 599088 422358 599140
rect 512822 599088 512828 599140
rect 512880 599128 512886 599140
rect 542446 599128 542452 599140
rect 512880 599100 542452 599128
rect 512880 599088 512886 599100
rect 542446 599088 542452 599100
rect 542504 599088 542510 599140
rect 334710 599020 334716 599072
rect 334768 599060 334774 599072
rect 537018 599060 537024 599072
rect 334768 599032 537024 599060
rect 334768 599020 334774 599032
rect 537018 599020 537024 599032
rect 537076 599020 537082 599072
rect 80698 598952 80704 599004
rect 80756 598992 80762 599004
rect 534074 598992 534080 599004
rect 80756 598964 534080 598992
rect 80756 598952 80762 598964
rect 534074 598952 534080 598964
rect 534132 598952 534138 599004
rect 414382 598204 414388 598256
rect 414440 598244 414446 598256
rect 482002 598244 482008 598256
rect 414440 598216 482008 598244
rect 414440 598204 414446 598216
rect 482002 598204 482008 598216
rect 482060 598204 482066 598256
rect 140222 597864 140228 597916
rect 140280 597904 140286 597916
rect 407298 597904 407304 597916
rect 140280 597876 407304 597904
rect 140280 597864 140286 597876
rect 407298 597864 407304 597876
rect 407356 597864 407362 597916
rect 518158 597864 518164 597916
rect 518216 597904 518222 597916
rect 552014 597904 552020 597916
rect 518216 597876 552020 597904
rect 518216 597864 518222 597876
rect 552014 597864 552020 597876
rect 552072 597864 552078 597916
rect 333422 597796 333428 597848
rect 333480 597836 333486 597848
rect 345474 597836 345480 597848
rect 333480 597808 345480 597836
rect 333480 597796 333486 597808
rect 345474 597796 345480 597808
rect 345532 597796 345538 597848
rect 503622 597796 503628 597848
rect 503680 597836 503686 597848
rect 547874 597836 547880 597848
rect 503680 597808 547880 597836
rect 503680 597796 503686 597808
rect 547874 597796 547880 597808
rect 547932 597796 547938 597848
rect 326430 597728 326436 597780
rect 326488 597768 326494 597780
rect 367094 597768 367100 597780
rect 326488 597740 367100 597768
rect 326488 597728 326494 597740
rect 367094 597728 367100 597740
rect 367152 597728 367158 597780
rect 477402 597728 477408 597780
rect 477460 597768 477466 597780
rect 538306 597768 538312 597780
rect 477460 597740 538312 597768
rect 477460 597728 477466 597740
rect 538306 597728 538312 597740
rect 538364 597728 538370 597780
rect 339678 597660 339684 597712
rect 339736 597700 339742 597712
rect 405734 597700 405740 597712
rect 339736 597672 405740 597700
rect 339736 597660 339742 597672
rect 405734 597660 405740 597672
rect 405792 597660 405798 597712
rect 472986 597660 472992 597712
rect 473044 597700 473050 597712
rect 543734 597700 543740 597712
rect 473044 597672 543740 597700
rect 473044 597660 473050 597672
rect 543734 597660 543740 597672
rect 543792 597660 543798 597712
rect 279418 597592 279424 597644
rect 279476 597632 279482 597644
rect 369302 597632 369308 597644
rect 279476 597604 369308 597632
rect 279476 597592 279482 597604
rect 369302 597592 369308 597604
rect 369360 597592 369366 597644
rect 486878 597592 486884 597644
rect 486936 597632 486942 597644
rect 574738 597632 574744 597644
rect 486936 597604 574744 597632
rect 486936 597592 486942 597604
rect 574738 597592 574744 597604
rect 574796 597592 574802 597644
rect 407022 597524 407028 597576
rect 407080 597564 407086 597576
rect 527174 597564 527180 597576
rect 407080 597536 527180 597564
rect 407080 597524 407086 597536
rect 527174 597524 527180 597536
rect 527232 597524 527238 597576
rect 532602 597524 532608 597576
rect 532660 597564 532666 597576
rect 561674 597564 561680 597576
rect 532660 597536 561680 597564
rect 532660 597524 532666 597536
rect 561674 597524 561680 597536
rect 561732 597524 561738 597576
rect 235994 597456 236000 597508
rect 236052 597496 236058 597508
rect 236638 597496 236644 597508
rect 236052 597468 236644 597496
rect 236052 597456 236058 597468
rect 236638 597456 236644 597468
rect 236696 597456 236702 597508
rect 90358 596776 90364 596828
rect 90416 596816 90422 596828
rect 102778 596816 102784 596828
rect 90416 596788 102784 596816
rect 90416 596776 90422 596788
rect 102778 596776 102784 596788
rect 102836 596776 102842 596828
rect 323578 596504 323584 596556
rect 323636 596544 323642 596556
rect 465258 596544 465264 596556
rect 323636 596516 465264 596544
rect 323636 596504 323642 596516
rect 465258 596504 465264 596516
rect 465316 596504 465322 596556
rect 329190 596436 329196 596488
rect 329248 596476 329254 596488
rect 539686 596476 539692 596488
rect 329248 596448 539692 596476
rect 329248 596436 329254 596448
rect 539686 596436 539692 596448
rect 539744 596436 539750 596488
rect 309042 596368 309048 596420
rect 309100 596408 309106 596420
rect 535546 596408 535552 596420
rect 309100 596380 535552 596408
rect 309100 596368 309106 596380
rect 535546 596368 535552 596380
rect 535604 596368 535610 596420
rect 153838 596300 153844 596352
rect 153896 596340 153902 596352
rect 383654 596340 383660 596352
rect 153896 596312 383660 596340
rect 153896 596300 153902 596312
rect 383654 596300 383660 596312
rect 383712 596300 383718 596352
rect 331030 596232 331036 596284
rect 331088 596272 331094 596284
rect 582374 596272 582380 596284
rect 331088 596244 582380 596272
rect 331088 596232 331094 596244
rect 582374 596232 582380 596244
rect 582432 596232 582438 596284
rect 38562 596164 38568 596216
rect 38620 596204 38626 596216
rect 143534 596204 143540 596216
rect 38620 596176 143540 596204
rect 38620 596164 38626 596176
rect 143534 596164 143540 596176
rect 143592 596164 143598 596216
rect 235994 596164 236000 596216
rect 236052 596204 236058 596216
rect 256602 596204 256608 596216
rect 236052 596176 256608 596204
rect 236052 596164 236058 596176
rect 256602 596164 256608 596176
rect 256660 596204 256666 596216
rect 529934 596204 529940 596216
rect 256660 596176 529940 596204
rect 256660 596164 256666 596176
rect 529934 596164 529940 596176
rect 529992 596164 529998 596216
rect 220722 596096 220728 596148
rect 220780 596136 220786 596148
rect 407022 596136 407028 596148
rect 220780 596108 407028 596136
rect 220780 596096 220786 596108
rect 407022 596096 407028 596108
rect 407080 596096 407086 596148
rect 569954 595620 569960 595672
rect 570012 595660 570018 595672
rect 570598 595660 570604 595672
rect 570012 595632 570604 595660
rect 570012 595620 570018 595632
rect 570598 595620 570604 595632
rect 570656 595620 570662 595672
rect 459554 595484 459560 595536
rect 459612 595524 459618 595536
rect 460428 595524 460434 595536
rect 459612 595496 460434 595524
rect 459612 595484 459618 595496
rect 460428 595484 460434 595496
rect 460486 595484 460492 595536
rect 92934 595416 92940 595468
rect 92992 595456 92998 595468
rect 317414 595456 317420 595468
rect 92992 595428 317420 595456
rect 92992 595416 92998 595428
rect 317414 595416 317420 595428
rect 317472 595416 317478 595468
rect 325050 595076 325056 595128
rect 325108 595116 325114 595128
rect 352558 595116 352564 595128
rect 325108 595088 352564 595116
rect 325108 595076 325114 595088
rect 352558 595076 352564 595088
rect 352616 595076 352622 595128
rect 460566 595076 460572 595128
rect 460624 595116 460630 595128
rect 544378 595116 544384 595128
rect 460624 595088 544384 595116
rect 460624 595076 460630 595088
rect 544378 595076 544384 595088
rect 544436 595076 544442 595128
rect 338850 595008 338856 595060
rect 338908 595048 338914 595060
rect 426618 595048 426624 595060
rect 338908 595020 426624 595048
rect 338908 595008 338914 595020
rect 426618 595008 426624 595020
rect 426676 595008 426682 595060
rect 456242 595008 456248 595060
rect 456300 595048 456306 595060
rect 553486 595048 553492 595060
rect 456300 595020 553492 595048
rect 456300 595008 456306 595020
rect 553486 595008 553492 595020
rect 553544 595008 553550 595060
rect 337838 594940 337844 594992
rect 337896 594980 337902 594992
rect 538858 594980 538864 594992
rect 337896 594952 538864 594980
rect 337896 594940 337902 594952
rect 538858 594940 538864 594952
rect 538916 594940 538922 594992
rect 318058 594872 318064 594924
rect 318116 594912 318122 594924
rect 535822 594912 535828 594924
rect 318116 594884 535828 594912
rect 318116 594872 318122 594884
rect 535822 594872 535828 594884
rect 535880 594872 535886 594924
rect 53558 594804 53564 594856
rect 53616 594844 53622 594856
rect 140590 594844 140596 594856
rect 53616 594816 140596 594844
rect 53616 594804 53622 594816
rect 140590 594804 140596 594816
rect 140648 594804 140654 594856
rect 331950 594804 331956 594856
rect 332008 594844 332014 594856
rect 569954 594844 569960 594856
rect 332008 594816 569960 594844
rect 332008 594804 332014 594816
rect 569954 594804 569960 594816
rect 570012 594804 570018 594856
rect 339494 594736 339500 594788
rect 339552 594776 339558 594788
rect 342898 594776 342904 594788
rect 339552 594748 342904 594776
rect 339552 594736 339558 594748
rect 342898 594736 342904 594748
rect 342956 594736 342962 594788
rect 535638 594532 535644 594584
rect 535696 594572 535702 594584
rect 537110 594572 537116 594584
rect 535696 594544 537116 594572
rect 535696 594532 535702 594544
rect 537110 594532 537116 594544
rect 537168 594532 537174 594584
rect 127618 594056 127624 594108
rect 127676 594096 127682 594108
rect 339494 594096 339500 594108
rect 127676 594068 339500 594096
rect 127676 594056 127682 594068
rect 339494 594056 339500 594068
rect 339552 594056 339558 594108
rect 54938 593376 54944 593428
rect 54996 593416 55002 593428
rect 169018 593416 169024 593428
rect 54996 593388 169024 593416
rect 54996 593376 55002 593388
rect 169018 593376 169024 593388
rect 169076 593416 169082 593428
rect 169570 593416 169576 593428
rect 169076 593388 169576 593416
rect 169076 593376 169082 593388
rect 169570 593376 169576 593388
rect 169628 593376 169634 593428
rect 143810 593308 143816 593360
rect 143868 593348 143874 593360
rect 339678 593348 339684 593360
rect 143868 593320 339684 593348
rect 143868 593308 143874 593320
rect 339678 593308 339684 593320
rect 339736 593308 339742 593360
rect 45462 592084 45468 592136
rect 45520 592124 45526 592136
rect 127618 592124 127624 592136
rect 45520 592096 127624 592124
rect 45520 592084 45526 592096
rect 127618 592084 127624 592096
rect 127676 592084 127682 592136
rect 39942 592016 39948 592068
rect 40000 592056 40006 592068
rect 163222 592056 163228 592068
rect 40000 592028 163228 592056
rect 40000 592016 40006 592028
rect 163222 592016 163228 592028
rect 163280 592016 163286 592068
rect 55030 591268 55036 591320
rect 55088 591308 55094 591320
rect 327902 591308 327908 591320
rect 55088 591280 327908 591308
rect 55088 591268 55094 591280
rect 327902 591268 327908 591280
rect 327960 591268 327966 591320
rect 562318 591268 562324 591320
rect 562376 591308 562382 591320
rect 579798 591308 579804 591320
rect 562376 591280 579804 591308
rect 562376 591268 562382 591280
rect 579798 591268 579804 591280
rect 579856 591268 579862 591320
rect 59998 590860 60004 590912
rect 60056 590900 60062 590912
rect 86218 590900 86224 590912
rect 60056 590872 86224 590900
rect 60056 590860 60062 590872
rect 86218 590860 86224 590872
rect 86276 590900 86282 590912
rect 86494 590900 86500 590912
rect 86276 590872 86500 590900
rect 86276 590860 86282 590872
rect 86494 590860 86500 590872
rect 86552 590860 86558 590912
rect 41322 590792 41328 590844
rect 41380 590832 41386 590844
rect 92934 590832 92940 590844
rect 41380 590804 92940 590832
rect 41380 590792 41386 590804
rect 92934 590792 92940 590804
rect 92992 590792 92998 590844
rect 48130 590724 48136 590776
rect 48188 590764 48194 590776
rect 159910 590764 159916 590776
rect 48188 590736 159916 590764
rect 48188 590724 48194 590736
rect 159910 590724 159916 590736
rect 159968 590724 159974 590776
rect 56318 590656 56324 590708
rect 56376 590696 56382 590708
rect 191098 590696 191104 590708
rect 56376 590668 191104 590696
rect 56376 590656 56382 590668
rect 191098 590656 191104 590668
rect 191156 590696 191162 590708
rect 191466 590696 191472 590708
rect 191156 590668 191472 590696
rect 191156 590656 191162 590668
rect 191466 590656 191472 590668
rect 191524 590656 191530 590708
rect 197262 590656 197268 590708
rect 197320 590696 197326 590708
rect 273990 590696 273996 590708
rect 197320 590668 273996 590696
rect 197320 590656 197326 590668
rect 273990 590656 273996 590668
rect 274048 590656 274054 590708
rect 535638 590656 535644 590708
rect 535696 590696 535702 590708
rect 554038 590696 554044 590708
rect 535696 590668 554044 590696
rect 535696 590656 535702 590668
rect 554038 590656 554044 590668
rect 554096 590656 554102 590708
rect 106182 589908 106188 589960
rect 106240 589948 106246 589960
rect 336550 589948 336556 589960
rect 106240 589920 336556 589948
rect 106240 589908 106246 589920
rect 336550 589908 336556 589920
rect 336608 589908 336614 589960
rect 38470 589500 38476 589552
rect 38528 589540 38534 589552
rect 105814 589540 105820 589552
rect 38528 589512 105820 589540
rect 38528 589500 38534 589512
rect 105814 589500 105820 589512
rect 105872 589540 105878 589552
rect 106182 589540 106188 589552
rect 105872 589512 106188 589540
rect 105872 589500 105878 589512
rect 106182 589500 106188 589512
rect 106240 589500 106246 589552
rect 99374 589432 99380 589484
rect 99432 589472 99438 589484
rect 251818 589472 251824 589484
rect 99432 589444 251824 589472
rect 99432 589432 99438 589444
rect 251818 589432 251824 589444
rect 251876 589432 251882 589484
rect 35802 589364 35808 589416
rect 35860 589404 35866 589416
rect 77478 589404 77484 589416
rect 35860 589376 77484 589404
rect 35860 589364 35866 589376
rect 77478 589364 77484 589376
rect 77536 589404 77542 589416
rect 257338 589404 257344 589416
rect 77536 589376 257344 589404
rect 77536 589364 77542 589376
rect 257338 589364 257344 589376
rect 257396 589364 257402 589416
rect 59078 589296 59084 589348
rect 59136 589336 59142 589348
rect 309778 589336 309784 589348
rect 59136 589308 309784 589336
rect 59136 589296 59142 589308
rect 309778 589296 309784 589308
rect 309836 589296 309842 589348
rect 50338 588276 50344 588328
rect 50396 588316 50402 588328
rect 197262 588316 197268 588328
rect 50396 588288 197268 588316
rect 50396 588276 50402 588288
rect 197262 588276 197268 588288
rect 197320 588276 197326 588328
rect 57698 588208 57704 588260
rect 57756 588248 57762 588260
rect 90358 588248 90364 588260
rect 57756 588220 90364 588248
rect 57756 588208 57762 588220
rect 90358 588208 90364 588220
rect 90416 588208 90422 588260
rect 59262 588140 59268 588192
rect 59320 588180 59326 588192
rect 112438 588180 112444 588192
rect 59320 588152 112444 588180
rect 59320 588140 59326 588152
rect 112438 588140 112444 588152
rect 112496 588140 112502 588192
rect 56226 588072 56232 588124
rect 56284 588112 56290 588124
rect 130378 588112 130384 588124
rect 56284 588084 130384 588112
rect 56284 588072 56290 588084
rect 130378 588072 130384 588084
rect 130436 588072 130442 588124
rect 214098 588072 214104 588124
rect 214156 588112 214162 588124
rect 248506 588112 248512 588124
rect 214156 588084 248512 588112
rect 214156 588072 214162 588084
rect 248506 588072 248512 588084
rect 248564 588072 248570 588124
rect 194778 588004 194784 588056
rect 194836 588044 194842 588056
rect 253290 588044 253296 588056
rect 194836 588016 253296 588044
rect 194836 588004 194842 588016
rect 253290 588004 253296 588016
rect 253348 588004 253354 588056
rect 60550 587936 60556 587988
rect 60608 587976 60614 587988
rect 153838 587976 153844 587988
rect 60608 587948 153844 587976
rect 60608 587936 60614 587948
rect 153838 587936 153844 587948
rect 153896 587936 153902 587988
rect 163222 587936 163228 587988
rect 163280 587976 163286 587988
rect 318150 587976 318156 587988
rect 163280 587948 318156 587976
rect 163280 587936 163286 587948
rect 318150 587936 318156 587948
rect 318208 587936 318214 587988
rect 8938 587868 8944 587920
rect 8996 587908 9002 587920
rect 172882 587908 172888 587920
rect 8996 587880 172888 587908
rect 8996 587868 9002 587880
rect 172882 587868 172888 587880
rect 172940 587908 172946 587920
rect 266354 587908 266360 587920
rect 172940 587880 266360 587908
rect 172940 587868 172946 587880
rect 266354 587868 266360 587880
rect 266412 587868 266418 587920
rect 324958 587868 324964 587920
rect 325016 587908 325022 587920
rect 337654 587908 337660 587920
rect 325016 587880 337660 587908
rect 325016 587868 325022 587880
rect 337654 587868 337660 587880
rect 337712 587868 337718 587920
rect 197262 587528 197268 587580
rect 197320 587568 197326 587580
rect 197998 587568 198004 587580
rect 197320 587540 198004 587568
rect 197320 587528 197326 587540
rect 197998 587528 198004 587540
rect 198056 587528 198062 587580
rect 299382 587120 299388 587172
rect 299440 587160 299446 587172
rect 337102 587160 337108 587172
rect 299440 587132 337108 587160
rect 299440 587120 299446 587132
rect 337102 587120 337108 587132
rect 337160 587120 337166 587172
rect 49602 586848 49608 586900
rect 49660 586888 49666 586900
rect 83366 586888 83372 586900
rect 49660 586860 83372 586888
rect 49660 586848 49666 586860
rect 83366 586848 83372 586860
rect 83424 586848 83430 586900
rect 49510 586780 49516 586832
rect 49568 586820 49574 586832
rect 96246 586820 96252 586832
rect 49568 586792 96252 586820
rect 49568 586780 49574 586792
rect 96246 586780 96252 586792
rect 96304 586780 96310 586832
rect 122006 586780 122012 586832
rect 122064 586820 122070 586832
rect 244918 586820 244924 586832
rect 122064 586792 244924 586820
rect 122064 586780 122070 586792
rect 244918 586780 244924 586792
rect 244976 586780 244982 586832
rect 63218 586712 63224 586764
rect 63276 586752 63282 586764
rect 137462 586752 137468 586764
rect 63276 586724 137468 586752
rect 63276 586712 63282 586724
rect 137462 586712 137468 586724
rect 137520 586712 137526 586764
rect 217318 586712 217324 586764
rect 217376 586752 217382 586764
rect 245102 586752 245108 586764
rect 217376 586724 245108 586752
rect 217376 586712 217382 586724
rect 245102 586712 245108 586724
rect 245160 586712 245166 586764
rect 57238 586644 57244 586696
rect 57296 586684 57302 586696
rect 166258 586684 166264 586696
rect 57296 586656 166264 586684
rect 57296 586644 57302 586656
rect 166258 586644 166264 586656
rect 166316 586644 166322 586696
rect 201218 586644 201224 586696
rect 201276 586684 201282 586696
rect 217226 586684 217232 586696
rect 201276 586656 217232 586684
rect 201276 586644 201282 586656
rect 217226 586644 217232 586656
rect 217284 586644 217290 586696
rect 239214 586644 239220 586696
rect 239272 586684 239278 586696
rect 277394 586684 277400 586696
rect 239272 586656 277400 586684
rect 239272 586644 239278 586656
rect 277394 586644 277400 586656
rect 277452 586644 277458 586696
rect 31018 586576 31024 586628
rect 31076 586616 31082 586628
rect 147122 586616 147128 586628
rect 31076 586588 147128 586616
rect 31076 586576 31082 586588
rect 147122 586576 147128 586588
rect 147180 586576 147186 586628
rect 181898 586576 181904 586628
rect 181956 586616 181962 586628
rect 243078 586616 243084 586628
rect 181956 586588 243084 586616
rect 181956 586576 181962 586588
rect 243078 586576 243084 586588
rect 243136 586576 243142 586628
rect 44082 586508 44088 586560
rect 44140 586548 44146 586560
rect 125226 586548 125232 586560
rect 44140 586520 125232 586548
rect 44140 586508 44146 586520
rect 125226 586508 125232 586520
rect 125284 586508 125290 586560
rect 50982 585488 50988 585540
rect 51040 585528 51046 585540
rect 67910 585528 67916 585540
rect 51040 585500 67916 585528
rect 51040 585488 51046 585500
rect 67910 585488 67916 585500
rect 67968 585488 67974 585540
rect 46842 585420 46848 585472
rect 46900 585460 46906 585472
rect 102686 585460 102692 585472
rect 46900 585432 102692 585460
rect 46900 585420 46906 585432
rect 102686 585420 102692 585432
rect 102744 585420 102750 585472
rect 15102 585352 15108 585404
rect 15160 585392 15166 585404
rect 71130 585392 71136 585404
rect 15160 585364 71136 585392
rect 15160 585352 15166 585364
rect 71130 585352 71136 585364
rect 71188 585352 71194 585404
rect 226334 585352 226340 585404
rect 226392 585392 226398 585404
rect 227622 585392 227628 585404
rect 226392 585364 227628 585392
rect 226392 585352 226398 585364
rect 227622 585352 227628 585364
rect 227680 585392 227686 585404
rect 247770 585392 247776 585404
rect 227680 585364 247776 585392
rect 227680 585352 227686 585364
rect 247770 585352 247776 585364
rect 247828 585352 247834 585404
rect 60734 585284 60740 585336
rect 60792 585324 60798 585336
rect 150342 585324 150348 585336
rect 60792 585296 150348 585324
rect 60792 585284 60798 585296
rect 150342 585284 150348 585296
rect 150400 585284 150406 585336
rect 185118 585284 185124 585336
rect 185176 585324 185182 585336
rect 185578 585324 185584 585336
rect 185176 585296 185584 585324
rect 185176 585284 185182 585296
rect 185578 585284 185584 585296
rect 185636 585324 185642 585336
rect 247678 585324 247684 585336
rect 185636 585296 247684 585324
rect 185636 585284 185642 585296
rect 247678 585284 247684 585296
rect 247736 585284 247742 585336
rect 48222 585216 48228 585268
rect 48280 585256 48286 585268
rect 109126 585256 109132 585268
rect 48280 585228 109132 585256
rect 48280 585216 48286 585228
rect 109126 585216 109132 585228
rect 109184 585216 109190 585268
rect 137462 585216 137468 585268
rect 137520 585256 137526 585268
rect 260190 585256 260196 585268
rect 137520 585228 260196 585256
rect 137520 585216 137526 585228
rect 260190 585216 260196 585228
rect 260248 585216 260254 585268
rect 35158 585148 35164 585200
rect 35216 585188 35222 585200
rect 255314 585188 255320 585200
rect 35216 585160 255320 585188
rect 35216 585148 35222 585160
rect 255314 585148 255320 585160
rect 255372 585148 255378 585200
rect 333238 585148 333244 585200
rect 333296 585188 333302 585200
rect 337654 585188 337660 585200
rect 333296 585160 337660 585188
rect 333296 585148 333302 585160
rect 337654 585148 337660 585160
rect 337712 585148 337718 585200
rect 217226 585080 217232 585132
rect 217284 585120 217290 585132
rect 295334 585120 295340 585132
rect 217284 585092 295340 585120
rect 217284 585080 217290 585092
rect 295334 585080 295340 585092
rect 295392 585080 295398 585132
rect 295334 584604 295340 584656
rect 295392 584644 295398 584656
rect 295978 584644 295984 584656
rect 295392 584616 295984 584644
rect 295392 584604 295398 584616
rect 295978 584604 295984 584616
rect 296036 584604 296042 584656
rect 61470 584536 61476 584588
rect 61528 584576 61534 584588
rect 245930 584576 245936 584588
rect 61528 584548 245936 584576
rect 61528 584536 61534 584548
rect 245930 584536 245936 584548
rect 245988 584536 245994 584588
rect 292482 583720 292488 583772
rect 292540 583760 292546 583772
rect 337654 583760 337660 583772
rect 292540 583732 337660 583760
rect 292540 583720 292546 583732
rect 337654 583720 337660 583732
rect 337712 583720 337718 583772
rect 245746 582360 245752 582412
rect 245804 582400 245810 582412
rect 318794 582400 318800 582412
rect 245804 582372 318800 582400
rect 245804 582360 245810 582372
rect 318794 582360 318800 582372
rect 318852 582400 318858 582412
rect 320082 582400 320088 582412
rect 318852 582372 320088 582400
rect 318852 582360 318858 582372
rect 320082 582360 320088 582372
rect 320140 582360 320146 582412
rect 245746 582224 245752 582276
rect 245804 582264 245810 582276
rect 245930 582264 245936 582276
rect 245804 582236 245936 582264
rect 245804 582224 245810 582236
rect 245930 582224 245936 582236
rect 245988 582224 245994 582276
rect 297358 581000 297364 581052
rect 297416 581040 297422 581052
rect 337654 581040 337660 581052
rect 297416 581012 337660 581040
rect 297416 581000 297422 581012
rect 337654 581000 337660 581012
rect 337712 581000 337718 581052
rect 535730 581000 535736 581052
rect 535788 581040 535794 581052
rect 563698 581040 563704 581052
rect 535788 581012 563704 581040
rect 535788 581000 535794 581012
rect 563698 581000 563704 581012
rect 563756 581000 563762 581052
rect 244182 580932 244188 580984
rect 244240 580972 244246 580984
rect 336090 580972 336096 580984
rect 244240 580944 336096 580972
rect 244240 580932 244246 580944
rect 336090 580932 336096 580944
rect 336148 580932 336154 580984
rect 242986 580524 242992 580576
rect 243044 580564 243050 580576
rect 243538 580564 243544 580576
rect 243044 580536 243544 580564
rect 243044 580524 243050 580536
rect 243538 580524 243544 580536
rect 243596 580524 243602 580576
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 57606 579680 57612 579692
rect 3384 579652 57612 579680
rect 3384 579640 3390 579652
rect 57606 579640 57612 579652
rect 57664 579680 57670 579692
rect 60734 579680 60740 579692
rect 57664 579652 60740 579680
rect 57664 579640 57670 579652
rect 60734 579640 60740 579652
rect 60792 579640 60798 579692
rect 242986 579640 242992 579692
rect 243044 579680 243050 579692
rect 244182 579680 244188 579692
rect 243044 579652 244188 579680
rect 243044 579640 243050 579652
rect 244182 579640 244188 579652
rect 244240 579640 244246 579692
rect 535730 579164 535736 579216
rect 535788 579204 535794 579216
rect 538214 579204 538220 579216
rect 535788 579176 538220 579204
rect 535788 579164 535794 579176
rect 538214 579164 538220 579176
rect 538272 579164 538278 579216
rect 245102 578892 245108 578944
rect 245160 578932 245166 578944
rect 276014 578932 276020 578944
rect 245160 578904 276020 578932
rect 245160 578892 245166 578904
rect 276014 578892 276020 578904
rect 276072 578892 276078 578944
rect 276014 578212 276020 578264
rect 276072 578252 276078 578264
rect 276658 578252 276664 578264
rect 276072 578224 276664 578252
rect 276072 578212 276078 578224
rect 276658 578212 276664 578224
rect 276716 578252 276722 578264
rect 337654 578252 337660 578264
rect 276716 578224 337660 578252
rect 276716 578212 276722 578224
rect 337654 578212 337660 578224
rect 337712 578212 337718 578264
rect 329742 576852 329748 576904
rect 329800 576892 329806 576904
rect 337654 576892 337660 576904
rect 329800 576864 337660 576892
rect 329800 576852 329806 576864
rect 337654 576852 337660 576864
rect 337712 576852 337718 576904
rect 535730 576852 535736 576904
rect 535788 576892 535794 576904
rect 539594 576892 539600 576904
rect 535788 576864 539600 576892
rect 535788 576852 535794 576864
rect 539594 576852 539600 576864
rect 539652 576852 539658 576904
rect 560938 576852 560944 576904
rect 560996 576892 561002 576904
rect 580166 576892 580172 576904
rect 560996 576864 580172 576892
rect 560996 576852 561002 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 245654 576512 245660 576564
rect 245712 576552 245718 576564
rect 245930 576552 245936 576564
rect 245712 576524 245936 576552
rect 245712 576512 245718 576524
rect 245930 576512 245936 576524
rect 245988 576512 245994 576564
rect 314930 576104 314936 576156
rect 314988 576144 314994 576156
rect 339034 576144 339040 576156
rect 314988 576116 339040 576144
rect 314988 576104 314994 576116
rect 339034 576104 339040 576116
rect 339092 576104 339098 576156
rect 59170 575492 59176 575544
rect 59228 575532 59234 575544
rect 61562 575532 61568 575544
rect 59228 575504 61568 575532
rect 59228 575492 59234 575504
rect 61562 575492 61568 575504
rect 61620 575492 61626 575544
rect 245654 575492 245660 575544
rect 245712 575532 245718 575544
rect 314746 575532 314752 575544
rect 245712 575504 314752 575532
rect 245712 575492 245718 575504
rect 314746 575492 314752 575504
rect 314804 575532 314810 575544
rect 314930 575532 314936 575544
rect 314804 575504 314936 575532
rect 314804 575492 314810 575504
rect 314930 575492 314936 575504
rect 314988 575492 314994 575544
rect 331030 572636 331036 572688
rect 331088 572676 331094 572688
rect 337654 572676 337660 572688
rect 331088 572648 337660 572676
rect 331088 572636 331094 572648
rect 337654 572636 337660 572648
rect 337712 572636 337718 572688
rect 245654 571956 245660 572008
rect 245712 571996 245718 572008
rect 293954 571996 293960 572008
rect 245712 571968 293960 571996
rect 245712 571956 245718 571968
rect 293954 571956 293960 571968
rect 294012 571956 294018 572008
rect 55122 571344 55128 571396
rect 55180 571384 55186 571396
rect 60734 571384 60740 571396
rect 55180 571356 60740 571384
rect 55180 571344 55186 571356
rect 60734 571344 60740 571356
rect 60792 571344 60798 571396
rect 293954 571276 293960 571328
rect 294012 571316 294018 571328
rect 295242 571316 295248 571328
rect 294012 571288 295248 571316
rect 294012 571276 294018 571288
rect 295242 571276 295248 571288
rect 295300 571316 295306 571328
rect 327718 571316 327724 571328
rect 295300 571288 327724 571316
rect 295300 571276 295306 571288
rect 327718 571276 327724 571288
rect 327776 571276 327782 571328
rect 337838 570528 337844 570580
rect 337896 570568 337902 570580
rect 338758 570568 338764 570580
rect 337896 570540 338764 570568
rect 337896 570528 337902 570540
rect 338758 570528 338764 570540
rect 338816 570528 338822 570580
rect 245654 569168 245660 569220
rect 245712 569208 245718 569220
rect 245930 569208 245936 569220
rect 245712 569180 245936 569208
rect 245712 569168 245718 569180
rect 245930 569168 245936 569180
rect 245988 569208 245994 569220
rect 262214 569208 262220 569220
rect 245988 569180 262220 569208
rect 245988 569168 245994 569180
rect 262214 569168 262220 569180
rect 262272 569168 262278 569220
rect 535454 569168 535460 569220
rect 535512 569208 535518 569220
rect 538398 569208 538404 569220
rect 535512 569180 538404 569208
rect 535512 569168 535518 569180
rect 538398 569168 538404 569180
rect 538456 569168 538462 569220
rect 304258 568624 304264 568676
rect 304316 568664 304322 568676
rect 337654 568664 337660 568676
rect 304316 568636 337660 568664
rect 304316 568624 304322 568636
rect 337654 568624 337660 568636
rect 337712 568624 337718 568676
rect 53650 568556 53656 568608
rect 53708 568596 53714 568608
rect 60734 568596 60740 568608
rect 53708 568568 60740 568596
rect 53708 568556 53714 568568
rect 60734 568556 60740 568568
rect 60792 568556 60798 568608
rect 262214 568556 262220 568608
rect 262272 568596 262278 568608
rect 325142 568596 325148 568608
rect 262272 568568 325148 568596
rect 262272 568556 262278 568568
rect 325142 568556 325148 568568
rect 325200 568556 325206 568608
rect 243538 568488 243544 568540
rect 243596 568528 243602 568540
rect 305638 568528 305644 568540
rect 243596 568500 305644 568528
rect 243596 568488 243602 568500
rect 305638 568488 305644 568500
rect 305696 568488 305702 568540
rect 315298 566448 315304 566500
rect 315356 566488 315362 566500
rect 333330 566488 333336 566500
rect 315356 566460 333336 566488
rect 315356 566448 315362 566460
rect 333330 566448 333336 566460
rect 333388 566448 333394 566500
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 22738 565876 22744 565888
rect 3476 565848 22744 565876
rect 3476 565836 3482 565848
rect 22738 565836 22744 565848
rect 22796 565836 22802 565888
rect 245930 565836 245936 565888
rect 245988 565876 245994 565888
rect 314654 565876 314660 565888
rect 245988 565848 314660 565876
rect 245988 565836 245994 565848
rect 314654 565836 314660 565848
rect 314712 565876 314718 565888
rect 315298 565876 315304 565888
rect 314712 565848 315304 565876
rect 314712 565836 314718 565848
rect 315298 565836 315304 565848
rect 315356 565836 315362 565888
rect 27522 564408 27528 564460
rect 27580 564448 27586 564460
rect 60734 564448 60740 564460
rect 27580 564420 60740 564448
rect 27580 564408 27586 564420
rect 60734 564408 60740 564420
rect 60792 564408 60798 564460
rect 535454 563864 535460 563916
rect 535512 563904 535518 563916
rect 538214 563904 538220 563916
rect 535512 563876 538220 563904
rect 535512 563864 535518 563876
rect 538214 563864 538220 563876
rect 538272 563864 538278 563916
rect 538858 563660 538864 563712
rect 538916 563700 538922 563712
rect 575474 563700 575480 563712
rect 538916 563672 575480 563700
rect 538916 563660 538922 563672
rect 575474 563660 575480 563672
rect 575532 563660 575538 563712
rect 575474 563048 575480 563100
rect 575532 563088 575538 563100
rect 579798 563088 579804 563100
rect 575532 563060 579804 563088
rect 575532 563048 575538 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 244918 562300 244924 562352
rect 244976 562340 244982 562352
rect 317322 562340 317328 562352
rect 244976 562312 317328 562340
rect 244976 562300 244982 562312
rect 317322 562300 317328 562312
rect 317380 562300 317386 562352
rect 317322 561688 317328 561740
rect 317380 561728 317386 561740
rect 337378 561728 337384 561740
rect 317380 561700 337384 561728
rect 317380 561688 317386 561700
rect 337378 561688 337384 561700
rect 337436 561688 337442 561740
rect 244918 561620 244924 561672
rect 244976 561660 244982 561672
rect 245562 561660 245568 561672
rect 244976 561632 245568 561660
rect 244976 561620 244982 561632
rect 245562 561620 245568 561632
rect 245620 561660 245626 561672
rect 329190 561660 329196 561672
rect 245620 561632 329196 561660
rect 245620 561620 245626 561632
rect 329190 561620 329196 561632
rect 329248 561620 329254 561672
rect 250438 560260 250444 560312
rect 250496 560300 250502 560312
rect 337654 560300 337660 560312
rect 250496 560272 337660 560300
rect 250496 560260 250502 560272
rect 337654 560260 337660 560272
rect 337712 560260 337718 560312
rect 318150 560192 318156 560244
rect 318208 560232 318214 560244
rect 336918 560232 336924 560244
rect 318208 560204 336924 560232
rect 318208 560192 318214 560204
rect 336918 560192 336924 560204
rect 336976 560192 336982 560244
rect 269022 559512 269028 559564
rect 269080 559552 269086 559564
rect 334802 559552 334808 559564
rect 269080 559524 334808 559552
rect 269080 559512 269086 559524
rect 334802 559512 334808 559524
rect 334860 559512 334866 559564
rect 245930 558900 245936 558952
rect 245988 558940 245994 558952
rect 267734 558940 267740 558952
rect 245988 558912 267740 558940
rect 245988 558900 245994 558912
rect 267734 558900 267740 558912
rect 267792 558940 267798 558952
rect 269022 558940 269028 558952
rect 267792 558912 269028 558940
rect 267792 558900 267798 558912
rect 269022 558900 269028 558912
rect 269080 558900 269086 558952
rect 249702 556792 249708 556844
rect 249760 556832 249766 556844
rect 337930 556832 337936 556844
rect 249760 556804 337936 556832
rect 249760 556792 249766 556804
rect 337930 556792 337936 556804
rect 337988 556792 337994 556844
rect 59078 556112 59084 556164
rect 59136 556152 59142 556164
rect 60734 556152 60740 556164
rect 59136 556124 60740 556152
rect 59136 556112 59142 556124
rect 60734 556112 60740 556124
rect 60792 556112 60798 556164
rect 35710 555432 35716 555484
rect 35768 555472 35774 555484
rect 59078 555472 59084 555484
rect 35768 555444 59084 555472
rect 35768 555432 35774 555444
rect 59078 555432 59084 555444
rect 59136 555432 59142 555484
rect 3142 554684 3148 554736
rect 3200 554724 3206 554736
rect 35158 554724 35164 554736
rect 3200 554696 35164 554724
rect 3200 554684 3206 554696
rect 35158 554684 35164 554696
rect 35216 554684 35222 554736
rect 535454 554684 535460 554736
rect 535512 554724 535518 554736
rect 562318 554724 562324 554736
rect 535512 554696 562324 554724
rect 535512 554684 535518 554696
rect 562318 554684 562324 554696
rect 562376 554684 562382 554736
rect 257246 552644 257252 552696
rect 257304 552684 257310 552696
rect 338942 552684 338948 552696
rect 257304 552656 338948 552684
rect 257304 552644 257310 552656
rect 338942 552644 338948 552656
rect 339000 552644 339006 552696
rect 39850 552032 39856 552084
rect 39908 552072 39914 552084
rect 60734 552072 60740 552084
rect 39908 552044 60740 552072
rect 39908 552032 39914 552044
rect 60734 552032 60740 552044
rect 60792 552032 60798 552084
rect 245930 552032 245936 552084
rect 245988 552072 245994 552084
rect 256694 552072 256700 552084
rect 245988 552044 256700 552072
rect 245988 552032 245994 552044
rect 256694 552032 256700 552044
rect 256752 552072 256758 552084
rect 257246 552072 257252 552084
rect 256752 552044 257252 552072
rect 256752 552032 256758 552044
rect 257246 552032 257252 552044
rect 257304 552032 257310 552084
rect 245654 551284 245660 551336
rect 245712 551324 245718 551336
rect 269758 551324 269764 551336
rect 245712 551296 269764 551324
rect 245712 551284 245718 551296
rect 269758 551284 269764 551296
rect 269816 551284 269822 551336
rect 245930 549244 245936 549296
rect 245988 549284 245994 549296
rect 255222 549284 255228 549296
rect 245988 549256 255228 549284
rect 245988 549244 245994 549256
rect 255222 549244 255228 549256
rect 255280 549244 255286 549296
rect 255240 549216 255268 549244
rect 331950 549216 331956 549228
rect 255240 549188 331956 549216
rect 331950 549176 331956 549188
rect 332008 549176 332014 549228
rect 37182 547884 37188 547936
rect 37240 547924 37246 547936
rect 60734 547924 60740 547936
rect 37240 547896 60740 547924
rect 37240 547884 37246 547896
rect 60734 547884 60740 547896
rect 60792 547884 60798 547936
rect 307202 547884 307208 547936
rect 307260 547924 307266 547936
rect 337654 547924 337660 547936
rect 307260 547896 337660 547924
rect 307260 547884 307266 547896
rect 337654 547884 337660 547896
rect 337712 547884 337718 547936
rect 245930 546456 245936 546508
rect 245988 546496 245994 546508
rect 264330 546496 264336 546508
rect 245988 546468 264336 546496
rect 245988 546456 245994 546468
rect 264330 546456 264336 546468
rect 264388 546456 264394 546508
rect 56502 545776 56508 545828
rect 56560 545816 56566 545828
rect 60734 545816 60740 545828
rect 56560 545788 60740 545816
rect 56560 545776 56566 545788
rect 60734 545776 60740 545788
rect 60792 545776 60798 545828
rect 245286 543668 245292 543720
rect 245344 543708 245350 543720
rect 329098 543708 329104 543720
rect 245344 543680 329104 543708
rect 245344 543668 245350 543680
rect 329098 543668 329104 543680
rect 329156 543668 329162 543720
rect 40678 542376 40684 542428
rect 40736 542416 40742 542428
rect 42794 542416 42800 542428
rect 40736 542388 42800 542416
rect 40736 542376 40742 542388
rect 42794 542376 42800 542388
rect 42852 542416 42858 542428
rect 60734 542416 60740 542428
rect 42852 542388 60740 542416
rect 42852 542376 42858 542388
rect 60734 542376 60740 542388
rect 60792 542376 60798 542428
rect 311158 542376 311164 542428
rect 311216 542416 311222 542428
rect 337654 542416 337660 542428
rect 311216 542388 337660 542416
rect 311216 542376 311222 542388
rect 337654 542376 337660 542388
rect 337712 542376 337718 542428
rect 290458 540948 290464 541000
rect 290516 540988 290522 541000
rect 337470 540988 337476 541000
rect 290516 540960 337476 540988
rect 290516 540948 290522 540960
rect 337470 540948 337476 540960
rect 337528 540948 337534 541000
rect 322198 539520 322204 539572
rect 322256 539560 322262 539572
rect 337654 539560 337660 539572
rect 322256 539532 337660 539560
rect 322256 539520 322262 539532
rect 337654 539520 337660 539532
rect 337712 539520 337718 539572
rect 41230 538228 41236 538280
rect 41288 538268 41294 538280
rect 60734 538268 60740 538280
rect 41288 538240 60740 538268
rect 41288 538228 41294 538240
rect 60734 538228 60740 538240
rect 60792 538228 60798 538280
rect 574738 538160 574744 538212
rect 574796 538200 574802 538212
rect 580166 538200 580172 538212
rect 574796 538172 580172 538200
rect 574796 538160 574802 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 309778 536732 309784 536784
rect 309836 536772 309842 536784
rect 337286 536772 337292 536784
rect 309836 536744 337292 536772
rect 309836 536732 309842 536744
rect 337286 536732 337292 536744
rect 337344 536732 337350 536784
rect 245838 536052 245844 536104
rect 245896 536092 245902 536104
rect 311710 536092 311716 536104
rect 245896 536064 311716 536092
rect 245896 536052 245902 536064
rect 311710 536052 311716 536064
rect 311768 536092 311774 536104
rect 338850 536092 338856 536104
rect 311768 536064 338856 536092
rect 311768 536052 311774 536064
rect 338850 536052 338856 536064
rect 338908 536052 338914 536104
rect 59078 535440 59084 535492
rect 59136 535480 59142 535492
rect 61562 535480 61568 535492
rect 59136 535452 61568 535480
rect 59136 535440 59142 535452
rect 61562 535440 61568 535452
rect 61620 535440 61626 535492
rect 244182 534012 244188 534064
rect 244240 534052 244246 534064
rect 334710 534052 334716 534064
rect 244240 534024 334716 534052
rect 244240 534012 244246 534024
rect 334710 534012 334716 534024
rect 334768 534012 334774 534064
rect 535546 533400 535552 533452
rect 535604 533440 535610 533452
rect 539686 533440 539692 533452
rect 535604 533412 539692 533440
rect 535604 533400 535610 533412
rect 539686 533400 539692 533412
rect 539744 533400 539750 533452
rect 242986 532720 242992 532772
rect 243044 532760 243050 532772
rect 244182 532760 244188 532772
rect 243044 532732 244188 532760
rect 243044 532720 243050 532732
rect 244182 532720 244188 532732
rect 244240 532720 244246 532772
rect 326338 532720 326344 532772
rect 326396 532760 326402 532772
rect 337654 532760 337660 532772
rect 326396 532732 337660 532760
rect 326396 532720 326402 532732
rect 337654 532720 337660 532732
rect 337712 532720 337718 532772
rect 54478 531972 54484 532024
rect 54536 532012 54542 532024
rect 58986 532012 58992 532024
rect 54536 531984 58992 532012
rect 54536 531972 54542 531984
rect 58986 531972 58992 531984
rect 59044 532012 59050 532024
rect 60734 532012 60740 532024
rect 59044 531984 60740 532012
rect 59044 531972 59050 531984
rect 60734 531972 60740 531984
rect 60792 531972 60798 532024
rect 264330 531972 264336 532024
rect 264388 532012 264394 532024
rect 336826 532012 336832 532024
rect 264388 531984 336832 532012
rect 264388 531972 264394 531984
rect 336826 531972 336832 531984
rect 336884 531972 336890 532024
rect 7558 529184 7564 529236
rect 7616 529224 7622 529236
rect 43898 529224 43904 529236
rect 7616 529196 43904 529224
rect 7616 529184 7622 529196
rect 43898 529184 43904 529196
rect 43956 529184 43962 529236
rect 246942 529184 246948 529236
rect 247000 529224 247006 529236
rect 321554 529224 321560 529236
rect 247000 529196 321560 529224
rect 247000 529184 247006 529196
rect 321554 529184 321560 529196
rect 321612 529184 321618 529236
rect 329098 528912 329104 528964
rect 329156 528952 329162 528964
rect 336826 528952 336832 528964
rect 329156 528924 336832 528952
rect 329156 528912 329162 528924
rect 336826 528912 336832 528924
rect 336884 528912 336890 528964
rect 43898 528572 43904 528624
rect 43956 528612 43962 528624
rect 60734 528612 60740 528624
rect 43956 528584 60740 528612
rect 43956 528572 43962 528584
rect 60734 528572 60740 528584
rect 60792 528572 60798 528624
rect 535546 528572 535552 528624
rect 535604 528612 535610 528624
rect 537110 528612 537116 528624
rect 535604 528584 537116 528612
rect 535604 528572 535610 528584
rect 537110 528572 537116 528584
rect 537168 528572 537174 528624
rect 246850 528504 246856 528556
rect 246908 528544 246914 528556
rect 335998 528544 336004 528556
rect 246908 528516 336004 528544
rect 246908 528504 246914 528516
rect 335998 528504 336004 528516
rect 336056 528504 336062 528556
rect 249058 527824 249064 527876
rect 249116 527864 249122 527876
rect 309042 527864 309048 527876
rect 249116 527836 309048 527864
rect 249116 527824 249122 527836
rect 309042 527824 309048 527836
rect 309100 527824 309106 527876
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 48958 527184 48964 527196
rect 3476 527156 6914 527184
rect 3476 527144 3482 527156
rect 6886 526436 6914 527156
rect 21376 527156 48964 527184
rect 21376 527128 21404 527156
rect 48958 527144 48964 527156
rect 49016 527144 49022 527196
rect 246298 527144 246304 527196
rect 246356 527184 246362 527196
rect 246850 527184 246856 527196
rect 246356 527156 246856 527184
rect 246356 527144 246362 527156
rect 246850 527144 246856 527156
rect 246908 527144 246914 527196
rect 309042 527144 309048 527196
rect 309100 527184 309106 527196
rect 309778 527184 309784 527196
rect 309100 527156 309784 527184
rect 309100 527144 309106 527156
rect 309778 527144 309784 527156
rect 309836 527144 309842 527196
rect 21358 527076 21364 527128
rect 21416 527076 21422 527128
rect 269758 527076 269764 527128
rect 269816 527116 269822 527128
rect 317230 527116 317236 527128
rect 269816 527088 317236 527116
rect 269816 527076 269822 527088
rect 317230 527076 317236 527088
rect 317288 527076 317294 527128
rect 21358 526436 21364 526448
rect 6886 526408 21364 526436
rect 21358 526396 21364 526408
rect 21416 526396 21422 526448
rect 314838 526396 314844 526448
rect 314896 526436 314902 526448
rect 337838 526436 337844 526448
rect 314896 526408 337844 526436
rect 314896 526396 314902 526408
rect 337838 526396 337844 526408
rect 337896 526396 337902 526448
rect 264330 525784 264336 525836
rect 264388 525824 264394 525836
rect 314838 525824 314844 525836
rect 264388 525796 314844 525824
rect 264388 525784 264394 525796
rect 314838 525784 314844 525796
rect 314896 525824 314902 525836
rect 315298 525824 315304 525836
rect 314896 525796 315304 525824
rect 314896 525784 314902 525796
rect 315298 525784 315304 525796
rect 315356 525784 315362 525836
rect 317230 525784 317236 525836
rect 317288 525824 317294 525836
rect 317414 525824 317420 525836
rect 317288 525796 317420 525824
rect 317288 525784 317294 525796
rect 317414 525784 317420 525796
rect 317472 525784 317478 525836
rect 53834 525716 53840 525768
rect 53892 525756 53898 525768
rect 55030 525756 55036 525768
rect 53892 525728 55036 525756
rect 53892 525716 53898 525728
rect 55030 525716 55036 525728
rect 55088 525756 55094 525768
rect 60734 525756 60740 525768
rect 55088 525728 60740 525756
rect 55088 525716 55094 525728
rect 60734 525716 60740 525728
rect 60792 525716 60798 525768
rect 544470 525716 544476 525768
rect 544528 525756 544534 525768
rect 579798 525756 579804 525768
rect 544528 525728 579804 525756
rect 544528 525716 544534 525728
rect 579798 525716 579804 525728
rect 579856 525716 579862 525768
rect 33042 525036 33048 525088
rect 33100 525076 33106 525088
rect 53834 525076 53840 525088
rect 33100 525048 53840 525076
rect 33100 525036 33106 525048
rect 53834 525036 53840 525048
rect 53892 525036 53898 525088
rect 300118 525036 300124 525088
rect 300176 525076 300182 525088
rect 337378 525076 337384 525088
rect 300176 525048 337384 525076
rect 300176 525036 300182 525048
rect 337378 525036 337384 525048
rect 337436 525036 337442 525088
rect 55030 524288 55036 524340
rect 55088 524328 55094 524340
rect 57238 524328 57244 524340
rect 55088 524300 57244 524328
rect 55088 524288 55094 524300
rect 57238 524288 57244 524300
rect 57296 524288 57302 524340
rect 535822 523676 535828 523728
rect 535880 523716 535886 523728
rect 536834 523716 536840 523728
rect 535880 523688 536840 523716
rect 535880 523676 535886 523688
rect 536834 523676 536840 523688
rect 536892 523716 536898 523728
rect 558178 523716 558184 523728
rect 536892 523688 558184 523716
rect 536892 523676 536898 523688
rect 558178 523676 558184 523688
rect 558236 523676 558242 523728
rect 307110 522996 307116 523048
rect 307168 523036 307174 523048
rect 337470 523036 337476 523048
rect 307168 523008 337476 523036
rect 307168 522996 307174 523008
rect 337470 522996 337476 523008
rect 337528 522996 337534 523048
rect 245838 521636 245844 521688
rect 245896 521676 245902 521688
rect 303522 521676 303528 521688
rect 245896 521648 303528 521676
rect 245896 521636 245902 521648
rect 303522 521636 303528 521648
rect 303580 521636 303586 521688
rect 314010 520276 314016 520328
rect 314068 520316 314074 520328
rect 337470 520316 337476 520328
rect 314068 520288 337476 520316
rect 314068 520276 314074 520288
rect 337470 520276 337476 520288
rect 337528 520276 337534 520328
rect 535546 520276 535552 520328
rect 535604 520316 535610 520328
rect 549346 520316 549352 520328
rect 535604 520288 549352 520316
rect 535604 520276 535610 520288
rect 549346 520276 549352 520288
rect 549404 520276 549410 520328
rect 245838 518916 245844 518968
rect 245896 518956 245902 518968
rect 270494 518956 270500 518968
rect 245896 518928 270500 518956
rect 245896 518916 245902 518928
rect 270494 518916 270500 518928
rect 270552 518956 270558 518968
rect 335998 518956 336004 518968
rect 270552 518928 336004 518956
rect 270552 518916 270558 518928
rect 335998 518916 336004 518928
rect 336056 518916 336062 518968
rect 535546 518848 535552 518900
rect 535604 518888 535610 518900
rect 549254 518888 549260 518900
rect 535604 518860 549260 518888
rect 535604 518848 535610 518860
rect 549254 518848 549260 518860
rect 549312 518848 549318 518900
rect 3418 516060 3424 516112
rect 3476 516100 3482 516112
rect 61470 516100 61476 516112
rect 3476 516072 61476 516100
rect 3476 516060 3482 516072
rect 61470 516060 61476 516072
rect 61528 516060 61534 516112
rect 535546 515040 535552 515092
rect 535604 515080 535610 515092
rect 538398 515080 538404 515092
rect 535604 515052 538404 515080
rect 535604 515040 535610 515052
rect 538398 515040 538404 515052
rect 538456 515040 538462 515092
rect 250530 514768 250536 514820
rect 250588 514808 250594 514820
rect 337654 514808 337660 514820
rect 250588 514780 337660 514808
rect 250588 514768 250594 514780
rect 337654 514768 337660 514780
rect 337712 514768 337718 514820
rect 305730 513340 305736 513392
rect 305788 513380 305794 513392
rect 337654 513380 337660 513392
rect 305788 513352 337660 513380
rect 305788 513340 305794 513352
rect 337654 513340 337660 513352
rect 337712 513340 337718 513392
rect 535546 513340 535552 513392
rect 535604 513380 535610 513392
rect 548518 513380 548524 513392
rect 535604 513352 548524 513380
rect 535604 513340 535610 513352
rect 548518 513340 548524 513352
rect 548576 513340 548582 513392
rect 245654 513272 245660 513324
rect 245712 513312 245718 513324
rect 264330 513312 264336 513324
rect 245712 513284 264336 513312
rect 245712 513272 245718 513284
rect 264330 513272 264336 513284
rect 264388 513272 264394 513324
rect 563698 511232 563704 511284
rect 563756 511272 563762 511284
rect 579614 511272 579620 511284
rect 563756 511244 579620 511272
rect 563756 511232 563762 511244
rect 579614 511232 579620 511244
rect 579672 511232 579678 511284
rect 330570 510620 330576 510672
rect 330628 510660 330634 510672
rect 337654 510660 337660 510672
rect 330628 510632 337660 510660
rect 330628 510620 330634 510632
rect 337654 510620 337660 510632
rect 337712 510620 337718 510672
rect 245838 509872 245844 509924
rect 245896 509912 245902 509924
rect 251082 509912 251088 509924
rect 245896 509884 251088 509912
rect 245896 509872 245902 509884
rect 251082 509872 251088 509884
rect 251140 509912 251146 509924
rect 259454 509912 259460 509924
rect 251140 509884 259460 509912
rect 251140 509872 251146 509884
rect 259454 509872 259460 509884
rect 259512 509872 259518 509924
rect 535546 507832 535552 507884
rect 535604 507872 535610 507884
rect 550634 507872 550640 507884
rect 535604 507844 550640 507872
rect 535604 507832 535610 507844
rect 550634 507832 550640 507844
rect 550692 507832 550698 507884
rect 255222 507356 255228 507408
rect 255280 507396 255286 507408
rect 258074 507396 258080 507408
rect 255280 507368 258080 507396
rect 255280 507356 255286 507368
rect 258074 507356 258080 507368
rect 258132 507356 258138 507408
rect 535546 506404 535552 506456
rect 535604 506444 535610 506456
rect 569954 506444 569960 506456
rect 535604 506416 569960 506444
rect 535604 506404 535610 506416
rect 569954 506404 569960 506416
rect 570012 506404 570018 506456
rect 245838 505724 245844 505776
rect 245896 505764 245902 505776
rect 255314 505764 255320 505776
rect 245896 505736 255320 505764
rect 245896 505724 245902 505736
rect 255314 505724 255320 505736
rect 255372 505724 255378 505776
rect 260190 505724 260196 505776
rect 260248 505764 260254 505776
rect 310422 505764 310428 505776
rect 260248 505736 310428 505764
rect 260248 505724 260254 505736
rect 310422 505724 310428 505736
rect 310480 505724 310486 505776
rect 310422 505112 310428 505164
rect 310480 505152 310486 505164
rect 337102 505152 337108 505164
rect 310480 505124 337108 505152
rect 310480 505112 310486 505124
rect 337102 505112 337108 505124
rect 337160 505112 337166 505164
rect 57790 504500 57796 504552
rect 57848 504540 57854 504552
rect 62298 504540 62304 504552
rect 57848 504512 62304 504540
rect 57848 504500 57854 504512
rect 62298 504500 62304 504512
rect 62356 504500 62362 504552
rect 255314 504364 255320 504416
rect 255372 504404 255378 504416
rect 311894 504404 311900 504416
rect 255372 504376 311900 504404
rect 255372 504364 255378 504376
rect 311894 504364 311900 504376
rect 311952 504364 311958 504416
rect 311894 503684 311900 503736
rect 311952 503724 311958 503736
rect 312630 503724 312636 503736
rect 311952 503696 312636 503724
rect 311952 503684 311958 503696
rect 312630 503684 312636 503696
rect 312688 503724 312694 503736
rect 337746 503724 337752 503736
rect 312688 503696 337752 503724
rect 312688 503684 312694 503696
rect 337746 503684 337752 503696
rect 337804 503684 337810 503736
rect 251818 502936 251824 502988
rect 251876 502976 251882 502988
rect 303614 502976 303620 502988
rect 251876 502948 303620 502976
rect 251876 502936 251882 502948
rect 303614 502936 303620 502948
rect 303672 502936 303678 502988
rect 303614 502324 303620 502376
rect 303672 502364 303678 502376
rect 304350 502364 304356 502376
rect 303672 502336 304356 502364
rect 303672 502324 303678 502336
rect 304350 502324 304356 502336
rect 304408 502364 304414 502376
rect 337654 502364 337660 502376
rect 304408 502336 337660 502364
rect 304408 502324 304414 502336
rect 337654 502324 337660 502336
rect 337712 502324 337718 502376
rect 535546 502324 535552 502376
rect 535604 502364 535610 502376
rect 546494 502364 546500 502376
rect 535604 502336 546500 502364
rect 535604 502324 535610 502336
rect 546494 502324 546500 502336
rect 546552 502324 546558 502376
rect 246942 501576 246948 501628
rect 247000 501616 247006 501628
rect 322934 501616 322940 501628
rect 247000 501588 322940 501616
rect 247000 501576 247006 501588
rect 322934 501576 322940 501588
rect 322992 501576 322998 501628
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 50430 501004 50436 501016
rect 3108 500976 50436 501004
rect 3108 500964 3114 500976
rect 50430 500964 50436 500976
rect 50488 500964 50494 501016
rect 245838 500488 245844 500540
rect 245896 500528 245902 500540
rect 249058 500528 249064 500540
rect 245896 500500 249064 500528
rect 245896 500488 245902 500500
rect 249058 500488 249064 500500
rect 249116 500488 249122 500540
rect 535546 499536 535552 499588
rect 535604 499576 535610 499588
rect 547966 499576 547972 499588
rect 535604 499548 547972 499576
rect 535604 499536 535610 499548
rect 547966 499536 547972 499548
rect 548024 499536 548030 499588
rect 278038 496816 278044 496868
rect 278096 496856 278102 496868
rect 337654 496856 337660 496868
rect 278096 496828 337660 496856
rect 278096 496816 278102 496828
rect 337654 496816 337660 496828
rect 337712 496816 337718 496868
rect 245838 495456 245844 495508
rect 245896 495496 245902 495508
rect 265710 495496 265716 495508
rect 245896 495468 265716 495496
rect 245896 495456 245902 495468
rect 265710 495456 265716 495468
rect 265768 495456 265774 495508
rect 333330 495456 333336 495508
rect 333388 495496 333394 495508
rect 337470 495496 337476 495508
rect 333388 495468 337476 495496
rect 333388 495456 333394 495468
rect 337470 495456 337476 495468
rect 337528 495456 337534 495508
rect 535546 495456 535552 495508
rect 535604 495496 535610 495508
rect 546586 495496 546592 495508
rect 535604 495468 546592 495496
rect 535604 495456 535610 495468
rect 546586 495456 546592 495468
rect 546644 495456 546650 495508
rect 535546 492668 535552 492720
rect 535604 492708 535610 492720
rect 550726 492708 550732 492720
rect 535604 492680 550732 492708
rect 535604 492668 535610 492680
rect 550726 492668 550732 492680
rect 550784 492668 550790 492720
rect 57882 491308 57888 491360
rect 57940 491348 57946 491360
rect 60734 491348 60740 491360
rect 57940 491320 60740 491348
rect 57940 491308 57946 491320
rect 60734 491308 60740 491320
rect 60792 491308 60798 491360
rect 269758 491308 269764 491360
rect 269816 491348 269822 491360
rect 328270 491348 328276 491360
rect 269816 491320 328276 491348
rect 269816 491308 269822 491320
rect 328270 491308 328276 491320
rect 328328 491348 328334 491360
rect 337470 491348 337476 491360
rect 328328 491320 337476 491348
rect 328328 491308 328334 491320
rect 337470 491308 337476 491320
rect 337528 491308 337534 491360
rect 249058 489880 249064 489932
rect 249116 489920 249122 489932
rect 337654 489920 337660 489932
rect 249116 489892 337660 489920
rect 249116 489880 249122 489892
rect 337654 489880 337660 489892
rect 337712 489880 337718 489932
rect 56410 488520 56416 488572
rect 56468 488560 56474 488572
rect 60734 488560 60740 488572
rect 56468 488532 60740 488560
rect 56468 488520 56474 488532
rect 60734 488520 60740 488532
rect 60792 488520 60798 488572
rect 247770 487772 247776 487824
rect 247828 487812 247834 487824
rect 256786 487812 256792 487824
rect 247828 487784 256792 487812
rect 247828 487772 247834 487784
rect 256786 487772 256792 487784
rect 256844 487772 256850 487824
rect 256786 487160 256792 487212
rect 256844 487200 256850 487212
rect 339310 487200 339316 487212
rect 256844 487172 339316 487200
rect 256844 487160 256850 487172
rect 339310 487160 339316 487172
rect 339368 487160 339374 487212
rect 245838 485800 245844 485852
rect 245896 485840 245902 485852
rect 289170 485840 289176 485852
rect 245896 485812 289176 485840
rect 245896 485800 245902 485812
rect 289170 485800 289176 485812
rect 289228 485800 289234 485852
rect 327718 485800 327724 485852
rect 327776 485840 327782 485852
rect 328270 485840 328276 485852
rect 327776 485812 328276 485840
rect 327776 485800 327782 485812
rect 328270 485800 328276 485812
rect 328328 485800 328334 485852
rect 253290 485052 253296 485104
rect 253348 485092 253354 485104
rect 337746 485092 337752 485104
rect 253348 485064 337752 485092
rect 253348 485052 253354 485064
rect 337746 485052 337752 485064
rect 337804 485052 337810 485104
rect 48038 484372 48044 484424
rect 48096 484412 48102 484424
rect 60734 484412 60740 484424
rect 48096 484384 60740 484412
rect 48096 484372 48102 484384
rect 60734 484372 60740 484384
rect 60792 484372 60798 484424
rect 535546 484372 535552 484424
rect 535604 484412 535610 484424
rect 549438 484412 549444 484424
rect 535604 484384 549444 484412
rect 535604 484372 535610 484384
rect 549438 484372 549444 484384
rect 549496 484372 549502 484424
rect 247678 484304 247684 484356
rect 247736 484344 247742 484356
rect 337930 484344 337936 484356
rect 247736 484316 337936 484344
rect 247736 484304 247742 484316
rect 337930 484304 337936 484316
rect 337988 484304 337994 484356
rect 535546 483012 535552 483064
rect 535604 483052 535610 483064
rect 553394 483052 553400 483064
rect 535604 483024 553400 483052
rect 535604 483012 535610 483024
rect 553394 483012 553400 483024
rect 553452 483012 553458 483064
rect 535546 482876 535552 482928
rect 535604 482916 535610 482928
rect 535730 482916 535736 482928
rect 535604 482888 535736 482916
rect 535604 482876 535610 482888
rect 535730 482876 535736 482888
rect 535788 482876 535794 482928
rect 245746 482264 245752 482316
rect 245804 482304 245810 482316
rect 247678 482304 247684 482316
rect 245804 482276 247684 482304
rect 245804 482264 245810 482276
rect 247678 482264 247684 482276
rect 247736 482304 247742 482316
rect 331858 482304 331864 482316
rect 247736 482276 331864 482304
rect 247736 482264 247742 482276
rect 331858 482264 331864 482276
rect 331916 482264 331922 482316
rect 45370 481652 45376 481704
rect 45428 481692 45434 481704
rect 60734 481692 60740 481704
rect 45428 481664 60740 481692
rect 45428 481652 45434 481664
rect 60734 481652 60740 481664
rect 60792 481652 60798 481704
rect 327902 479476 327908 479528
rect 327960 479516 327966 479528
rect 336734 479516 336740 479528
rect 327960 479488 336740 479516
rect 327960 479476 327966 479488
rect 336734 479476 336740 479488
rect 336792 479476 336798 479528
rect 8202 477504 8208 477556
rect 8260 477544 8266 477556
rect 60734 477544 60740 477556
rect 8260 477516 60740 477544
rect 8260 477504 8266 477516
rect 60734 477504 60740 477516
rect 60792 477504 60798 477556
rect 535730 477504 535736 477556
rect 535788 477544 535794 477556
rect 549254 477544 549260 477556
rect 535788 477516 549260 477544
rect 535788 477504 535794 477516
rect 549254 477504 549260 477516
rect 549312 477504 549318 477556
rect 3878 475328 3884 475380
rect 3936 475368 3942 475380
rect 4798 475368 4804 475380
rect 3936 475340 4804 475368
rect 3936 475328 3942 475340
rect 4798 475328 4804 475340
rect 4856 475368 4862 475380
rect 17218 475368 17224 475380
rect 4856 475340 17224 475368
rect 4856 475328 4862 475340
rect 17218 475328 17224 475340
rect 17276 475328 17282 475380
rect 245746 474716 245752 474768
rect 245804 474756 245810 474768
rect 280798 474756 280804 474768
rect 245804 474728 280804 474756
rect 245804 474716 245810 474728
rect 280798 474716 280804 474728
rect 280856 474716 280862 474768
rect 310422 474716 310428 474768
rect 310480 474756 310486 474768
rect 337654 474756 337660 474768
rect 310480 474728 337660 474756
rect 310480 474716 310486 474728
rect 337654 474716 337660 474728
rect 337712 474716 337718 474768
rect 535730 474716 535736 474768
rect 535788 474756 535794 474768
rect 543826 474756 543832 474768
rect 535788 474728 543832 474756
rect 535788 474716 535794 474728
rect 543826 474716 543832 474728
rect 543884 474716 543890 474768
rect 329282 474104 329288 474156
rect 329340 474144 329346 474156
rect 337746 474144 337752 474156
rect 329340 474116 337752 474144
rect 329340 474104 329346 474116
rect 337746 474104 337752 474116
rect 337804 474104 337810 474156
rect 535730 472200 535736 472252
rect 535788 472240 535794 472252
rect 538490 472240 538496 472252
rect 535788 472212 538496 472240
rect 535788 472200 535794 472212
rect 538490 472200 538496 472212
rect 538548 472200 538554 472252
rect 245838 471996 245844 472048
rect 245896 472036 245902 472048
rect 269206 472036 269212 472048
rect 245896 472008 269212 472036
rect 245896 471996 245902 472008
rect 269206 471996 269212 472008
rect 269264 471996 269270 472048
rect 58986 471656 58992 471708
rect 59044 471696 59050 471708
rect 63402 471696 63408 471708
rect 59044 471668 63408 471696
rect 59044 471656 59050 471668
rect 63402 471656 63408 471668
rect 63460 471656 63466 471708
rect 535730 470568 535736 470620
rect 535788 470608 535794 470620
rect 545206 470608 545212 470620
rect 535788 470580 545212 470608
rect 535788 470568 535794 470580
rect 545206 470568 545212 470580
rect 545264 470568 545270 470620
rect 297910 469820 297916 469872
rect 297968 469860 297974 469872
rect 336734 469860 336740 469872
rect 297968 469832 336740 469860
rect 297968 469820 297974 469832
rect 336734 469820 336740 469832
rect 336792 469820 336798 469872
rect 245838 469140 245844 469192
rect 245896 469180 245902 469192
rect 269758 469180 269764 469192
rect 245896 469152 269764 469180
rect 245896 469140 245902 469152
rect 269758 469140 269764 469152
rect 269816 469140 269822 469192
rect 269206 468460 269212 468512
rect 269264 468500 269270 468512
rect 318702 468500 318708 468512
rect 269264 468472 318708 468500
rect 269264 468460 269270 468472
rect 318702 468460 318708 468472
rect 318760 468500 318766 468512
rect 338022 468500 338028 468512
rect 318760 468472 338028 468500
rect 318760 468460 318766 468472
rect 338022 468460 338028 468472
rect 338080 468460 338086 468512
rect 535730 467984 535736 468036
rect 535788 468024 535794 468036
rect 539686 468024 539692 468036
rect 535788 467996 539692 468024
rect 535788 467984 535794 467996
rect 539686 467984 539692 467996
rect 539744 467984 539750 468036
rect 31662 467848 31668 467900
rect 31720 467888 31726 467900
rect 60734 467888 60740 467900
rect 31720 467860 60740 467888
rect 31720 467848 31726 467860
rect 60734 467848 60740 467860
rect 60792 467848 60798 467900
rect 331950 467440 331956 467492
rect 332008 467480 332014 467492
rect 336826 467480 336832 467492
rect 332008 467452 336832 467480
rect 332008 467440 332014 467452
rect 336826 467440 336832 467452
rect 336884 467440 336890 467492
rect 41138 466420 41144 466472
rect 41196 466460 41202 466472
rect 42794 466460 42800 466472
rect 41196 466432 42800 466460
rect 41196 466420 41202 466432
rect 42794 466420 42800 466432
rect 42852 466420 42858 466472
rect 245838 465060 245844 465112
rect 245896 465100 245902 465112
rect 255314 465100 255320 465112
rect 245896 465072 255320 465100
rect 245896 465060 245902 465072
rect 255314 465060 255320 465072
rect 255372 465060 255378 465112
rect 535730 465060 535736 465112
rect 535788 465100 535794 465112
rect 545298 465100 545304 465112
rect 535788 465072 545304 465100
rect 535788 465060 535794 465072
rect 545298 465060 545304 465072
rect 545356 465060 545362 465112
rect 37090 464312 37096 464364
rect 37148 464352 37154 464364
rect 58986 464352 58992 464364
rect 37148 464324 58992 464352
rect 37148 464312 37154 464324
rect 58986 464312 58992 464324
rect 59044 464312 59050 464364
rect 49418 463700 49424 463752
rect 49476 463740 49482 463752
rect 60734 463740 60740 463752
rect 49476 463712 60740 463740
rect 49476 463700 49482 463712
rect 60734 463700 60740 463712
rect 60792 463700 60798 463752
rect 3418 462612 3424 462664
rect 3476 462652 3482 462664
rect 8938 462652 8944 462664
rect 3476 462624 8944 462652
rect 3476 462612 3482 462624
rect 8938 462612 8944 462624
rect 8996 462612 9002 462664
rect 293954 462340 293960 462392
rect 294012 462380 294018 462392
rect 297358 462380 297364 462392
rect 294012 462352 297364 462380
rect 294012 462340 294018 462352
rect 297358 462340 297364 462352
rect 297416 462340 297422 462392
rect 535730 462340 535736 462392
rect 535788 462380 535794 462392
rect 540974 462380 540980 462392
rect 535788 462352 540980 462380
rect 535788 462340 535794 462352
rect 540974 462340 540980 462352
rect 541032 462340 541038 462392
rect 245838 461592 245844 461644
rect 245896 461632 245902 461644
rect 293954 461632 293960 461644
rect 245896 461604 293960 461632
rect 245896 461592 245902 461604
rect 293954 461592 293960 461604
rect 294012 461592 294018 461644
rect 301498 461592 301504 461644
rect 301556 461632 301562 461644
rect 337654 461632 337660 461644
rect 301556 461604 337660 461632
rect 301556 461592 301562 461604
rect 337654 461592 337660 461604
rect 337712 461592 337718 461644
rect 8938 460912 8944 460964
rect 8996 460952 9002 460964
rect 63126 460952 63132 460964
rect 8996 460924 63132 460952
rect 8996 460912 9002 460924
rect 63126 460912 63132 460924
rect 63184 460912 63190 460964
rect 335262 459552 335268 459604
rect 335320 459592 335326 459604
rect 337654 459592 337660 459604
rect 335320 459564 337660 459592
rect 335320 459552 335326 459564
rect 337654 459552 337660 459564
rect 337712 459552 337718 459604
rect 535730 459552 535736 459604
rect 535788 459592 535794 459604
rect 552106 459592 552112 459604
rect 535788 459564 552112 459592
rect 535788 459552 535794 459564
rect 552106 459552 552112 459564
rect 552164 459552 552170 459604
rect 280062 458804 280068 458856
rect 280120 458844 280126 458856
rect 305730 458844 305736 458856
rect 280120 458816 305736 458844
rect 280120 458804 280126 458816
rect 305730 458804 305736 458816
rect 305788 458804 305794 458856
rect 245838 458192 245844 458244
rect 245896 458232 245902 458244
rect 279510 458232 279516 458244
rect 245896 458204 279516 458232
rect 245896 458192 245902 458204
rect 279510 458192 279516 458204
rect 279568 458232 279574 458244
rect 280062 458232 280068 458244
rect 279568 458204 280068 458232
rect 279568 458192 279574 458204
rect 280062 458192 280068 458204
rect 280120 458192 280126 458244
rect 43806 456764 43812 456816
rect 43864 456804 43870 456816
rect 60734 456804 60740 456816
rect 43864 456776 60740 456804
rect 43864 456764 43870 456776
rect 60734 456764 60740 456776
rect 60792 456764 60798 456816
rect 331858 456764 331864 456816
rect 331916 456804 331922 456816
rect 337654 456804 337660 456816
rect 331916 456776 337660 456804
rect 331916 456764 331922 456776
rect 337654 456764 337660 456776
rect 337712 456764 337718 456816
rect 535730 456764 535736 456816
rect 535788 456804 535794 456816
rect 543918 456804 543924 456816
rect 535788 456776 543924 456804
rect 535788 456764 535794 456776
rect 543918 456764 543924 456776
rect 543976 456764 543982 456816
rect 556798 456764 556804 456816
rect 556856 456804 556862 456816
rect 580902 456804 580908 456816
rect 556856 456776 580908 456804
rect 556856 456764 556862 456776
rect 580902 456764 580908 456776
rect 580960 456764 580966 456816
rect 265526 456016 265532 456068
rect 265584 456056 265590 456068
rect 327810 456056 327816 456068
rect 265584 456028 327816 456056
rect 265584 456016 265590 456028
rect 327810 456016 327816 456028
rect 327868 456016 327874 456068
rect 245838 455404 245844 455456
rect 245896 455444 245902 455456
rect 264974 455444 264980 455456
rect 245896 455416 264980 455444
rect 245896 455404 245902 455416
rect 264974 455404 264980 455416
rect 265032 455444 265038 455456
rect 265526 455444 265532 455456
rect 265032 455416 265532 455444
rect 265032 455404 265038 455416
rect 265526 455404 265532 455416
rect 265584 455404 265590 455456
rect 245838 454044 245844 454096
rect 245896 454084 245902 454096
rect 308490 454084 308496 454096
rect 245896 454056 308496 454084
rect 245896 454044 245902 454056
rect 308490 454044 308496 454056
rect 308548 454044 308554 454096
rect 330478 454044 330484 454096
rect 330536 454084 330542 454096
rect 337654 454084 337660 454096
rect 330536 454056 337660 454084
rect 330536 454044 330542 454056
rect 337654 454044 337660 454056
rect 337712 454044 337718 454096
rect 535730 452616 535736 452668
rect 535788 452656 535794 452668
rect 541066 452656 541072 452668
rect 535788 452628 541072 452656
rect 535788 452616 535794 452628
rect 541066 452616 541072 452628
rect 541124 452616 541130 452668
rect 327810 451868 327816 451920
rect 327868 451908 327874 451920
rect 337562 451908 337568 451920
rect 327868 451880 337568 451908
rect 327868 451868 327874 451880
rect 337562 451868 337568 451880
rect 337620 451868 337626 451920
rect 34422 451256 34428 451308
rect 34480 451296 34486 451308
rect 60734 451296 60740 451308
rect 34480 451268 60740 451296
rect 34480 451256 34486 451268
rect 60734 451256 60740 451268
rect 60792 451256 60798 451308
rect 52178 450508 52184 450560
rect 52236 450548 52242 450560
rect 59998 450548 60004 450560
rect 52236 450520 60004 450548
rect 52236 450508 52242 450520
rect 59998 450508 60004 450520
rect 60056 450508 60062 450560
rect 254578 449896 254584 449948
rect 254636 449936 254642 449948
rect 337286 449936 337292 449948
rect 254636 449908 337292 449936
rect 254636 449896 254642 449908
rect 337286 449896 337292 449908
rect 337344 449896 337350 449948
rect 3418 449556 3424 449608
rect 3476 449596 3482 449608
rect 8938 449596 8944 449608
rect 3476 449568 8944 449596
rect 3476 449556 3482 449568
rect 8938 449556 8944 449568
rect 8996 449556 9002 449608
rect 60366 448536 60372 448588
rect 60424 448576 60430 448588
rect 61470 448576 61476 448588
rect 60424 448548 61476 448576
rect 60424 448536 60430 448548
rect 61470 448536 61476 448548
rect 61528 448536 61534 448588
rect 535730 447108 535736 447160
rect 535788 447148 535794 447160
rect 542538 447148 542544 447160
rect 535788 447120 542544 447148
rect 535788 447108 535794 447120
rect 542538 447108 542544 447120
rect 542596 447108 542602 447160
rect 305730 446360 305736 446412
rect 305788 446400 305794 446412
rect 337102 446400 337108 446412
rect 305788 446372 337108 446400
rect 305788 446360 305794 446372
rect 337102 446360 337108 446372
rect 337160 446360 337166 446412
rect 245838 445748 245844 445800
rect 245896 445788 245902 445800
rect 261570 445788 261576 445800
rect 245896 445760 261576 445788
rect 245896 445748 245902 445760
rect 261570 445748 261576 445760
rect 261628 445788 261634 445800
rect 265618 445788 265624 445800
rect 261628 445760 265624 445788
rect 261628 445748 261634 445760
rect 265618 445748 265624 445760
rect 265676 445748 265682 445800
rect 42610 444388 42616 444440
rect 42668 444428 42674 444440
rect 60734 444428 60740 444440
rect 42668 444400 60740 444428
rect 42668 444388 42674 444400
rect 60734 444388 60740 444400
rect 60792 444388 60798 444440
rect 535730 444388 535736 444440
rect 535788 444428 535794 444440
rect 550818 444428 550824 444440
rect 535788 444400 550824 444428
rect 535788 444388 535794 444400
rect 550818 444388 550824 444400
rect 550876 444388 550882 444440
rect 336090 443096 336096 443148
rect 336148 443136 336154 443148
rect 338022 443136 338028 443148
rect 336148 443108 338028 443136
rect 336148 443096 336154 443108
rect 338022 443096 338028 443108
rect 338080 443096 338086 443148
rect 46566 441600 46572 441652
rect 46624 441640 46630 441652
rect 60734 441640 60740 441652
rect 46624 441612 60740 441640
rect 46624 441600 46630 441612
rect 60734 441600 60740 441612
rect 60792 441600 60798 441652
rect 535730 441600 535736 441652
rect 535788 441640 535794 441652
rect 548150 441640 548156 441652
rect 535788 441612 548156 441640
rect 535788 441600 535794 441612
rect 548150 441600 548156 441612
rect 548208 441600 548214 441652
rect 245838 438880 245844 438932
rect 245896 438920 245902 438932
rect 283650 438920 283656 438932
rect 245896 438892 283656 438920
rect 245896 438880 245902 438892
rect 283650 438880 283656 438892
rect 283708 438880 283714 438932
rect 329190 438880 329196 438932
rect 329248 438920 329254 438932
rect 337286 438920 337292 438932
rect 329248 438892 337292 438920
rect 329248 438880 329254 438892
rect 337286 438880 337292 438892
rect 337344 438880 337350 438932
rect 247770 436092 247776 436144
rect 247828 436132 247834 436144
rect 337286 436132 337292 436144
rect 247828 436104 337292 436132
rect 247828 436092 247834 436104
rect 337286 436092 337292 436104
rect 337344 436092 337350 436144
rect 245746 434732 245752 434784
rect 245804 434772 245810 434784
rect 322198 434772 322204 434784
rect 245804 434744 322204 434772
rect 245804 434732 245810 434744
rect 322198 434732 322204 434744
rect 322256 434732 322262 434784
rect 535730 434732 535736 434784
rect 535788 434772 535794 434784
rect 546678 434772 546684 434784
rect 535788 434744 546684 434772
rect 535788 434732 535794 434744
rect 546678 434732 546684 434744
rect 546736 434732 546742 434784
rect 288618 433236 288624 433288
rect 288676 433276 288682 433288
rect 289078 433276 289084 433288
rect 288676 433248 289084 433276
rect 288676 433236 288682 433248
rect 289078 433236 289084 433248
rect 289136 433236 289142 433288
rect 245838 432556 245844 432608
rect 245896 432596 245902 432608
rect 288618 432596 288624 432608
rect 245896 432568 288624 432596
rect 245896 432556 245902 432568
rect 288618 432556 288624 432568
rect 288676 432556 288682 432608
rect 253290 431944 253296 431996
rect 253348 431984 253354 431996
rect 317506 431984 317512 431996
rect 253348 431956 317512 431984
rect 253348 431944 253354 431956
rect 317506 431944 317512 431956
rect 317564 431984 317570 431996
rect 337654 431984 337660 431996
rect 317564 431956 337660 431984
rect 317564 431944 317570 431956
rect 337654 431944 337660 431956
rect 337712 431944 337718 431996
rect 288618 431332 288624 431384
rect 288676 431372 288682 431384
rect 293034 431372 293040 431384
rect 288676 431344 293040 431372
rect 288676 431332 288682 431344
rect 293034 431332 293040 431344
rect 293092 431332 293098 431384
rect 326522 431196 326528 431248
rect 326580 431236 326586 431248
rect 337378 431236 337384 431248
rect 326580 431208 337384 431236
rect 326580 431196 326586 431208
rect 337378 431196 337384 431208
rect 337436 431196 337442 431248
rect 548518 431196 548524 431248
rect 548576 431236 548582 431248
rect 571242 431236 571248 431248
rect 548576 431208 571248 431236
rect 548576 431196 548582 431208
rect 571242 431196 571248 431208
rect 571300 431196 571306 431248
rect 53466 430584 53472 430636
rect 53524 430624 53530 430636
rect 60734 430624 60740 430636
rect 53524 430596 60740 430624
rect 53524 430584 53530 430596
rect 60734 430584 60740 430596
rect 60792 430584 60798 430636
rect 570598 429836 570604 429888
rect 570656 429876 570662 429888
rect 571242 429876 571248 429888
rect 570656 429848 571248 429876
rect 570656 429836 570662 429848
rect 571242 429836 571248 429848
rect 571300 429876 571306 429888
rect 580166 429876 580172 429888
rect 571300 429848 580172 429876
rect 571300 429836 571306 429848
rect 580166 429836 580172 429848
rect 580224 429836 580230 429888
rect 282822 429156 282828 429208
rect 282880 429196 282886 429208
rect 336918 429196 336924 429208
rect 282880 429168 336924 429196
rect 282880 429156 282886 429168
rect 336918 429156 336924 429168
rect 336976 429156 336982 429208
rect 4798 428408 4804 428460
rect 4856 428448 4862 428460
rect 51074 428448 51080 428460
rect 4856 428420 51080 428448
rect 4856 428408 4862 428420
rect 51074 428408 51080 428420
rect 51132 428408 51138 428460
rect 51074 427796 51080 427848
rect 51132 427836 51138 427848
rect 52086 427836 52092 427848
rect 51132 427808 52092 427836
rect 51132 427796 51138 427808
rect 52086 427796 52092 427808
rect 52144 427836 52150 427848
rect 60734 427836 60740 427848
rect 52144 427808 60740 427836
rect 52144 427796 52150 427808
rect 60734 427796 60740 427808
rect 60792 427796 60798 427848
rect 245746 427796 245752 427848
rect 245804 427836 245810 427848
rect 323670 427836 323676 427848
rect 245804 427808 323676 427836
rect 245804 427796 245810 427808
rect 323670 427796 323676 427808
rect 323728 427796 323734 427848
rect 256510 426436 256516 426488
rect 256568 426476 256574 426488
rect 336918 426476 336924 426488
rect 256568 426448 336924 426476
rect 256568 426436 256574 426448
rect 336918 426436 336924 426448
rect 336976 426436 336982 426488
rect 535822 426436 535828 426488
rect 535880 426476 535886 426488
rect 548058 426476 548064 426488
rect 535880 426448 548064 426476
rect 535880 426436 535886 426448
rect 548058 426436 548064 426448
rect 548116 426436 548122 426488
rect 245838 425076 245844 425128
rect 245896 425116 245902 425128
rect 251910 425116 251916 425128
rect 245896 425088 251916 425116
rect 245896 425076 245902 425088
rect 251910 425076 251916 425088
rect 251968 425076 251974 425128
rect 264882 425076 264888 425128
rect 264940 425116 264946 425128
rect 337654 425116 337660 425128
rect 264940 425088 337660 425116
rect 264940 425076 264946 425088
rect 337654 425076 337660 425088
rect 337712 425076 337718 425128
rect 32950 423648 32956 423700
rect 33008 423688 33014 423700
rect 60734 423688 60740 423700
rect 33008 423660 60740 423688
rect 33008 423648 33014 423660
rect 60734 423648 60740 423660
rect 60792 423648 60798 423700
rect 251818 422288 251824 422340
rect 251876 422328 251882 422340
rect 337654 422328 337660 422340
rect 251876 422300 337660 422328
rect 251876 422288 251882 422300
rect 337654 422288 337660 422300
rect 337712 422288 337718 422340
rect 535822 422288 535828 422340
rect 535880 422328 535886 422340
rect 539778 422328 539784 422340
rect 535880 422300 539784 422328
rect 535880 422288 535886 422300
rect 539778 422288 539784 422300
rect 539836 422288 539842 422340
rect 50706 420928 50712 420980
rect 50764 420968 50770 420980
rect 60734 420968 60740 420980
rect 50764 420940 60740 420968
rect 50764 420928 50770 420940
rect 60734 420928 60740 420940
rect 60792 420928 60798 420980
rect 245746 420928 245752 420980
rect 245804 420968 245810 420980
rect 322290 420968 322296 420980
rect 245804 420940 322296 420968
rect 245804 420928 245810 420940
rect 322290 420928 322296 420940
rect 322348 420928 322354 420980
rect 251082 420180 251088 420232
rect 251140 420220 251146 420232
rect 307202 420220 307208 420232
rect 251140 420192 307208 420220
rect 251140 420180 251146 420192
rect 307202 420180 307208 420192
rect 307260 420180 307266 420232
rect 535822 419500 535828 419552
rect 535880 419540 535886 419552
rect 545390 419540 545396 419552
rect 535880 419512 545396 419540
rect 535880 419500 535886 419512
rect 545390 419500 545396 419512
rect 545448 419500 545454 419552
rect 558178 419432 558184 419484
rect 558236 419472 558242 419484
rect 580166 419472 580172 419484
rect 558236 419444 580172 419472
rect 558236 419432 558242 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 535822 417324 535828 417376
rect 535880 417364 535886 417376
rect 539870 417364 539876 417376
rect 535880 417336 539876 417364
rect 535880 417324 535886 417336
rect 539870 417324 539876 417336
rect 539928 417324 539934 417376
rect 4798 416780 4804 416832
rect 4856 416820 4862 416832
rect 61010 416820 61016 416832
rect 4856 416792 61016 416820
rect 4856 416780 4862 416792
rect 61010 416780 61016 416792
rect 61068 416780 61074 416832
rect 245838 415352 245844 415404
rect 245896 415392 245902 415404
rect 253290 415392 253296 415404
rect 245896 415364 253296 415392
rect 245896 415352 245902 415364
rect 253290 415352 253296 415364
rect 253348 415352 253354 415404
rect 257338 415352 257344 415404
rect 257396 415392 257402 415404
rect 336826 415392 336832 415404
rect 257396 415364 336832 415392
rect 257396 415352 257402 415364
rect 336826 415352 336832 415364
rect 336884 415352 336890 415404
rect 46750 413992 46756 414044
rect 46808 414032 46814 414044
rect 60826 414032 60832 414044
rect 46808 414004 60832 414032
rect 46808 413992 46814 414004
rect 60826 413992 60832 414004
rect 60884 413992 60890 414044
rect 535822 413992 535828 414044
rect 535880 414032 535886 414044
rect 563054 414032 563060 414044
rect 535880 414004 563060 414032
rect 535880 413992 535886 414004
rect 563054 413992 563060 414004
rect 563112 413992 563118 414044
rect 307662 411884 307668 411936
rect 307720 411924 307726 411936
rect 318058 411924 318064 411936
rect 307720 411896 318064 411924
rect 307720 411884 307726 411896
rect 318058 411884 318064 411896
rect 318116 411884 318122 411936
rect 307202 411380 307208 411392
rect 296686 411352 307208 411380
rect 58986 411272 58992 411324
rect 59044 411312 59050 411324
rect 61378 411312 61384 411324
rect 59044 411284 61384 411312
rect 59044 411272 59050 411284
rect 61378 411272 61384 411284
rect 61436 411272 61442 411324
rect 245838 411272 245844 411324
rect 245896 411312 245902 411324
rect 296686 411312 296714 411352
rect 307202 411340 307208 411352
rect 307260 411380 307266 411392
rect 307662 411380 307668 411392
rect 307260 411352 307668 411380
rect 307260 411340 307266 411352
rect 307662 411340 307668 411352
rect 307720 411340 307726 411392
rect 245896 411284 296714 411312
rect 245896 411272 245902 411284
rect 306558 411272 306564 411324
rect 306616 411312 306622 411324
rect 320818 411312 320824 411324
rect 306616 411284 320824 411312
rect 306616 411272 306622 411284
rect 320818 411272 320824 411284
rect 320876 411272 320882 411324
rect 535822 411272 535828 411324
rect 535880 411312 535886 411324
rect 541158 411312 541164 411324
rect 535880 411284 541164 411312
rect 535880 411272 535886 411284
rect 541158 411272 541164 411284
rect 541216 411272 541222 411324
rect 25682 410524 25688 410576
rect 25740 410564 25746 410576
rect 50338 410564 50344 410576
rect 25740 410536 50344 410564
rect 25740 410524 25746 410536
rect 50338 410524 50344 410536
rect 50396 410524 50402 410576
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 25682 409884 25688 409896
rect 3200 409856 25688 409884
rect 3200 409844 3206 409856
rect 25682 409844 25688 409856
rect 25740 409884 25746 409896
rect 26142 409884 26148 409896
rect 25740 409856 26148 409884
rect 25740 409844 25746 409856
rect 26142 409844 26148 409856
rect 26200 409844 26206 409896
rect 271138 409844 271144 409896
rect 271196 409884 271202 409896
rect 337470 409884 337476 409896
rect 271196 409856 337476 409884
rect 271196 409844 271202 409856
rect 337470 409844 337476 409856
rect 337528 409844 337534 409896
rect 245838 409096 245844 409148
rect 245896 409136 245902 409148
rect 269114 409136 269120 409148
rect 245896 409108 269120 409136
rect 245896 409096 245902 409108
rect 269114 409096 269120 409108
rect 269172 409136 269178 409148
rect 269758 409136 269764 409148
rect 269172 409108 269764 409136
rect 269172 409096 269178 409108
rect 269758 409096 269764 409108
rect 269816 409096 269822 409148
rect 335354 408484 335360 408536
rect 335412 408524 335418 408536
rect 336918 408524 336924 408536
rect 335412 408496 336924 408524
rect 335412 408484 335418 408496
rect 336918 408484 336924 408496
rect 336976 408484 336982 408536
rect 53742 407736 53748 407788
rect 53800 407776 53806 407788
rect 60734 407776 60740 407788
rect 53800 407748 60740 407776
rect 53800 407736 53806 407748
rect 60734 407736 60740 407748
rect 60792 407736 60798 407788
rect 300302 407124 300308 407176
rect 300360 407164 300366 407176
rect 335170 407164 335176 407176
rect 300360 407136 335176 407164
rect 300360 407124 300366 407136
rect 335170 407124 335176 407136
rect 335228 407164 335234 407176
rect 337654 407164 337660 407176
rect 335228 407136 337660 407164
rect 335228 407124 335234 407136
rect 337654 407124 337660 407136
rect 337712 407124 337718 407176
rect 245838 406376 245844 406428
rect 245896 406416 245902 406428
rect 306558 406416 306564 406428
rect 245896 406388 306564 406416
rect 245896 406376 245902 406388
rect 306558 406376 306564 406388
rect 306616 406376 306622 406428
rect 554038 406376 554044 406428
rect 554096 406416 554102 406428
rect 576854 406416 576860 406428
rect 554096 406388 576860 406416
rect 554096 406376 554102 406388
rect 576854 406376 576860 406388
rect 576912 406376 576918 406428
rect 328454 405628 328460 405680
rect 328512 405668 328518 405680
rect 329282 405668 329288 405680
rect 328512 405640 329288 405668
rect 328512 405628 328518 405640
rect 329282 405628 329288 405640
rect 329340 405628 329346 405680
rect 333974 405628 333980 405680
rect 334032 405668 334038 405680
rect 335354 405668 335360 405680
rect 334032 405640 335360 405668
rect 334032 405628 334038 405640
rect 335354 405628 335360 405640
rect 335412 405628 335418 405680
rect 57698 405016 57704 405068
rect 57756 405056 57762 405068
rect 68278 405056 68284 405068
rect 57756 405028 68284 405056
rect 57756 405016 57762 405028
rect 68278 405016 68284 405028
rect 68336 405016 68342 405068
rect 159358 405016 159364 405068
rect 159416 405056 159422 405068
rect 271138 405056 271144 405068
rect 159416 405028 271144 405056
rect 159416 405016 159422 405028
rect 271138 405016 271144 405028
rect 271196 405016 271202 405068
rect 61930 404948 61936 405000
rect 61988 404988 61994 405000
rect 328454 404988 328460 405000
rect 61988 404960 328460 404988
rect 61988 404948 61994 404960
rect 328454 404948 328460 404960
rect 328512 404948 328518 405000
rect 574738 404948 574744 405000
rect 574796 404988 574802 405000
rect 576854 404988 576860 405000
rect 574796 404960 576860 404988
rect 574796 404948 574802 404960
rect 576854 404948 576860 404960
rect 576912 404988 576918 405000
rect 579706 404988 579712 405000
rect 576912 404960 579712 404988
rect 576912 404948 576918 404960
rect 579706 404948 579712 404960
rect 579764 404948 579770 405000
rect 4062 404472 4068 404524
rect 4120 404512 4126 404524
rect 9582 404512 9588 404524
rect 4120 404484 9588 404512
rect 4120 404472 4126 404484
rect 9582 404472 9588 404484
rect 9640 404512 9646 404524
rect 75914 404512 75920 404524
rect 9640 404484 75920 404512
rect 9640 404472 9646 404484
rect 75914 404472 75920 404484
rect 75972 404472 75978 404524
rect 50430 404404 50436 404456
rect 50488 404444 50494 404456
rect 178034 404444 178040 404456
rect 50488 404416 178040 404444
rect 50488 404404 50494 404416
rect 178034 404404 178040 404416
rect 178092 404404 178098 404456
rect 201402 404404 201408 404456
rect 201460 404444 201466 404456
rect 249058 404444 249064 404456
rect 201460 404416 249064 404444
rect 201460 404404 201466 404416
rect 249058 404404 249064 404416
rect 249116 404404 249122 404456
rect 46198 404336 46204 404388
rect 46256 404376 46262 404388
rect 117958 404376 117964 404388
rect 46256 404348 117964 404376
rect 46256 404336 46262 404348
rect 117958 404336 117964 404348
rect 118016 404376 118022 404388
rect 120718 404376 120724 404388
rect 118016 404348 120724 404376
rect 118016 404336 118022 404348
rect 120718 404336 120724 404348
rect 120776 404336 120782 404388
rect 171594 404336 171600 404388
rect 171652 404376 171658 404388
rect 333974 404376 333980 404388
rect 171652 404348 333980 404376
rect 171652 404336 171658 404348
rect 333974 404336 333980 404348
rect 334032 404336 334038 404388
rect 334802 404336 334808 404388
rect 334860 404376 334866 404388
rect 337746 404376 337752 404388
rect 334860 404348 337752 404376
rect 334860 404336 334866 404348
rect 337746 404336 337752 404348
rect 337804 404336 337810 404388
rect 535454 404336 535460 404388
rect 535512 404376 535518 404388
rect 542354 404376 542360 404388
rect 535512 404348 542360 404376
rect 535512 404336 535518 404348
rect 542354 404336 542360 404348
rect 542412 404336 542418 404388
rect 22738 404268 22744 404320
rect 22796 404308 22802 404320
rect 241790 404308 241796 404320
rect 22796 404280 241796 404308
rect 22796 404268 22802 404280
rect 241790 404268 241796 404280
rect 241848 404268 241854 404320
rect 48958 404200 48964 404252
rect 49016 404240 49022 404252
rect 200574 404240 200580 404252
rect 49016 404212 200580 404240
rect 49016 404200 49022 404212
rect 200574 404200 200580 404212
rect 200632 404240 200638 404252
rect 201402 404240 201408 404252
rect 200632 404212 201408 404240
rect 200632 404200 200638 404212
rect 201402 404200 201408 404212
rect 201460 404200 201466 404252
rect 241790 404064 241796 404116
rect 241848 404104 241854 404116
rect 242802 404104 242808 404116
rect 241848 404076 242808 404104
rect 241848 404064 241854 404076
rect 242802 404064 242808 404076
rect 242860 404064 242866 404116
rect 232498 403792 232504 403844
rect 232556 403832 232562 403844
rect 249794 403832 249800 403844
rect 232556 403804 249800 403832
rect 232556 403792 232562 403804
rect 249794 403792 249800 403804
rect 249852 403792 249858 403844
rect 168282 403724 168288 403776
rect 168340 403764 168346 403776
rect 253934 403764 253940 403776
rect 168340 403736 253940 403764
rect 168340 403724 168346 403736
rect 253934 403724 253940 403736
rect 253992 403724 253998 403776
rect 56226 403656 56232 403708
rect 56284 403696 56290 403708
rect 66898 403696 66904 403708
rect 56284 403668 66904 403696
rect 56284 403656 56290 403668
rect 66898 403656 66904 403668
rect 66956 403656 66962 403708
rect 232130 403656 232136 403708
rect 232188 403696 232194 403708
rect 339126 403696 339132 403708
rect 232188 403668 339132 403696
rect 232188 403656 232194 403668
rect 339126 403656 339132 403668
rect 339184 403656 339190 403708
rect 56318 403588 56324 403640
rect 56376 403628 56382 403640
rect 104158 403628 104164 403640
rect 56376 403600 104164 403628
rect 56376 403588 56382 403600
rect 104158 403588 104164 403600
rect 104216 403588 104222 403640
rect 169018 403588 169024 403640
rect 169076 403628 169082 403640
rect 194134 403628 194140 403640
rect 169076 403600 194140 403628
rect 169076 403588 169082 403600
rect 194134 403588 194140 403600
rect 194192 403628 194198 403640
rect 338574 403628 338580 403640
rect 194192 403600 338580 403628
rect 194192 403588 194198 403600
rect 338574 403588 338580 403600
rect 338632 403588 338638 403640
rect 252462 402976 252468 403028
rect 252520 403016 252526 403028
rect 298094 403016 298100 403028
rect 252520 402988 298100 403016
rect 252520 402976 252526 402988
rect 298094 402976 298100 402988
rect 298152 402976 298158 403028
rect 75914 402908 75920 402960
rect 75972 402948 75978 402960
rect 181438 402948 181444 402960
rect 75972 402920 181444 402948
rect 75972 402908 75978 402920
rect 181438 402908 181444 402920
rect 181496 402908 181502 402960
rect 219342 402908 219348 402960
rect 219400 402948 219406 402960
rect 247034 402948 247040 402960
rect 219400 402920 247040 402948
rect 219400 402908 219406 402920
rect 247034 402908 247040 402920
rect 247092 402948 247098 402960
rect 323578 402948 323584 402960
rect 247092 402920 323584 402948
rect 247092 402908 247098 402920
rect 323578 402908 323584 402920
rect 323636 402908 323642 402960
rect 18598 402840 18604 402892
rect 18656 402880 18662 402892
rect 79318 402880 79324 402892
rect 18656 402852 79324 402880
rect 18656 402840 18662 402852
rect 79318 402840 79324 402852
rect 79376 402840 79382 402892
rect 222470 402840 222476 402892
rect 222528 402880 222534 402892
rect 252462 402880 252468 402892
rect 222528 402852 252468 402880
rect 222528 402840 222534 402852
rect 252462 402840 252468 402852
rect 252520 402840 252526 402892
rect 238662 402772 238668 402824
rect 238720 402812 238726 402824
rect 253198 402812 253204 402824
rect 238720 402784 253204 402812
rect 238720 402772 238726 402784
rect 253198 402772 253204 402784
rect 253256 402772 253262 402824
rect 52270 402432 52276 402484
rect 52328 402472 52334 402484
rect 73798 402472 73804 402484
rect 52328 402444 73804 402472
rect 52328 402432 52334 402444
rect 73798 402432 73804 402444
rect 73856 402432 73862 402484
rect 60550 402364 60556 402416
rect 60608 402404 60614 402416
rect 82814 402404 82820 402416
rect 60608 402376 82820 402404
rect 60608 402364 60614 402376
rect 82814 402364 82820 402376
rect 82872 402364 82878 402416
rect 48130 402296 48136 402348
rect 48188 402336 48194 402348
rect 83458 402336 83464 402348
rect 48188 402308 83464 402336
rect 48188 402296 48194 402308
rect 83458 402296 83464 402308
rect 83516 402296 83522 402348
rect 117498 402296 117504 402348
rect 117556 402336 117562 402348
rect 144914 402336 144920 402348
rect 117556 402308 144920 402336
rect 117556 402296 117562 402308
rect 144914 402296 144920 402308
rect 144972 402296 144978 402348
rect 172422 402296 172428 402348
rect 172480 402336 172486 402348
rect 187694 402336 187700 402348
rect 172480 402308 187700 402336
rect 172480 402296 172486 402308
rect 187694 402296 187700 402308
rect 187752 402296 187758 402348
rect 57606 402228 57612 402280
rect 57664 402268 57670 402280
rect 121454 402268 121460 402280
rect 57664 402240 121460 402268
rect 57664 402228 57670 402240
rect 121454 402228 121460 402240
rect 121512 402228 121518 402280
rect 130378 402228 130384 402280
rect 130436 402268 130442 402280
rect 135898 402268 135904 402280
rect 130436 402240 135904 402268
rect 130436 402228 130442 402240
rect 135898 402228 135904 402240
rect 135956 402228 135962 402280
rect 155862 402228 155868 402280
rect 155920 402268 155926 402280
rect 190914 402268 190920 402280
rect 155920 402240 190920 402268
rect 155920 402228 155926 402240
rect 190914 402228 190920 402240
rect 190972 402228 190978 402280
rect 191742 402228 191748 402280
rect 191800 402268 191806 402280
rect 248506 402268 248512 402280
rect 191800 402240 248512 402268
rect 191800 402228 191806 402240
rect 248506 402228 248512 402240
rect 248564 402228 248570 402280
rect 146478 402024 146484 402076
rect 146536 402064 146542 402076
rect 147674 402064 147680 402076
rect 146536 402036 147680 402064
rect 146536 402024 146542 402036
rect 147674 402024 147680 402036
rect 147732 402024 147738 402076
rect 102778 401616 102784 401668
rect 102836 401656 102842 401668
rect 105262 401656 105268 401668
rect 102836 401628 105268 401656
rect 102836 401616 102842 401628
rect 105262 401616 105268 401628
rect 105320 401616 105326 401668
rect 129642 401616 129648 401668
rect 129700 401656 129706 401668
rect 130378 401656 130384 401668
rect 129700 401628 130384 401656
rect 129700 401616 129706 401628
rect 130378 401616 130384 401628
rect 130436 401616 130442 401668
rect 157978 401616 157984 401668
rect 158036 401656 158042 401668
rect 158714 401656 158720 401668
rect 158036 401628 158720 401656
rect 158036 401616 158042 401628
rect 158714 401616 158720 401628
rect 158772 401616 158778 401668
rect 535822 401616 535828 401668
rect 535880 401656 535886 401668
rect 541250 401656 541256 401668
rect 535880 401628 541256 401656
rect 535880 401616 535886 401628
rect 541250 401616 541256 401628
rect 541308 401616 541314 401668
rect 63126 401004 63132 401056
rect 63184 401044 63190 401056
rect 71130 401044 71136 401056
rect 63184 401016 71136 401044
rect 63184 401004 63190 401016
rect 71130 401004 71136 401016
rect 71188 401004 71194 401056
rect 53558 400936 53564 400988
rect 53616 400976 53622 400988
rect 86218 400976 86224 400988
rect 53616 400948 86224 400976
rect 53616 400936 53622 400948
rect 86218 400936 86224 400948
rect 86276 400936 86282 400988
rect 119338 400936 119344 400988
rect 119396 400976 119402 400988
rect 251174 400976 251180 400988
rect 119396 400948 251180 400976
rect 119396 400936 119402 400948
rect 251174 400936 251180 400948
rect 251232 400936 251238 400988
rect 50890 400868 50896 400920
rect 50948 400908 50954 400920
rect 76282 400908 76288 400920
rect 50948 400880 76288 400908
rect 50948 400868 50954 400880
rect 76282 400868 76288 400880
rect 76340 400908 76346 400920
rect 339862 400908 339868 400920
rect 76340 400880 339868 400908
rect 76340 400868 76346 400880
rect 339862 400868 339868 400880
rect 339920 400868 339926 400920
rect 533982 400596 533988 400648
rect 534040 400636 534046 400648
rect 538306 400636 538312 400648
rect 534040 400608 538312 400636
rect 534040 400596 534046 400608
rect 538306 400596 538312 400608
rect 538364 400596 538370 400648
rect 339494 399780 339500 399832
rect 339552 399820 339558 399832
rect 340000 399820 340006 399832
rect 339552 399792 340006 399820
rect 339552 399780 339558 399792
rect 340000 399780 340006 399792
rect 340058 399780 340064 399832
rect 347866 399780 347872 399832
rect 347924 399820 347930 399832
rect 349016 399820 349022 399832
rect 347924 399792 349022 399820
rect 347924 399780 347930 399792
rect 349016 399780 349022 399792
rect 349074 399780 349080 399832
rect 357434 399780 357440 399832
rect 357492 399820 357498 399832
rect 358676 399820 358682 399832
rect 357492 399792 358682 399820
rect 357492 399780 357498 399792
rect 358676 399780 358682 399792
rect 358734 399780 358740 399832
rect 367094 399780 367100 399832
rect 367152 399820 367158 399832
rect 368336 399820 368342 399832
rect 367152 399792 368342 399820
rect 367152 399780 367158 399792
rect 368336 399780 368342 399792
rect 368394 399780 368400 399832
rect 386414 399780 386420 399832
rect 386472 399820 386478 399832
rect 387656 399820 387662 399832
rect 386472 399792 387662 399820
rect 386472 399780 386478 399792
rect 387656 399780 387662 399792
rect 387714 399780 387720 399832
rect 396074 399780 396080 399832
rect 396132 399820 396138 399832
rect 397316 399820 397322 399832
rect 396132 399792 397322 399820
rect 396132 399780 396138 399792
rect 397316 399780 397322 399792
rect 397374 399780 397380 399832
rect 405734 399780 405740 399832
rect 405792 399820 405798 399832
rect 406976 399820 406982 399832
rect 405792 399792 406982 399820
rect 405792 399780 405798 399792
rect 406976 399780 406982 399792
rect 407034 399780 407040 399832
rect 474734 399780 474740 399832
rect 474792 399820 474798 399832
rect 475884 399820 475890 399832
rect 474792 399792 475890 399820
rect 474792 399780 474798 399792
rect 475884 399780 475890 399792
rect 475942 399780 475948 399832
rect 494054 399780 494060 399832
rect 494112 399820 494118 399832
rect 495204 399820 495210 399832
rect 494112 399792 495210 399820
rect 494112 399780 494118 399792
rect 495204 399780 495210 399792
rect 495262 399780 495268 399832
rect 503714 399780 503720 399832
rect 503772 399820 503778 399832
rect 504864 399820 504870 399832
rect 503772 399792 504870 399820
rect 503772 399780 503778 399792
rect 504864 399780 504870 399792
rect 504922 399780 504928 399832
rect 513374 399780 513380 399832
rect 513432 399820 513438 399832
rect 514524 399820 514530 399832
rect 513432 399792 514530 399820
rect 513432 399780 513438 399792
rect 514524 399780 514530 399792
rect 514582 399780 514588 399832
rect 523034 399780 523040 399832
rect 523092 399820 523098 399832
rect 524184 399820 524190 399832
rect 523092 399792 524190 399820
rect 523092 399780 523098 399792
rect 524184 399780 524190 399792
rect 524242 399780 524248 399832
rect 339126 399576 339132 399628
rect 339184 399616 339190 399628
rect 359274 399616 359280 399628
rect 339184 399588 359280 399616
rect 339184 399576 339190 399588
rect 359274 399576 359280 399588
rect 359332 399576 359338 399628
rect 45462 399508 45468 399560
rect 45520 399548 45526 399560
rect 75914 399548 75920 399560
rect 45520 399520 75920 399548
rect 45520 399508 45526 399520
rect 75914 399508 75920 399520
rect 75972 399508 75978 399560
rect 132402 399508 132408 399560
rect 132460 399548 132466 399560
rect 246298 399548 246304 399560
rect 132460 399520 246304 399548
rect 132460 399508 132466 399520
rect 246298 399508 246304 399520
rect 246356 399508 246362 399560
rect 325142 399508 325148 399560
rect 325200 399548 325206 399560
rect 368382 399548 368388 399560
rect 325200 399520 368388 399548
rect 325200 399508 325206 399520
rect 368382 399508 368388 399520
rect 368440 399508 368446 399560
rect 38470 399440 38476 399492
rect 38528 399480 38534 399492
rect 71038 399480 71044 399492
rect 38528 399452 71044 399480
rect 38528 399440 38534 399452
rect 71038 399440 71044 399452
rect 71096 399440 71102 399492
rect 111058 399440 111064 399492
rect 111116 399480 111122 399492
rect 126974 399480 126980 399492
rect 111116 399452 126980 399480
rect 111116 399440 111122 399452
rect 126974 399440 126980 399452
rect 127032 399440 127038 399492
rect 151078 399440 151084 399492
rect 151136 399480 151142 399492
rect 174814 399480 174820 399492
rect 151136 399452 174820 399480
rect 151136 399440 151142 399452
rect 174814 399440 174820 399452
rect 174872 399480 174878 399492
rect 380618 399480 380624 399492
rect 174872 399452 380624 399480
rect 174872 399440 174878 399452
rect 380618 399440 380624 399452
rect 380676 399440 380682 399492
rect 526438 399440 526444 399492
rect 526496 399480 526502 399492
rect 543918 399480 543924 399492
rect 526496 399452 543924 399480
rect 526496 399440 526502 399452
rect 543918 399440 543924 399452
rect 543976 399440 543982 399492
rect 368382 398964 368388 399016
rect 368440 399004 368446 399016
rect 428182 399004 428188 399016
rect 368440 398976 428188 399004
rect 368440 398964 368446 398976
rect 428182 398964 428188 398976
rect 428240 398964 428246 399016
rect 168374 398896 168380 398948
rect 168432 398936 168438 398948
rect 169754 398936 169760 398948
rect 168432 398908 169760 398936
rect 168432 398896 168438 398908
rect 169754 398896 169760 398908
rect 169812 398896 169818 398948
rect 242802 398896 242808 398948
rect 242860 398936 242866 398948
rect 440326 398936 440332 398948
rect 242860 398908 440332 398936
rect 242860 398896 242866 398908
rect 440326 398896 440332 398908
rect 440384 398896 440390 398948
rect 64690 398828 64696 398880
rect 64748 398868 64754 398880
rect 339494 398868 339500 398880
rect 64748 398840 339500 398868
rect 64748 398828 64754 398840
rect 339494 398828 339500 398840
rect 339552 398828 339558 398880
rect 358814 398828 358820 398880
rect 358872 398868 358878 398880
rect 359274 398868 359280 398880
rect 358872 398840 359280 398868
rect 358872 398828 358878 398840
rect 359274 398828 359280 398840
rect 359332 398868 359338 398880
rect 533430 398868 533436 398880
rect 359332 398840 533436 398868
rect 359332 398828 359338 398840
rect 533430 398828 533436 398840
rect 533488 398828 533494 398880
rect 127526 398760 127532 398812
rect 127584 398800 127590 398812
rect 411438 398800 411444 398812
rect 127584 398772 411444 398800
rect 127584 398760 127590 398772
rect 411438 398760 411444 398772
rect 411496 398760 411502 398812
rect 457254 398760 457260 398812
rect 457312 398800 457318 398812
rect 542998 398800 543004 398812
rect 457312 398772 543004 398800
rect 457312 398760 457318 398772
rect 542998 398760 543004 398772
rect 543056 398760 543062 398812
rect 169754 398692 169760 398744
rect 169812 398732 169818 398744
rect 454586 398732 454592 398744
rect 169812 398704 454592 398732
rect 169812 398692 169818 398704
rect 454586 398692 454592 398704
rect 454644 398692 454650 398744
rect 511994 398692 512000 398744
rect 512052 398732 512058 398744
rect 560938 398732 560944 398744
rect 512052 398704 560944 398732
rect 512052 398692 512058 398704
rect 560938 398692 560944 398704
rect 560996 398692 561002 398744
rect 100018 398624 100024 398676
rect 100076 398664 100082 398676
rect 102042 398664 102048 398676
rect 100076 398636 102048 398664
rect 100076 398624 100082 398636
rect 102042 398624 102048 398636
rect 102100 398664 102106 398676
rect 380526 398664 380532 398676
rect 102100 398636 380532 398664
rect 102100 398624 102106 398636
rect 380526 398624 380532 398636
rect 380584 398624 380590 398676
rect 380618 398624 380624 398676
rect 380676 398664 380682 398676
rect 464246 398664 464252 398676
rect 380676 398636 464252 398664
rect 380676 398624 380682 398636
rect 464246 398624 464252 398636
rect 464304 398624 464310 398676
rect 338574 398556 338580 398608
rect 338632 398596 338638 398608
rect 485498 398596 485504 398608
rect 338632 398568 485504 398596
rect 338632 398556 338638 398568
rect 485498 398556 485504 398568
rect 485556 398556 485562 398608
rect 335998 398488 336004 398540
rect 336056 398528 336062 398540
rect 385126 398528 385132 398540
rect 336056 398500 385132 398528
rect 336056 398488 336062 398500
rect 385126 398488 385132 398500
rect 385184 398488 385190 398540
rect 440326 398488 440332 398540
rect 440384 398528 440390 398540
rect 497734 398528 497740 398540
rect 440384 398500 497740 398528
rect 440384 398488 440390 398500
rect 497734 398488 497740 398500
rect 497792 398488 497798 398540
rect 339862 398420 339868 398472
rect 339920 398460 339926 398472
rect 353386 398460 353392 398472
rect 339920 398432 353392 398460
rect 339920 398420 339926 398432
rect 353386 398420 353392 398432
rect 353444 398460 353450 398472
rect 354122 398460 354128 398472
rect 353444 398432 354128 398460
rect 353444 398420 353450 398432
rect 354122 398420 354128 398432
rect 354180 398420 354186 398472
rect 530578 398216 530584 398268
rect 530636 398256 530642 398268
rect 539870 398256 539876 398268
rect 530636 398228 539876 398256
rect 530636 398216 530642 398228
rect 539870 398216 539876 398228
rect 539928 398216 539934 398268
rect 41322 398148 41328 398200
rect 41380 398188 41386 398200
rect 75178 398188 75184 398200
rect 41380 398160 75184 398188
rect 41380 398148 41386 398160
rect 75178 398148 75184 398160
rect 75236 398148 75242 398200
rect 120718 398148 120724 398200
rect 120776 398188 120782 398200
rect 127526 398188 127532 398200
rect 120776 398160 127532 398188
rect 120776 398148 120782 398160
rect 127526 398148 127532 398160
rect 127584 398148 127590 398200
rect 530670 398148 530676 398200
rect 530728 398188 530734 398200
rect 541066 398188 541072 398200
rect 530728 398160 541072 398188
rect 530728 398148 530734 398160
rect 541066 398148 541072 398160
rect 541124 398148 541130 398200
rect 3970 398080 3976 398132
rect 4028 398120 4034 398132
rect 31018 398120 31024 398132
rect 4028 398092 31024 398120
rect 4028 398080 4034 398092
rect 31018 398080 31024 398092
rect 31076 398080 31082 398132
rect 62114 398080 62120 398132
rect 62172 398120 62178 398132
rect 63310 398120 63316 398132
rect 62172 398092 63316 398120
rect 62172 398080 62178 398092
rect 63310 398080 63316 398092
rect 63368 398120 63374 398132
rect 331214 398120 331220 398132
rect 63368 398092 331220 398120
rect 63368 398080 63374 398092
rect 331214 398080 331220 398092
rect 331272 398120 331278 398132
rect 331950 398120 331956 398132
rect 331272 398092 331956 398120
rect 331272 398080 331278 398092
rect 331950 398080 331956 398092
rect 332008 398080 332014 398132
rect 356790 398080 356796 398132
rect 356848 398120 356854 398132
rect 452010 398120 452016 398132
rect 356848 398092 452016 398120
rect 356848 398080 356854 398092
rect 452010 398080 452016 398092
rect 452068 398080 452074 398132
rect 502978 398080 502984 398132
rect 503036 398120 503042 398132
rect 539686 398120 539692 398132
rect 503036 398092 539692 398120
rect 503036 398080 503042 398092
rect 539686 398080 539692 398092
rect 539744 398080 539750 398132
rect 355226 397468 355232 397520
rect 355284 397508 355290 397520
rect 356698 397508 356704 397520
rect 355284 397480 356704 397508
rect 355284 397468 355290 397480
rect 356698 397468 356704 397480
rect 356756 397468 356762 397520
rect 385126 397468 385132 397520
rect 385184 397508 385190 397520
rect 385678 397508 385684 397520
rect 385184 397480 385684 397508
rect 385184 397468 385190 397480
rect 385678 397468 385684 397480
rect 385736 397468 385742 397520
rect 464338 397468 464344 397520
rect 464396 397508 464402 397520
rect 466178 397508 466184 397520
rect 464396 397480 466184 397508
rect 464396 397468 464402 397480
rect 466178 397468 466184 397480
rect 466236 397468 466242 397520
rect 500218 397468 500224 397520
rect 500276 397508 500282 397520
rect 502334 397508 502340 397520
rect 500276 397480 502340 397508
rect 500276 397468 500282 397480
rect 502334 397468 502340 397480
rect 502392 397468 502398 397520
rect 511994 397468 512000 397520
rect 512052 397508 512058 397520
rect 512638 397508 512644 397520
rect 512052 397480 512644 397508
rect 512052 397468 512058 397480
rect 512638 397468 512644 397480
rect 512696 397468 512702 397520
rect 525058 397468 525064 397520
rect 525116 397508 525122 397520
rect 526070 397508 526076 397520
rect 525116 397480 526076 397508
rect 525116 397468 525122 397480
rect 526070 397468 526076 397480
rect 526128 397468 526134 397520
rect 41138 397400 41144 397452
rect 41196 397440 41202 397452
rect 41322 397440 41328 397452
rect 41196 397412 41328 397440
rect 41196 397400 41202 397412
rect 41322 397400 41328 397412
rect 41380 397440 41386 397452
rect 545298 397440 545304 397452
rect 41380 397412 545304 397440
rect 41380 397400 41386 397412
rect 545298 397400 545304 397412
rect 545356 397400 545362 397452
rect 140590 397332 140596 397384
rect 140648 397372 140654 397384
rect 545206 397372 545212 397384
rect 140648 397344 545212 397372
rect 140648 397332 140654 397344
rect 545206 397332 545212 397344
rect 545264 397332 545270 397384
rect 161934 397264 161940 397316
rect 161992 397304 161998 397316
rect 162762 397304 162768 397316
rect 161992 397276 162768 397304
rect 161992 397264 161998 397276
rect 162762 397264 162768 397276
rect 162820 397304 162826 397316
rect 283558 397304 283564 397316
rect 162820 397276 283564 397304
rect 162820 397264 162826 397276
rect 283558 397264 283564 397276
rect 283616 397264 283622 397316
rect 322290 397264 322296 397316
rect 322348 397304 322354 397316
rect 322750 397304 322756 397316
rect 322348 397276 322756 397304
rect 322348 397264 322354 397276
rect 322750 397264 322756 397276
rect 322808 397304 322814 397316
rect 552106 397304 552112 397316
rect 322808 397276 552112 397304
rect 322808 397264 322814 397276
rect 552106 397264 552112 397276
rect 552164 397264 552170 397316
rect 265710 397196 265716 397248
rect 265768 397236 265774 397248
rect 331306 397236 331312 397248
rect 265768 397208 331312 397236
rect 265768 397196 265774 397208
rect 331306 397196 331312 397208
rect 331364 397196 331370 397248
rect 54938 396856 54944 396908
rect 54996 396896 55002 396908
rect 89714 396896 89720 396908
rect 54996 396868 89720 396896
rect 54996 396856 55002 396868
rect 89714 396856 89720 396868
rect 89772 396856 89778 396908
rect 335262 396856 335268 396908
rect 335320 396896 335326 396908
rect 347774 396896 347780 396908
rect 335320 396868 347780 396896
rect 335320 396856 335326 396868
rect 347774 396856 347780 396868
rect 347832 396856 347838 396908
rect 45462 396788 45468 396840
rect 45520 396828 45526 396840
rect 85942 396828 85948 396840
rect 45520 396800 85948 396828
rect 45520 396788 45526 396800
rect 85942 396788 85948 396800
rect 86000 396788 86006 396840
rect 163498 396788 163504 396840
rect 163556 396828 163562 396840
rect 206370 396828 206376 396840
rect 163556 396800 206376 396828
rect 163556 396788 163562 396800
rect 206370 396788 206376 396800
rect 206428 396788 206434 396840
rect 227622 396788 227628 396840
rect 227680 396828 227686 396840
rect 250530 396828 250536 396840
rect 227680 396800 250536 396828
rect 227680 396788 227686 396800
rect 250530 396788 250536 396800
rect 250588 396788 250594 396840
rect 331306 396788 331312 396840
rect 331364 396828 331370 396840
rect 332410 396828 332416 396840
rect 331364 396800 332416 396828
rect 331364 396788 331370 396800
rect 332410 396788 332416 396800
rect 332468 396828 332474 396840
rect 332468 396800 364334 396828
rect 332468 396788 332474 396800
rect 48130 396720 48136 396772
rect 48188 396760 48194 396772
rect 95602 396760 95608 396772
rect 48188 396732 95608 396760
rect 48188 396720 48194 396732
rect 95602 396720 95608 396732
rect 95660 396720 95666 396772
rect 195238 396720 195244 396772
rect 195296 396760 195302 396772
rect 256786 396760 256792 396772
rect 195296 396732 256792 396760
rect 195296 396720 195302 396732
rect 256786 396720 256792 396732
rect 256844 396720 256850 396772
rect 273990 396720 273996 396772
rect 274048 396760 274054 396772
rect 341518 396760 341524 396772
rect 274048 396732 341524 396760
rect 274048 396720 274054 396732
rect 341518 396720 341524 396732
rect 341576 396760 341582 396772
rect 355226 396760 355232 396772
rect 341576 396732 355232 396760
rect 341576 396720 341582 396732
rect 355226 396720 355232 396732
rect 355284 396720 355290 396772
rect 364306 396760 364334 396800
rect 365070 396760 365076 396772
rect 364306 396732 365076 396760
rect 365070 396720 365076 396732
rect 365128 396760 365134 396772
rect 408862 396760 408868 396772
rect 365128 396732 408868 396760
rect 365128 396720 365134 396732
rect 408862 396720 408868 396732
rect 408920 396720 408926 396772
rect 414106 396720 414112 396772
rect 414164 396760 414170 396772
rect 425606 396760 425612 396772
rect 414164 396732 425612 396760
rect 414164 396720 414170 396732
rect 425606 396720 425612 396732
rect 425664 396720 425670 396772
rect 489178 396720 489184 396772
rect 489236 396760 489242 396772
rect 546586 396760 546592 396772
rect 489236 396732 546592 396760
rect 489236 396720 489242 396732
rect 546586 396720 546592 396732
rect 546644 396720 546650 396772
rect 37090 395972 37096 396024
rect 37148 396012 37154 396024
rect 540974 396012 540980 396024
rect 37148 395984 540980 396012
rect 37148 395972 37154 395984
rect 540974 395972 540980 395984
rect 541032 395972 541038 396024
rect 308490 395904 308496 395956
rect 308548 395944 308554 395956
rect 309042 395944 309048 395956
rect 308548 395916 309048 395944
rect 308548 395904 308554 395916
rect 309042 395904 309048 395916
rect 309100 395944 309106 395956
rect 538490 395944 538496 395956
rect 309100 395916 538496 395944
rect 309100 395904 309106 395916
rect 538490 395904 538496 395916
rect 538548 395904 538554 395956
rect 322198 395836 322204 395888
rect 322256 395876 322262 395888
rect 322842 395876 322848 395888
rect 322256 395848 322848 395876
rect 322256 395836 322262 395848
rect 322842 395836 322848 395848
rect 322900 395876 322906 395888
rect 549438 395876 549444 395888
rect 322900 395848 549444 395876
rect 322900 395836 322906 395848
rect 549438 395836 549444 395848
rect 549496 395836 549502 395888
rect 260742 395768 260748 395820
rect 260800 395808 260806 395820
rect 363598 395808 363604 395820
rect 260800 395780 363604 395808
rect 260800 395768 260806 395780
rect 363598 395768 363604 395780
rect 363656 395768 363662 395820
rect 357342 395428 357348 395480
rect 357400 395468 357406 395480
rect 375374 395468 375380 395480
rect 357400 395440 375380 395468
rect 357400 395428 357406 395440
rect 375374 395428 375380 395440
rect 375432 395428 375438 395480
rect 173158 395360 173164 395412
rect 173216 395400 173222 395412
rect 259454 395400 259460 395412
rect 173216 395372 259460 395400
rect 173216 395360 173222 395372
rect 259454 395360 259460 395372
rect 259512 395400 259518 395412
rect 260742 395400 260748 395412
rect 259512 395372 260748 395400
rect 259512 395360 259518 395372
rect 260742 395360 260748 395372
rect 260800 395360 260806 395412
rect 371970 395360 371976 395412
rect 372028 395400 372034 395412
rect 382458 395400 382464 395412
rect 372028 395372 382464 395400
rect 372028 395360 372034 395372
rect 382458 395360 382464 395372
rect 382516 395360 382522 395412
rect 391198 395360 391204 395412
rect 391256 395400 391262 395412
rect 414014 395400 414020 395412
rect 391256 395372 414020 395400
rect 391256 395360 391262 395372
rect 414014 395360 414020 395372
rect 414072 395360 414078 395412
rect 520918 395360 520924 395412
rect 520976 395400 520982 395412
rect 542446 395400 542452 395412
rect 520976 395372 542452 395400
rect 520976 395360 520982 395372
rect 542446 395360 542452 395372
rect 542504 395360 542510 395412
rect 168190 395292 168196 395344
rect 168248 395332 168254 395344
rect 197354 395332 197360 395344
rect 168248 395304 197360 395332
rect 168248 395292 168254 395304
rect 197354 395292 197360 395304
rect 197412 395292 197418 395344
rect 214558 395292 214564 395344
rect 214616 395332 214622 395344
rect 244366 395332 244372 395344
rect 214616 395304 244372 395332
rect 214616 395292 214622 395304
rect 244366 395292 244372 395304
rect 244424 395332 244430 395344
rect 357342 395332 357348 395344
rect 244424 395304 357348 395332
rect 244424 395292 244430 395304
rect 357342 395292 357348 395304
rect 357400 395292 357406 395344
rect 369670 395292 369676 395344
rect 369728 395332 369734 395344
rect 401778 395332 401784 395344
rect 369728 395304 401784 395332
rect 369728 395292 369734 395304
rect 401778 395292 401784 395304
rect 401836 395292 401842 395344
rect 416038 395292 416044 395344
rect 416096 395332 416102 395344
rect 452838 395332 452844 395344
rect 416096 395304 452844 395332
rect 416096 395292 416102 395304
rect 452838 395292 452844 395304
rect 452896 395292 452902 395344
rect 522298 395292 522304 395344
rect 522356 395332 522362 395344
rect 545114 395332 545120 395344
rect 522356 395304 545120 395332
rect 522356 395292 522362 395304
rect 545114 395292 545120 395304
rect 545172 395292 545178 395344
rect 61838 394612 61844 394664
rect 61896 394652 61902 394664
rect 62022 394652 62028 394664
rect 61896 394624 62028 394652
rect 61896 394612 61902 394624
rect 62022 394612 62028 394624
rect 62080 394612 62086 394664
rect 246390 394612 246396 394664
rect 246448 394652 246454 394664
rect 246942 394652 246948 394664
rect 246448 394624 246948 394652
rect 246448 394612 246454 394624
rect 246942 394612 246948 394624
rect 247000 394652 247006 394664
rect 542538 394652 542544 394664
rect 247000 394624 542544 394652
rect 247000 394612 247006 394624
rect 542538 394612 542544 394624
rect 542596 394612 542602 394664
rect 251910 394544 251916 394596
rect 251968 394584 251974 394596
rect 252462 394584 252468 394596
rect 251968 394556 252468 394584
rect 251968 394544 251974 394556
rect 252462 394544 252468 394556
rect 252520 394544 252526 394596
rect 335170 394544 335176 394596
rect 335228 394584 335234 394596
rect 582466 394584 582472 394596
rect 335228 394556 582472 394584
rect 335228 394544 335234 394556
rect 582466 394544 582472 394556
rect 582524 394544 582530 394596
rect 337930 394476 337936 394528
rect 337988 394516 337994 394528
rect 434806 394516 434812 394528
rect 337988 394488 434812 394516
rect 337988 394476 337994 394488
rect 434806 394476 434812 394488
rect 434864 394516 434870 394528
rect 580258 394516 580264 394528
rect 434864 394488 580264 394516
rect 434864 394476 434870 394488
rect 580258 394476 580264 394488
rect 580316 394476 580322 394528
rect 323670 394408 323676 394460
rect 323728 394448 323734 394460
rect 550818 394448 550824 394460
rect 323728 394420 550824 394448
rect 323728 394408 323734 394420
rect 550818 394408 550824 394420
rect 550876 394408 550882 394460
rect 178034 394340 178040 394392
rect 178092 394380 178098 394392
rect 178678 394380 178684 394392
rect 178092 394352 178684 394380
rect 178092 394340 178098 394352
rect 178678 394340 178684 394352
rect 178736 394340 178742 394392
rect 46658 394068 46664 394120
rect 46716 394108 46722 394120
rect 88334 394108 88340 394120
rect 46716 394080 88340 394108
rect 46716 394068 46722 394080
rect 88334 394068 88340 394080
rect 88392 394068 88398 394120
rect 189718 394068 189724 394120
rect 189776 394108 189782 394120
rect 262214 394108 262220 394120
rect 189776 394080 262220 394108
rect 189776 394068 189782 394080
rect 262214 394068 262220 394080
rect 262272 394068 262278 394120
rect 43990 394000 43996 394052
rect 44048 394040 44054 394052
rect 133874 394040 133880 394052
rect 44048 394012 133880 394040
rect 44048 394000 44054 394012
rect 133874 394000 133880 394012
rect 133932 394000 133938 394052
rect 179322 394000 179328 394052
rect 179380 394040 179386 394052
rect 337378 394040 337384 394052
rect 179380 394012 337384 394040
rect 179380 394000 179386 394012
rect 337378 394000 337384 394012
rect 337436 394000 337442 394052
rect 62022 393932 62028 393984
rect 62080 393972 62086 393984
rect 335354 393972 335360 393984
rect 62080 393944 335360 393972
rect 62080 393932 62086 393944
rect 335354 393932 335360 393944
rect 335412 393972 335418 393984
rect 336090 393972 336096 393984
rect 335412 393944 336096 393972
rect 335412 393932 335418 393944
rect 336090 393932 336096 393944
rect 336148 393932 336154 393984
rect 355502 393932 355508 393984
rect 355560 393972 355566 393984
rect 421098 393972 421104 393984
rect 355560 393944 421104 393972
rect 355560 393932 355566 393944
rect 421098 393932 421104 393944
rect 421156 393932 421162 393984
rect 472618 393932 472624 393984
rect 472676 393972 472682 393984
rect 492674 393972 492680 393984
rect 472676 393944 492680 393972
rect 472676 393932 472682 393944
rect 492674 393932 492680 393944
rect 492732 393932 492738 393984
rect 496078 393932 496084 393984
rect 496136 393972 496142 393984
rect 531314 393972 531320 393984
rect 496136 393944 531320 393972
rect 496136 393932 496142 393944
rect 531314 393932 531320 393944
rect 531372 393932 531378 393984
rect 160738 393320 160744 393372
rect 160796 393360 160802 393372
rect 178678 393360 178684 393372
rect 160796 393332 178684 393360
rect 160796 393320 160802 393332
rect 178678 393320 178684 393332
rect 178736 393320 178742 393372
rect 252462 393320 252468 393372
rect 252520 393360 252526 393372
rect 252520 393332 372660 393360
rect 252520 393320 252526 393332
rect 372632 393292 372660 393332
rect 373902 393292 373908 393304
rect 372632 393264 373908 393292
rect 373902 393252 373908 393264
rect 373960 393292 373966 393304
rect 457438 393292 457444 393304
rect 373960 393264 457444 393292
rect 373960 393252 373966 393264
rect 457438 393252 457444 393264
rect 457496 393252 457502 393304
rect 329742 392776 329748 392828
rect 329800 392816 329806 392828
rect 346486 392816 346492 392828
rect 329800 392788 346492 392816
rect 329800 392776 329806 392788
rect 346486 392776 346492 392788
rect 346544 392776 346550 392828
rect 321462 392708 321468 392760
rect 321520 392748 321526 392760
rect 343818 392748 343824 392760
rect 321520 392720 343824 392748
rect 321520 392708 321526 392720
rect 343818 392708 343824 392720
rect 343876 392708 343882 392760
rect 374638 392708 374644 392760
rect 374696 392748 374702 392760
rect 405734 392748 405740 392760
rect 374696 392720 405740 392748
rect 374696 392708 374702 392720
rect 405734 392708 405740 392720
rect 405792 392708 405798 392760
rect 171042 392640 171048 392692
rect 171100 392680 171106 392692
rect 252462 392680 252468 392692
rect 171100 392652 252468 392680
rect 171100 392640 171106 392652
rect 252462 392640 252468 392652
rect 252520 392640 252526 392692
rect 324222 392640 324228 392692
rect 324280 392680 324286 392692
rect 351914 392680 351920 392692
rect 324280 392652 351920 392680
rect 324280 392640 324286 392652
rect 351914 392640 351920 392652
rect 351972 392640 351978 392692
rect 377398 392640 377404 392692
rect 377456 392680 377462 392692
rect 418154 392680 418160 392692
rect 377456 392652 418160 392680
rect 377456 392640 377462 392652
rect 418154 392640 418160 392652
rect 418212 392640 418218 392692
rect 95878 392572 95884 392624
rect 95936 392612 95942 392624
rect 242894 392612 242900 392624
rect 95936 392584 242900 392612
rect 95936 392572 95942 392584
rect 242894 392572 242900 392584
rect 242952 392572 242958 392624
rect 292022 392572 292028 392624
rect 292080 392612 292086 392624
rect 300210 392612 300216 392624
rect 292080 392584 300216 392612
rect 292080 392572 292086 392584
rect 300210 392572 300216 392584
rect 300268 392572 300274 392624
rect 337838 392572 337844 392624
rect 337896 392612 337902 392624
rect 368474 392612 368480 392624
rect 337896 392584 368480 392612
rect 337896 392572 337902 392584
rect 368474 392572 368480 392584
rect 368532 392572 368538 392624
rect 379422 392572 379428 392624
rect 379480 392612 379486 392624
rect 579614 392612 579620 392624
rect 379480 392584 579620 392612
rect 379480 392572 379486 392584
rect 579614 392572 579620 392584
rect 579672 392572 579678 392624
rect 238754 392028 238760 392080
rect 238812 392068 238818 392080
rect 292022 392068 292028 392080
rect 238812 392040 292028 392068
rect 238812 392028 238818 392040
rect 292022 392028 292028 392040
rect 292080 392028 292086 392080
rect 142798 391960 142804 392012
rect 142856 392000 142862 392012
rect 245654 392000 245660 392012
rect 142856 391972 245660 392000
rect 142856 391960 142862 391972
rect 245654 391960 245660 391972
rect 245712 391960 245718 392012
rect 292298 391960 292304 392012
rect 292356 392000 292362 392012
rect 350534 392000 350540 392012
rect 292356 391972 350540 392000
rect 292356 391960 292362 391972
rect 350534 391960 350540 391972
rect 350592 391960 350598 392012
rect 245672 391932 245700 391960
rect 541250 391932 541256 391944
rect 245672 391904 541256 391932
rect 541250 391892 541256 391904
rect 541308 391892 541314 391944
rect 135898 391348 135904 391400
rect 135956 391388 135962 391400
rect 205634 391388 205640 391400
rect 135956 391360 205640 391388
rect 135956 391348 135962 391360
rect 205634 391348 205640 391360
rect 205692 391348 205698 391400
rect 197354 391280 197360 391332
rect 197412 391320 197418 391332
rect 292298 391320 292304 391332
rect 197412 391292 292304 391320
rect 197412 391280 197418 391292
rect 292298 391280 292304 391292
rect 292356 391280 292362 391332
rect 158622 391212 158628 391264
rect 158680 391252 158686 391264
rect 258074 391252 258080 391264
rect 158680 391224 258080 391252
rect 158680 391212 158686 391224
rect 258074 391212 258080 391224
rect 258132 391212 258138 391264
rect 166810 389784 166816 389836
rect 166868 389824 166874 389836
rect 267734 389824 267740 389836
rect 166868 389796 267740 389824
rect 166868 389784 166874 389796
rect 267734 389784 267740 389796
rect 267792 389784 267798 389836
rect 286962 389784 286968 389836
rect 287020 389824 287026 389836
rect 343726 389824 343732 389836
rect 287020 389796 343732 389824
rect 287020 389784 287026 389796
rect 343726 389784 343732 389796
rect 343784 389784 343790 389836
rect 409782 389784 409788 389836
rect 409840 389824 409846 389836
rect 539778 389824 539784 389836
rect 409840 389796 539784 389824
rect 409840 389784 409846 389796
rect 539778 389784 539784 389796
rect 539836 389784 539842 389836
rect 245010 389172 245016 389224
rect 245068 389212 245074 389224
rect 531958 389212 531964 389224
rect 245068 389184 531964 389212
rect 245068 389172 245074 389184
rect 531958 389172 531964 389184
rect 532016 389172 532022 389224
rect 52086 388492 52092 388544
rect 52144 388532 52150 388544
rect 153194 388532 153200 388544
rect 52144 388504 153200 388532
rect 52144 388492 52150 388504
rect 153194 388492 153200 388504
rect 153252 388532 153258 388544
rect 154114 388532 154120 388544
rect 153252 388504 154120 388532
rect 153252 388492 153258 388504
rect 154114 388492 154120 388504
rect 154172 388492 154178 388544
rect 152550 388424 152556 388476
rect 152608 388464 152614 388476
rect 270494 388464 270500 388476
rect 152608 388436 270500 388464
rect 152608 388424 152614 388436
rect 270494 388424 270500 388436
rect 270552 388424 270558 388476
rect 317230 388424 317236 388476
rect 317288 388464 317294 388476
rect 333422 388464 333428 388476
rect 317288 388436 333428 388464
rect 317288 388424 317294 388436
rect 333422 388424 333428 388436
rect 333480 388424 333486 388476
rect 339310 388424 339316 388476
rect 339368 388464 339374 388476
rect 406378 388464 406384 388476
rect 339368 388436 406384 388464
rect 339368 388424 339374 388436
rect 406378 388424 406384 388436
rect 406436 388424 406442 388476
rect 482278 388424 482284 388476
rect 482336 388464 482342 388476
rect 518894 388464 518900 388476
rect 482336 388436 518900 388464
rect 482336 388424 482342 388436
rect 518894 388424 518900 388436
rect 518952 388424 518958 388476
rect 154114 387880 154120 387932
rect 154172 387920 154178 387932
rect 202966 387920 202972 387932
rect 154172 387892 202972 387920
rect 154172 387880 154178 387892
rect 202966 387880 202972 387892
rect 203024 387880 203030 387932
rect 218698 387880 218704 387932
rect 218756 387920 218762 387932
rect 219342 387920 219348 387932
rect 218756 387892 219348 387920
rect 218756 387880 218762 387892
rect 219342 387880 219348 387892
rect 219400 387920 219406 387932
rect 270494 387920 270500 387932
rect 219400 387892 270500 387920
rect 219400 387880 219406 387892
rect 270494 387880 270500 387892
rect 270552 387880 270558 387932
rect 182174 387812 182180 387864
rect 182232 387852 182238 387864
rect 316034 387852 316040 387864
rect 182232 387824 316040 387852
rect 182232 387812 182238 387824
rect 316034 387812 316040 387824
rect 316092 387852 316098 387864
rect 317230 387852 317236 387864
rect 316092 387824 317236 387852
rect 316092 387812 316098 387824
rect 317230 387812 317236 387824
rect 317288 387812 317294 387864
rect 367002 387812 367008 387864
rect 367060 387852 367066 387864
rect 440510 387852 440516 387864
rect 367060 387824 440516 387852
rect 367060 387812 367066 387824
rect 440510 387812 440516 387824
rect 440568 387812 440574 387864
rect 60366 387744 60372 387796
rect 60424 387784 60430 387796
rect 60550 387784 60556 387796
rect 60424 387756 60556 387784
rect 60424 387744 60430 387756
rect 60550 387744 60556 387756
rect 60608 387744 60614 387796
rect 288342 387200 288348 387252
rect 288400 387240 288406 387252
rect 306466 387240 306472 387252
rect 288400 387212 306472 387240
rect 288400 387200 288406 387212
rect 306466 387200 306472 387212
rect 306524 387200 306530 387252
rect 181438 387132 181444 387184
rect 181496 387172 181502 387184
rect 241514 387172 241520 387184
rect 181496 387144 241520 387172
rect 181496 387132 181502 387144
rect 241514 387132 241520 387144
rect 241572 387172 241578 387184
rect 365714 387172 365720 387184
rect 241572 387144 365720 387172
rect 241572 387132 241578 387144
rect 365714 387132 365720 387144
rect 365772 387172 365778 387184
rect 367002 387172 367008 387184
rect 365772 387144 367008 387172
rect 365772 387132 365778 387144
rect 367002 387132 367008 387144
rect 367060 387132 367066 387184
rect 60550 387064 60556 387116
rect 60608 387104 60614 387116
rect 327166 387104 327172 387116
rect 60608 387076 327172 387104
rect 60608 387064 60614 387076
rect 327166 387064 327172 387076
rect 327224 387104 327230 387116
rect 327902 387104 327908 387116
rect 327224 387076 327908 387104
rect 327224 387064 327230 387076
rect 327902 387064 327908 387076
rect 327960 387064 327966 387116
rect 381538 387064 381544 387116
rect 381596 387104 381602 387116
rect 534350 387104 534356 387116
rect 381596 387076 534356 387104
rect 381596 387064 381602 387076
rect 534350 387064 534356 387076
rect 534408 387064 534414 387116
rect 125594 386384 125600 386436
rect 125652 386424 125658 386436
rect 273990 386424 273996 386436
rect 125652 386396 273996 386424
rect 125652 386384 125658 386396
rect 273990 386384 273996 386396
rect 274048 386384 274054 386436
rect 227714 386316 227720 386368
rect 227772 386356 227778 386368
rect 228358 386356 228364 386368
rect 227772 386328 228364 386356
rect 227772 386316 227778 386328
rect 228358 386316 228364 386328
rect 228416 386356 228422 386368
rect 545390 386356 545396 386368
rect 228416 386328 545396 386356
rect 228416 386316 228422 386328
rect 545390 386316 545396 386328
rect 545448 386316 545454 386368
rect 155954 386248 155960 386300
rect 156012 386288 156018 386300
rect 156414 386288 156420 386300
rect 156012 386260 156420 386288
rect 156012 386248 156018 386260
rect 156414 386248 156420 386260
rect 156472 386288 156478 386300
rect 440234 386288 440240 386300
rect 156472 386260 440240 386288
rect 156472 386248 156478 386260
rect 440234 386248 440240 386260
rect 440292 386248 440298 386300
rect 255314 386180 255320 386232
rect 255372 386220 255378 386232
rect 347866 386220 347872 386232
rect 255372 386192 347872 386220
rect 255372 386180 255378 386192
rect 347866 386180 347872 386192
rect 347924 386180 347930 386232
rect 79318 385636 79324 385688
rect 79376 385676 79382 385688
rect 118602 385676 118608 385688
rect 79376 385648 118608 385676
rect 79376 385636 79382 385648
rect 118602 385636 118608 385648
rect 118660 385636 118666 385688
rect 140682 385636 140688 385688
rect 140740 385676 140746 385688
rect 156414 385676 156420 385688
rect 140740 385648 156420 385676
rect 140740 385636 140746 385648
rect 156414 385636 156420 385648
rect 156472 385636 156478 385688
rect 202138 385636 202144 385688
rect 202196 385676 202202 385688
rect 255314 385676 255320 385688
rect 202196 385648 255320 385676
rect 202196 385636 202202 385648
rect 255314 385636 255320 385648
rect 255372 385636 255378 385688
rect 118602 385024 118608 385076
rect 118660 385064 118666 385076
rect 234706 385064 234712 385076
rect 118660 385036 234712 385064
rect 118660 385024 118666 385036
rect 234706 385024 234712 385036
rect 234764 385024 234770 385076
rect 52362 384956 52368 385008
rect 52420 384996 52426 385008
rect 113174 384996 113180 385008
rect 52420 384968 113180 384996
rect 52420 384956 52426 384968
rect 113174 384956 113180 384968
rect 113232 384996 113238 385008
rect 114462 384996 114468 385008
rect 113232 384968 114468 384996
rect 113232 384956 113238 384968
rect 114462 384956 114468 384968
rect 114520 384956 114526 385008
rect 320818 384956 320824 385008
rect 320876 384996 320882 385008
rect 321462 384996 321468 385008
rect 320876 384968 321468 384996
rect 320876 384956 320882 384968
rect 321462 384956 321468 384968
rect 321520 384996 321526 385008
rect 541158 384996 541164 385008
rect 321520 384968 541164 384996
rect 321520 384956 321526 384968
rect 541158 384956 541164 384968
rect 541216 384956 541222 385008
rect 179874 384412 179880 384464
rect 179932 384452 179938 384464
rect 260098 384452 260104 384464
rect 179932 384424 260104 384452
rect 179932 384412 179938 384424
rect 260098 384412 260104 384424
rect 260156 384412 260162 384464
rect 122742 384344 122748 384396
rect 122800 384384 122806 384396
rect 244274 384384 244280 384396
rect 122800 384356 244280 384384
rect 122800 384344 122806 384356
rect 244274 384344 244280 384356
rect 244332 384344 244338 384396
rect 63494 384276 63500 384328
rect 63552 384316 63558 384328
rect 98638 384316 98644 384328
rect 63552 384288 98644 384316
rect 63552 384276 63558 384288
rect 98638 384276 98644 384288
rect 98696 384276 98702 384328
rect 114462 384276 114468 384328
rect 114520 384316 114526 384328
rect 293310 384316 293316 384328
rect 114520 384288 293316 384316
rect 114520 384276 114526 384288
rect 293310 384276 293316 384288
rect 293368 384276 293374 384328
rect 531958 384276 531964 384328
rect 532016 384316 532022 384328
rect 563054 384316 563060 384328
rect 532016 384288 563060 384316
rect 532016 384276 532022 384288
rect 563054 384276 563060 384288
rect 563112 384276 563118 384328
rect 66254 383460 66260 383512
rect 66312 383500 66318 383512
rect 67266 383500 67272 383512
rect 66312 383472 67272 383500
rect 66312 383460 66318 383472
rect 67266 383460 67272 383472
rect 67324 383460 67330 383512
rect 135898 383052 135904 383104
rect 135956 383092 135962 383104
rect 183554 383092 183560 383104
rect 135956 383064 183560 383092
rect 135956 383052 135962 383064
rect 183554 383052 183560 383064
rect 183612 383092 183618 383104
rect 231118 383092 231124 383104
rect 183612 383064 231124 383092
rect 183612 383052 183618 383064
rect 231118 383052 231124 383064
rect 231176 383052 231182 383104
rect 234614 383052 234620 383104
rect 234672 383092 234678 383104
rect 323118 383092 323124 383104
rect 234672 383064 323124 383092
rect 234672 383052 234678 383064
rect 323118 383052 323124 383064
rect 323176 383092 323182 383104
rect 323176 383064 325694 383092
rect 323176 383052 323182 383064
rect 178678 382984 178684 383036
rect 178736 383024 178742 383036
rect 292574 383024 292580 383036
rect 178736 382996 292580 383024
rect 178736 382984 178742 382996
rect 292574 382984 292580 382996
rect 292632 382984 292638 383036
rect 293310 382984 293316 383036
rect 293368 383024 293374 383036
rect 302970 383024 302976 383036
rect 293368 382996 302976 383024
rect 293368 382984 293374 382996
rect 302970 382984 302976 382996
rect 303028 383024 303034 383036
rect 307018 383024 307024 383036
rect 303028 382996 307024 383024
rect 303028 382984 303034 382996
rect 307018 382984 307024 382996
rect 307076 382984 307082 383036
rect 325666 383024 325694 383064
rect 546678 383024 546684 383036
rect 325666 382996 546684 383024
rect 546678 382984 546684 382996
rect 546736 382984 546742 383036
rect 67266 382916 67272 382968
rect 67324 382956 67330 382968
rect 340966 382956 340972 382968
rect 67324 382928 340972 382956
rect 67324 382916 67330 382928
rect 340966 382916 340972 382928
rect 341024 382916 341030 382968
rect 292574 382168 292580 382220
rect 292632 382208 292638 382220
rect 293126 382208 293132 382220
rect 292632 382180 293132 382208
rect 292632 382168 292638 382180
rect 293126 382168 293132 382180
rect 293184 382208 293190 382220
rect 549346 382208 549352 382220
rect 293184 382180 549352 382208
rect 293184 382168 293190 382180
rect 549346 382168 549352 382180
rect 549404 382168 549410 382220
rect 219434 381624 219440 381676
rect 219492 381664 219498 381676
rect 244918 381664 244924 381676
rect 219492 381636 244924 381664
rect 219492 381624 219498 381636
rect 244918 381624 244924 381636
rect 244976 381624 244982 381676
rect 176562 381556 176568 381608
rect 176620 381596 176626 381608
rect 275278 381596 275284 381608
rect 176620 381568 275284 381596
rect 176620 381556 176626 381568
rect 275278 381556 275284 381568
rect 275336 381556 275342 381608
rect 166902 381488 166908 381540
rect 166960 381528 166966 381540
rect 290458 381528 290464 381540
rect 166960 381500 290464 381528
rect 166960 381488 166966 381500
rect 290458 381488 290464 381500
rect 290516 381488 290522 381540
rect 399478 381488 399484 381540
rect 399536 381528 399542 381540
rect 543826 381528 543832 381540
rect 399536 381500 543832 381528
rect 399536 381488 399542 381500
rect 543826 381488 543832 381500
rect 543884 381488 543890 381540
rect 177942 380196 177948 380248
rect 178000 380236 178006 380248
rect 247770 380236 247776 380248
rect 178000 380208 247776 380236
rect 178000 380196 178006 380208
rect 247770 380196 247776 380208
rect 247828 380196 247834 380248
rect 69106 380128 69112 380180
rect 69164 380168 69170 380180
rect 218698 380168 218704 380180
rect 69164 380140 218704 380168
rect 69164 380128 69170 380140
rect 218698 380128 218704 380140
rect 218756 380128 218762 380180
rect 269758 380128 269764 380180
rect 269816 380168 269822 380180
rect 311894 380168 311900 380180
rect 269816 380140 311900 380168
rect 269816 380128 269822 380140
rect 311894 380128 311900 380140
rect 311952 380128 311958 380180
rect 456794 380128 456800 380180
rect 456852 380168 456858 380180
rect 534258 380168 534264 380180
rect 456852 380140 534264 380168
rect 456852 380128 456858 380140
rect 534258 380128 534264 380140
rect 534316 380128 534322 380180
rect 222194 379584 222200 379636
rect 222252 379624 222258 379636
rect 273898 379624 273904 379636
rect 222252 379596 273904 379624
rect 222252 379584 222258 379596
rect 273898 379584 273904 379596
rect 273956 379584 273962 379636
rect 311894 379584 311900 379636
rect 311952 379624 311958 379636
rect 312722 379624 312728 379636
rect 311952 379596 312728 379624
rect 311952 379584 311958 379596
rect 312722 379584 312728 379596
rect 312780 379624 312786 379636
rect 389174 379624 389180 379636
rect 312780 379596 389180 379624
rect 312780 379584 312786 379596
rect 389174 379584 389180 379596
rect 389232 379624 389238 379636
rect 389818 379624 389824 379636
rect 389232 379596 389824 379624
rect 389232 379584 389238 379596
rect 389818 379584 389824 379596
rect 389876 379584 389882 379636
rect 209774 379516 209780 379568
rect 209832 379556 209838 379568
rect 456794 379556 456800 379568
rect 209832 379528 456800 379556
rect 209832 379516 209838 379528
rect 456794 379516 456800 379528
rect 456852 379516 456858 379568
rect 152918 379448 152924 379500
rect 152976 379488 152982 379500
rect 287698 379488 287704 379500
rect 152976 379460 287704 379488
rect 152976 379448 152982 379460
rect 287698 379448 287704 379460
rect 287756 379448 287762 379500
rect 563054 379448 563060 379500
rect 563112 379488 563118 379500
rect 580166 379488 580172 379500
rect 563112 379460 580172 379488
rect 563112 379448 563118 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 50798 378836 50804 378888
rect 50856 378876 50862 378888
rect 151814 378876 151820 378888
rect 50856 378848 151820 378876
rect 50856 378836 50862 378848
rect 151814 378836 151820 378848
rect 151872 378876 151878 378888
rect 152918 378876 152924 378888
rect 151872 378848 152924 378876
rect 151872 378836 151878 378848
rect 152918 378836 152924 378848
rect 152976 378836 152982 378888
rect 191098 378836 191104 378888
rect 191156 378876 191162 378888
rect 191742 378876 191748 378888
rect 191156 378848 191748 378876
rect 191156 378836 191162 378848
rect 191742 378836 191748 378848
rect 191800 378876 191806 378888
rect 380894 378876 380900 378888
rect 191800 378848 380900 378876
rect 191800 378836 191806 378848
rect 380894 378836 380900 378848
rect 380952 378876 380958 378888
rect 381538 378876 381544 378888
rect 380952 378848 381544 378876
rect 380952 378836 380958 378848
rect 381538 378836 381544 378848
rect 381596 378836 381602 378888
rect 111702 378768 111708 378820
rect 111760 378808 111766 378820
rect 252554 378808 252560 378820
rect 111760 378780 252560 378808
rect 111760 378768 111766 378780
rect 252554 378768 252560 378780
rect 252612 378768 252618 378820
rect 342990 378768 342996 378820
rect 343048 378808 343054 378820
rect 535638 378808 535644 378820
rect 343048 378780 535644 378808
rect 343048 378768 343054 378780
rect 535638 378768 535644 378780
rect 535696 378768 535702 378820
rect 200758 377612 200764 377664
rect 200816 377652 200822 377664
rect 265618 377652 265624 377664
rect 200816 377624 265624 377652
rect 200816 377612 200822 377624
rect 265618 377612 265624 377624
rect 265676 377612 265682 377664
rect 148318 377544 148324 377596
rect 148376 377584 148382 377596
rect 238018 377584 238024 377596
rect 148376 377556 238024 377584
rect 148376 377544 148382 377556
rect 238018 377544 238024 377556
rect 238076 377544 238082 377596
rect 234706 377476 234712 377528
rect 234764 377516 234770 377528
rect 404354 377516 404360 377528
rect 234764 377488 404360 377516
rect 234764 377476 234770 377488
rect 404354 377476 404360 377488
rect 404412 377516 404418 377528
rect 404998 377516 405004 377528
rect 404412 377488 405004 377516
rect 404412 377476 404418 377488
rect 404998 377476 405004 377488
rect 405056 377476 405062 377528
rect 139302 377408 139308 377460
rect 139360 377448 139366 377460
rect 256694 377448 256700 377460
rect 139360 377420 256700 377448
rect 139360 377408 139366 377420
rect 256694 377408 256700 377420
rect 256752 377408 256758 377460
rect 291102 377408 291108 377460
rect 291160 377448 291166 377460
rect 499574 377448 499580 377460
rect 291160 377420 499580 377448
rect 291160 377408 291166 377420
rect 499574 377408 499580 377420
rect 499632 377408 499638 377460
rect 36998 376728 37004 376780
rect 37056 376768 37062 376780
rect 62666 376768 62672 376780
rect 37056 376740 62672 376768
rect 37056 376728 37062 376740
rect 62666 376728 62672 376740
rect 62724 376728 62730 376780
rect 259454 376728 259460 376780
rect 259512 376768 259518 376780
rect 291102 376768 291108 376780
rect 259512 376740 291108 376768
rect 259512 376728 259518 376740
rect 291102 376728 291108 376740
rect 291160 376728 291166 376780
rect 164234 376660 164240 376712
rect 164292 376700 164298 376712
rect 164878 376700 164884 376712
rect 164292 376672 164884 376700
rect 164292 376660 164298 376672
rect 164878 376660 164884 376672
rect 164936 376660 164942 376712
rect 62666 376116 62672 376168
rect 62724 376156 62730 376168
rect 237374 376156 237380 376168
rect 62724 376128 237380 376156
rect 62724 376116 62730 376128
rect 237374 376116 237380 376128
rect 237432 376116 237438 376168
rect 164878 376048 164884 376100
rect 164936 376088 164942 376100
rect 356054 376088 356060 376100
rect 164936 376060 356060 376088
rect 164936 376048 164942 376060
rect 356054 376048 356060 376060
rect 356112 376088 356118 376100
rect 356698 376088 356704 376100
rect 356112 376060 356704 376088
rect 356112 376048 356118 376060
rect 356698 376048 356704 376060
rect 356756 376048 356762 376100
rect 186958 375980 186964 376032
rect 187016 376020 187022 376032
rect 548150 376020 548156 376032
rect 187016 375992 548156 376020
rect 187016 375980 187022 375992
rect 548150 375980 548156 375992
rect 548208 375980 548214 376032
rect 92382 375300 92388 375352
rect 92440 375340 92446 375352
rect 93762 375340 93768 375352
rect 92440 375312 93768 375340
rect 92440 375300 92446 375312
rect 93762 375300 93768 375312
rect 93820 375300 93826 375352
rect 215294 375300 215300 375352
rect 215352 375340 215358 375352
rect 279418 375340 279424 375352
rect 215352 375312 279424 375340
rect 215352 375300 215358 375312
rect 279418 375300 279424 375312
rect 279476 375300 279482 375352
rect 60458 374620 60464 374672
rect 60516 374660 60522 374672
rect 90358 374660 90364 374672
rect 60516 374632 90364 374660
rect 60516 374620 60522 374632
rect 90358 374620 90364 374632
rect 90416 374620 90422 374672
rect 160830 374620 160836 374672
rect 160888 374660 160894 374672
rect 264974 374660 264980 374672
rect 160888 374632 264980 374660
rect 160888 374620 160894 374632
rect 264974 374620 264980 374632
rect 265032 374620 265038 374672
rect 364978 374620 364984 374672
rect 365036 374660 365042 374672
rect 521654 374660 521660 374672
rect 365036 374632 521660 374660
rect 365036 374620 365042 374632
rect 521654 374620 521660 374632
rect 521712 374620 521718 374672
rect 157978 374076 157984 374128
rect 158036 374116 158042 374128
rect 160922 374116 160928 374128
rect 158036 374088 160928 374116
rect 158036 374076 158042 374088
rect 160922 374076 160928 374088
rect 160980 374076 160986 374128
rect 267734 374076 267740 374128
rect 267792 374116 267798 374128
rect 364978 374116 364984 374128
rect 267792 374088 364984 374116
rect 267792 374076 267798 374088
rect 364978 374076 364984 374088
rect 365036 374076 365042 374128
rect 93762 374008 93768 374060
rect 93820 374048 93826 374060
rect 295426 374048 295432 374060
rect 93820 374020 295432 374048
rect 93820 374008 93826 374020
rect 295426 374008 295432 374020
rect 295484 374008 295490 374060
rect 243078 373940 243084 373992
rect 243136 373980 243142 373992
rect 386414 373980 386420 373992
rect 243136 373952 386420 373980
rect 243136 373940 243142 373952
rect 386414 373940 386420 373952
rect 386472 373940 386478 373992
rect 172330 373328 172336 373380
rect 172388 373368 172394 373380
rect 243078 373368 243084 373380
rect 172388 373340 243084 373368
rect 172388 373328 172394 373340
rect 243078 373328 243084 373340
rect 243136 373328 243142 373380
rect 2958 373260 2964 373312
rect 3016 373300 3022 373312
rect 15102 373300 15108 373312
rect 3016 373272 15108 373300
rect 3016 373260 3022 373272
rect 15102 373260 15108 373272
rect 15160 373300 15166 373312
rect 130562 373300 130568 373312
rect 15160 373272 130568 373300
rect 15160 373260 15166 373272
rect 130562 373260 130568 373272
rect 130620 373300 130626 373312
rect 251818 373300 251824 373312
rect 130620 373272 251824 373300
rect 130620 373260 130626 373272
rect 251818 373260 251824 373272
rect 251876 373260 251882 373312
rect 384298 373260 384304 373312
rect 384356 373300 384362 373312
rect 473354 373300 473360 373312
rect 384356 373272 473360 373300
rect 384356 373260 384362 373272
rect 473354 373260 473360 373272
rect 473412 373260 473418 373312
rect 160922 371900 160928 371952
rect 160980 371940 160986 371952
rect 245654 371940 245660 371952
rect 160980 371912 245660 371940
rect 160980 371900 160986 371912
rect 245654 371900 245660 371912
rect 245712 371900 245718 371952
rect 237374 371832 237380 371884
rect 237432 371872 237438 371884
rect 444466 371872 444472 371884
rect 237432 371844 444472 371872
rect 237432 371832 237438 371844
rect 444466 371832 444472 371844
rect 444524 371832 444530 371884
rect 310238 371152 310244 371204
rect 310296 371192 310302 371204
rect 508498 371192 508504 371204
rect 310296 371164 508504 371192
rect 310296 371152 310302 371164
rect 508498 371152 508504 371164
rect 508556 371152 508562 371204
rect 208486 370676 208492 370728
rect 208544 370716 208550 370728
rect 245010 370716 245016 370728
rect 208544 370688 245016 370716
rect 208544 370676 208550 370688
rect 245010 370676 245016 370688
rect 245068 370676 245074 370728
rect 171778 370608 171784 370660
rect 171836 370648 171842 370660
rect 242802 370648 242808 370660
rect 171836 370620 242808 370648
rect 171836 370608 171842 370620
rect 242802 370608 242808 370620
rect 242860 370648 242866 370660
rect 262858 370648 262864 370660
rect 242860 370620 262864 370648
rect 242860 370608 242866 370620
rect 262858 370608 262864 370620
rect 262916 370608 262922 370660
rect 177758 370540 177764 370592
rect 177816 370580 177822 370592
rect 250438 370580 250444 370592
rect 177816 370552 250444 370580
rect 177816 370540 177822 370552
rect 250438 370540 250444 370552
rect 250496 370540 250502 370592
rect 281442 370540 281448 370592
rect 281500 370580 281506 370592
rect 320174 370580 320180 370592
rect 281500 370552 320180 370580
rect 281500 370540 281506 370552
rect 320174 370540 320180 370552
rect 320232 370540 320238 370592
rect 52362 370472 52368 370524
rect 52420 370512 52426 370524
rect 100018 370512 100024 370524
rect 52420 370484 100024 370512
rect 52420 370472 52426 370484
rect 100018 370472 100024 370484
rect 100076 370472 100082 370524
rect 110322 370472 110328 370524
rect 110380 370512 110386 370524
rect 232498 370512 232504 370524
rect 110380 370484 232504 370512
rect 110380 370472 110386 370484
rect 232498 370472 232504 370484
rect 232556 370472 232562 370524
rect 310330 370472 310336 370524
rect 310388 370512 310394 370524
rect 352558 370512 352564 370524
rect 310388 370484 352564 370512
rect 310388 370472 310394 370484
rect 352558 370472 352564 370484
rect 352616 370472 352622 370524
rect 274634 369928 274640 369980
rect 274692 369968 274698 369980
rect 309226 369968 309232 369980
rect 274692 369940 309232 369968
rect 274692 369928 274698 369940
rect 309226 369928 309232 369940
rect 309284 369968 309290 369980
rect 310238 369968 310244 369980
rect 309284 369940 310244 369968
rect 309284 369928 309290 369940
rect 310238 369928 310244 369940
rect 310296 369928 310302 369980
rect 255314 369860 255320 369912
rect 255372 369900 255378 369912
rect 256510 369900 256516 369912
rect 255372 369872 256516 369900
rect 255372 369860 255378 369872
rect 256510 369860 256516 369872
rect 256568 369900 256574 369912
rect 302234 369900 302240 369912
rect 256568 369872 302240 369900
rect 256568 369860 256574 369872
rect 302234 369860 302240 369872
rect 302292 369860 302298 369912
rect 276842 369792 276848 369844
rect 276900 369832 276906 369844
rect 278038 369832 278044 369844
rect 276900 369804 278044 369832
rect 276900 369792 276906 369804
rect 278038 369792 278044 369804
rect 278096 369792 278102 369844
rect 52178 369180 52184 369232
rect 52236 369220 52242 369232
rect 112438 369220 112444 369232
rect 52236 369192 112444 369220
rect 52236 369180 52242 369192
rect 112438 369180 112444 369192
rect 112496 369180 112502 369232
rect 224954 369180 224960 369232
rect 225012 369220 225018 369232
rect 255314 369220 255320 369232
rect 225012 369192 255320 369220
rect 225012 369180 225018 369192
rect 255314 369180 255320 369192
rect 255372 369180 255378 369232
rect 53742 369112 53748 369164
rect 53800 369152 53806 369164
rect 116670 369152 116676 369164
rect 53800 369124 116676 369152
rect 53800 369112 53806 369124
rect 116670 369112 116676 369124
rect 116728 369112 116734 369164
rect 125502 369112 125508 369164
rect 125560 369152 125566 369164
rect 246574 369152 246580 369164
rect 125560 369124 246580 369152
rect 125560 369112 125566 369124
rect 246574 369112 246580 369124
rect 246632 369112 246638 369164
rect 369118 369112 369124 369164
rect 369176 369152 369182 369164
rect 376754 369152 376760 369164
rect 369176 369124 376760 369152
rect 369176 369112 369182 369124
rect 376754 369112 376760 369124
rect 376812 369112 376818 369164
rect 379330 369112 379336 369164
rect 379388 369152 379394 369164
rect 523034 369152 523040 369164
rect 379388 369124 523040 369152
rect 379388 369112 379394 369124
rect 523034 369112 523040 369124
rect 523092 369112 523098 369164
rect 245654 368500 245660 368552
rect 245712 368540 245718 368552
rect 276842 368540 276848 368552
rect 245712 368512 276848 368540
rect 245712 368500 245718 368512
rect 276842 368500 276848 368512
rect 276900 368540 276906 368552
rect 277302 368540 277308 368552
rect 276900 368512 277308 368540
rect 276900 368500 276906 368512
rect 277302 368500 277308 368512
rect 277360 368500 277366 368552
rect 313274 368432 313280 368484
rect 313332 368472 313338 368484
rect 314010 368472 314016 368484
rect 313332 368444 314016 368472
rect 313332 368432 313338 368444
rect 314010 368432 314016 368444
rect 314068 368432 314074 368484
rect 208394 367820 208400 367872
rect 208452 367860 208458 367872
rect 260742 367860 260748 367872
rect 208452 367832 260748 367860
rect 208452 367820 208458 367832
rect 260742 367820 260748 367832
rect 260800 367860 260806 367872
rect 261478 367860 261484 367872
rect 260800 367832 261484 367860
rect 260800 367820 260806 367832
rect 261478 367820 261484 367832
rect 261536 367820 261542 367872
rect 50982 367752 50988 367804
rect 51040 367792 51046 367804
rect 120074 367792 120080 367804
rect 51040 367764 120080 367792
rect 51040 367752 51046 367764
rect 120074 367752 120080 367764
rect 120132 367752 120138 367804
rect 122098 367752 122104 367804
rect 122156 367792 122162 367804
rect 244182 367792 244188 367804
rect 122156 367764 244188 367792
rect 122156 367752 122162 367764
rect 244182 367752 244188 367764
rect 244240 367792 244246 367804
rect 319530 367792 319536 367804
rect 244240 367764 319536 367792
rect 244240 367752 244246 367764
rect 319530 367752 319536 367764
rect 319588 367752 319594 367804
rect 366358 367752 366364 367804
rect 366416 367792 366422 367804
rect 535730 367792 535736 367804
rect 366416 367764 535736 367792
rect 366416 367752 366422 367764
rect 535730 367752 535736 367764
rect 535788 367752 535794 367804
rect 263594 367276 263600 367328
rect 263652 367316 263658 367328
rect 264882 367316 264888 367328
rect 263652 367288 264888 367316
rect 263652 367276 263658 367288
rect 264882 367276 264888 367288
rect 264940 367316 264946 367328
rect 309962 367316 309968 367328
rect 264940 367288 309968 367316
rect 264940 367276 264946 367288
rect 309962 367276 309968 367288
rect 310020 367276 310026 367328
rect 218054 367208 218060 367260
rect 218112 367248 218118 367260
rect 313274 367248 313280 367260
rect 218112 367220 313280 367248
rect 218112 367208 218118 367220
rect 313274 367208 313280 367220
rect 313332 367208 313338 367260
rect 145558 367140 145564 367192
rect 145616 367180 145622 367192
rect 208486 367180 208492 367192
rect 145616 367152 208492 367180
rect 145616 367140 145622 367152
rect 208486 367140 208492 367152
rect 208544 367140 208550 367192
rect 255958 367140 255964 367192
rect 256016 367180 256022 367192
rect 256602 367180 256608 367192
rect 256016 367152 256608 367180
rect 256016 367140 256022 367152
rect 256602 367140 256608 367152
rect 256660 367180 256666 367192
rect 403618 367180 403624 367192
rect 256660 367152 403624 367180
rect 256660 367140 256666 367152
rect 403618 367140 403624 367152
rect 403676 367140 403682 367192
rect 300854 367112 300860 367124
rect 128372 367084 300860 367112
rect 128372 367056 128400 367084
rect 300854 367072 300860 367084
rect 300912 367072 300918 367124
rect 66898 367004 66904 367056
rect 66956 367044 66962 367056
rect 128354 367044 128360 367056
rect 66956 367016 128360 367044
rect 66956 367004 66962 367016
rect 128354 367004 128360 367016
rect 128412 367004 128418 367056
rect 301038 367004 301044 367056
rect 301096 367044 301102 367056
rect 301498 367044 301504 367056
rect 301096 367016 301504 367044
rect 301096 367004 301102 367016
rect 301498 367004 301504 367016
rect 301556 367004 301562 367056
rect 53466 366324 53472 366376
rect 53524 366364 53530 366376
rect 138014 366364 138020 366376
rect 53524 366336 138020 366364
rect 53524 366324 53530 366336
rect 138014 366324 138020 366336
rect 138072 366324 138078 366376
rect 216674 366324 216680 366376
rect 216732 366364 216738 366376
rect 263594 366364 263600 366376
rect 216732 366336 263600 366364
rect 216732 366324 216738 366336
rect 263594 366324 263600 366336
rect 263652 366324 263658 366376
rect 417418 366324 417424 366376
rect 417476 366364 417482 366376
rect 477494 366364 477500 366376
rect 417476 366336 477500 366364
rect 417476 366324 417482 366336
rect 477494 366324 477500 366336
rect 477552 366324 477558 366376
rect 283650 365916 283656 365968
rect 283708 365956 283714 365968
rect 423674 365956 423680 365968
rect 283708 365928 423680 365956
rect 283708 365916 283714 365928
rect 423674 365916 423680 365928
rect 423732 365956 423738 365968
rect 424318 365956 424324 365968
rect 423732 365928 424324 365956
rect 423732 365916 423738 365928
rect 424318 365916 424324 365928
rect 424376 365916 424382 365968
rect 189074 365848 189080 365900
rect 189132 365888 189138 365900
rect 338758 365888 338764 365900
rect 189132 365860 338764 365888
rect 189132 365848 189138 365860
rect 338758 365848 338764 365860
rect 338816 365848 338822 365900
rect 138014 365780 138020 365832
rect 138072 365820 138078 365832
rect 296806 365820 296812 365832
rect 138072 365792 296812 365820
rect 138072 365780 138078 365792
rect 296806 365780 296812 365792
rect 296864 365780 296870 365832
rect 101398 365712 101404 365764
rect 101456 365752 101462 365764
rect 301038 365752 301044 365764
rect 101456 365724 301044 365752
rect 101456 365712 101462 365724
rect 301038 365712 301044 365724
rect 301096 365712 301102 365764
rect 273990 365644 273996 365696
rect 274048 365684 274054 365696
rect 274542 365684 274548 365696
rect 274048 365656 274548 365684
rect 274048 365644 274054 365656
rect 274542 365644 274548 365656
rect 274600 365684 274606 365696
rect 300302 365684 300308 365696
rect 274600 365656 300308 365684
rect 274600 365644 274606 365656
rect 300302 365644 300308 365656
rect 300360 365644 300366 365696
rect 544378 365644 544384 365696
rect 544436 365684 544442 365696
rect 580166 365684 580172 365696
rect 544436 365656 580172 365684
rect 544436 365644 544442 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 314010 365208 314016 365220
rect 267706 365180 314016 365208
rect 179230 365100 179236 365152
rect 179288 365140 179294 365152
rect 264238 365140 264244 365152
rect 179288 365112 264244 365140
rect 179288 365100 179294 365112
rect 264238 365100 264244 365112
rect 264296 365140 264302 365152
rect 267706 365140 267734 365180
rect 314010 365168 314016 365180
rect 314068 365168 314074 365220
rect 264296 365112 267734 365140
rect 264296 365100 264302 365112
rect 300762 365100 300768 365152
rect 300820 365140 300826 365152
rect 372614 365140 372620 365152
rect 300820 365112 372620 365140
rect 300820 365100 300826 365112
rect 372614 365100 372620 365112
rect 372672 365100 372678 365152
rect 173710 365032 173716 365084
rect 173768 365072 173774 365084
rect 173768 365044 277394 365072
rect 173768 365032 173774 365044
rect 42610 364964 42616 365016
rect 42668 365004 42674 365016
rect 96614 365004 96620 365016
rect 42668 364976 96620 365004
rect 42668 364964 42674 364976
rect 96614 364964 96620 364976
rect 96672 364964 96678 365016
rect 126238 364964 126244 365016
rect 126296 365004 126302 365016
rect 245746 365004 245752 365016
rect 126296 364976 245752 365004
rect 126296 364964 126302 364976
rect 245746 364964 245752 364976
rect 245804 364964 245810 365016
rect 277366 365004 277394 365044
rect 363598 365032 363604 365084
rect 363656 365072 363662 365084
rect 440326 365072 440332 365084
rect 363656 365044 440332 365072
rect 363656 365032 363662 365044
rect 440326 365032 440332 365044
rect 440384 365032 440390 365084
rect 279510 365004 279516 365016
rect 277366 364976 279516 365004
rect 279510 364964 279516 364976
rect 279568 365004 279574 365016
rect 418798 365004 418804 365016
rect 279568 364976 418804 365004
rect 279568 364964 279574 364976
rect 418798 364964 418804 364976
rect 418856 364964 418862 365016
rect 96614 364420 96620 364472
rect 96672 364460 96678 364472
rect 300946 364460 300952 364472
rect 96672 364432 300952 364460
rect 96672 364420 96678 364432
rect 300946 364420 300952 364432
rect 301004 364420 301010 364472
rect 83458 364352 83464 364404
rect 83516 364392 83522 364404
rect 307846 364392 307852 364404
rect 83516 364364 307852 364392
rect 83516 364352 83522 364364
rect 307846 364352 307852 364364
rect 307904 364352 307910 364404
rect 273898 363808 273904 363860
rect 273956 363848 273962 363860
rect 298186 363848 298192 363860
rect 273956 363820 298192 363848
rect 273956 363808 273962 363820
rect 298186 363808 298192 363820
rect 298244 363808 298250 363860
rect 277302 363740 277308 363792
rect 277360 363780 277366 363792
rect 347038 363780 347044 363792
rect 277360 363752 347044 363780
rect 277360 363740 277366 363752
rect 347038 363740 347044 363752
rect 347096 363740 347102 363792
rect 228818 363672 228824 363724
rect 228876 363712 228882 363724
rect 336642 363712 336648 363724
rect 228876 363684 336648 363712
rect 228876 363672 228882 363684
rect 336642 363672 336648 363684
rect 336700 363672 336706 363724
rect 41230 363604 41236 363656
rect 41288 363644 41294 363656
rect 304994 363644 305000 363656
rect 41288 363616 305000 363644
rect 41288 363604 41294 363616
rect 304994 363604 305000 363616
rect 305052 363604 305058 363656
rect 389818 363604 389824 363656
rect 389876 363644 389882 363656
rect 431954 363644 431960 363656
rect 389876 363616 431960 363644
rect 389876 363604 389882 363616
rect 431954 363604 431960 363616
rect 432012 363604 432018 363656
rect 432046 363604 432052 363656
rect 432104 363644 432110 363656
rect 452654 363644 452660 363656
rect 432104 363616 452660 363644
rect 432104 363604 432110 363616
rect 452654 363604 452660 363616
rect 452712 363604 452718 363656
rect 304994 363400 305000 363452
rect 305052 363440 305058 363452
rect 305730 363440 305736 363452
rect 305052 363412 305736 363440
rect 305052 363400 305058 363412
rect 305730 363400 305736 363412
rect 305788 363400 305794 363452
rect 144178 362992 144184 363044
rect 144236 363032 144242 363044
rect 212534 363032 212540 363044
rect 144236 363004 212540 363032
rect 144236 362992 144242 363004
rect 212534 362992 212540 363004
rect 212592 362992 212598 363044
rect 245746 362992 245752 363044
rect 245804 363032 245810 363044
rect 246942 363032 246948 363044
rect 245804 363004 246948 363032
rect 245804 362992 245810 363004
rect 246942 362992 246948 363004
rect 247000 363032 247006 363044
rect 315390 363032 315396 363044
rect 247000 363004 315396 363032
rect 247000 362992 247006 363004
rect 315390 362992 315396 363004
rect 315448 362992 315454 363044
rect 162302 362924 162308 362976
rect 162360 362964 162366 362976
rect 162762 362964 162768 362976
rect 162360 362936 162768 362964
rect 162360 362924 162366 362936
rect 162762 362924 162768 362936
rect 162820 362964 162826 362976
rect 294046 362964 294052 362976
rect 162820 362936 294052 362964
rect 162820 362924 162826 362936
rect 294046 362924 294052 362936
rect 294104 362924 294110 362976
rect 336642 362924 336648 362976
rect 336700 362964 336706 362976
rect 340874 362964 340880 362976
rect 336700 362936 340880 362964
rect 336700 362924 336706 362936
rect 340874 362924 340880 362936
rect 340932 362924 340938 362976
rect 212534 362312 212540 362364
rect 212592 362352 212598 362364
rect 256694 362352 256700 362364
rect 212592 362324 256700 362352
rect 212592 362312 212598 362324
rect 256694 362312 256700 362324
rect 256752 362312 256758 362364
rect 140038 362244 140044 362296
rect 140096 362284 140102 362296
rect 245746 362284 245752 362296
rect 140096 362256 245752 362284
rect 140096 362244 140102 362256
rect 245746 362244 245752 362256
rect 245804 362244 245810 362296
rect 95142 362176 95148 362228
rect 95200 362216 95206 362228
rect 117958 362216 117964 362228
rect 95200 362188 117964 362216
rect 95200 362176 95206 362188
rect 117958 362176 117964 362188
rect 118016 362176 118022 362228
rect 122650 362176 122656 362228
rect 122708 362216 122714 362228
rect 242986 362216 242992 362228
rect 122708 362188 242992 362216
rect 122708 362176 122714 362188
rect 242986 362176 242992 362188
rect 243044 362176 243050 362228
rect 258902 362176 258908 362228
rect 258960 362216 258966 362228
rect 289722 362216 289728 362228
rect 258960 362188 289728 362216
rect 258960 362176 258966 362188
rect 289722 362176 289728 362188
rect 289780 362216 289786 362228
rect 336734 362216 336740 362228
rect 289780 362188 336740 362216
rect 289780 362176 289786 362188
rect 336734 362176 336740 362188
rect 336792 362176 336798 362228
rect 340138 361700 340144 361752
rect 340196 361740 340202 361752
rect 413278 361740 413284 361752
rect 340196 361712 413284 361740
rect 340196 361700 340202 361712
rect 413278 361700 413284 361712
rect 413336 361700 413342 361752
rect 153102 361632 153108 361684
rect 153160 361672 153166 361684
rect 201586 361672 201592 361684
rect 153160 361644 201592 361672
rect 153160 361632 153166 361644
rect 201586 361632 201592 361644
rect 201644 361672 201650 361684
rect 202138 361672 202144 361684
rect 201644 361644 202144 361672
rect 201644 361632 201650 361644
rect 202138 361632 202144 361644
rect 202196 361632 202202 361684
rect 227346 361632 227352 361684
rect 227404 361672 227410 361684
rect 227622 361672 227628 361684
rect 227404 361644 227628 361672
rect 227404 361632 227410 361644
rect 227622 361632 227628 361644
rect 227680 361672 227686 361684
rect 342254 361672 342260 361684
rect 227680 361644 342260 361672
rect 227680 361632 227686 361644
rect 342254 361632 342260 361644
rect 342312 361632 342318 361684
rect 175090 361564 175096 361616
rect 175148 361604 175154 361616
rect 359458 361604 359464 361616
rect 175148 361576 359464 361604
rect 175148 361564 175154 361576
rect 359458 361564 359464 361576
rect 359516 361564 359522 361616
rect 287698 360816 287704 360868
rect 287756 360856 287762 360868
rect 316126 360856 316132 360868
rect 287756 360828 316132 360856
rect 287756 360816 287762 360828
rect 316126 360816 316132 360828
rect 316184 360816 316190 360868
rect 250530 360340 250536 360392
rect 250588 360380 250594 360392
rect 251082 360380 251088 360392
rect 250588 360352 251088 360380
rect 250588 360340 250594 360352
rect 251082 360340 251088 360352
rect 251140 360380 251146 360392
rect 349430 360380 349436 360392
rect 251140 360352 349436 360380
rect 251140 360340 251146 360352
rect 349430 360340 349436 360352
rect 349488 360340 349494 360392
rect 113174 360272 113180 360324
rect 113232 360312 113238 360324
rect 317506 360312 317512 360324
rect 113232 360284 317512 360312
rect 113232 360272 113238 360284
rect 317506 360272 317512 360284
rect 317564 360272 317570 360324
rect 70394 360204 70400 360256
rect 70452 360244 70458 360256
rect 71130 360244 71136 360256
rect 70452 360216 71136 360244
rect 70452 360204 70458 360216
rect 71130 360204 71136 360216
rect 71188 360244 71194 360256
rect 291194 360244 291200 360256
rect 71188 360216 291200 360244
rect 71188 360204 71194 360216
rect 291194 360204 291200 360216
rect 291252 360204 291258 360256
rect 243906 359660 243912 359712
rect 243964 359700 243970 359712
rect 277394 359700 277400 359712
rect 243964 359672 277400 359700
rect 243964 359660 243970 359672
rect 277366 359660 277400 359672
rect 277452 359660 277458 359712
rect 177850 359592 177856 359644
rect 177908 359632 177914 359644
rect 254578 359632 254584 359644
rect 177908 359604 254584 359632
rect 177908 359592 177914 359604
rect 254578 359592 254584 359604
rect 254636 359592 254642 359644
rect 166626 359524 166632 359576
rect 166684 359564 166690 359576
rect 248414 359564 248420 359576
rect 166684 359536 248420 359564
rect 166684 359524 166690 359536
rect 248414 359524 248420 359536
rect 248472 359524 248478 359576
rect 170950 359456 170956 359508
rect 171008 359496 171014 359508
rect 255958 359496 255964 359508
rect 171008 359468 255964 359496
rect 171008 359456 171014 359468
rect 255958 359456 255964 359468
rect 256016 359456 256022 359508
rect 277366 359496 277394 359660
rect 375098 359496 375104 359508
rect 277366 359468 375104 359496
rect 375098 359456 375104 359468
rect 375156 359496 375162 359508
rect 391934 359496 391940 359508
rect 375156 359468 391940 359496
rect 375156 359456 375162 359468
rect 391934 359456 391940 359468
rect 391992 359456 391998 359508
rect 393958 359456 393964 359508
rect 394016 359496 394022 359508
rect 489914 359496 489920 359508
rect 394016 359468 489920 359496
rect 394016 359456 394022 359468
rect 489914 359456 489920 359468
rect 489972 359456 489978 359508
rect 68278 358912 68284 358964
rect 68336 358952 68342 358964
rect 193398 358952 193404 358964
rect 68336 358924 193404 358952
rect 68336 358912 68342 358924
rect 193398 358912 193404 358924
rect 193456 358912 193462 358964
rect 349798 358952 349804 358964
rect 277366 358924 349804 358952
rect 146938 358844 146944 358896
rect 146996 358884 147002 358896
rect 276658 358884 276664 358896
rect 146996 358856 276664 358884
rect 146996 358844 147002 358856
rect 276658 358844 276664 358856
rect 276716 358884 276722 358896
rect 277118 358884 277124 358896
rect 276716 358856 277124 358884
rect 276716 358844 276722 358856
rect 277118 358844 277124 358856
rect 277176 358884 277182 358896
rect 277366 358884 277394 358924
rect 349798 358912 349804 358924
rect 349856 358912 349862 358964
rect 277176 358856 277394 358884
rect 277176 358844 277182 358856
rect 279418 358844 279424 358896
rect 279476 358884 279482 358896
rect 454034 358884 454040 358896
rect 279476 358856 454040 358884
rect 279476 358844 279482 358856
rect 454034 358844 454040 358856
rect 454092 358844 454098 358896
rect 166258 358776 166264 358828
rect 166316 358816 166322 358828
rect 166810 358816 166816 358828
rect 166316 358788 166816 358816
rect 166316 358776 166322 358788
rect 166810 358776 166816 358788
rect 166868 358816 166874 358828
rect 445018 358816 445024 358828
rect 166868 358788 445024 358816
rect 166868 358776 166874 358788
rect 445018 358776 445024 358788
rect 445076 358776 445082 358828
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 4798 358476 4804 358488
rect 2832 358448 4804 358476
rect 2832 358436 2838 358448
rect 4798 358436 4804 358448
rect 4856 358436 4862 358488
rect 290458 358096 290464 358148
rect 290516 358136 290522 358148
rect 298002 358136 298008 358148
rect 290516 358108 298008 358136
rect 290516 358096 290522 358108
rect 298002 358096 298008 358108
rect 298060 358096 298066 358148
rect 175918 357756 175924 357808
rect 175976 357796 175982 357808
rect 195238 357796 195244 357808
rect 175976 357768 195244 357796
rect 175976 357756 175982 357768
rect 195238 357756 195244 357768
rect 195296 357756 195302 357808
rect 212350 357756 212356 357808
rect 212408 357796 212414 357808
rect 214558 357796 214564 357808
rect 212408 357768 214564 357796
rect 212408 357756 212414 357768
rect 214558 357756 214564 357768
rect 214616 357756 214622 357808
rect 285950 357756 285956 357808
rect 286008 357796 286014 357808
rect 286962 357796 286968 357808
rect 286008 357768 286968 357796
rect 286008 357756 286014 357768
rect 286962 357756 286968 357768
rect 287020 357796 287026 357808
rect 306374 357796 306380 357808
rect 287020 357768 306380 357796
rect 287020 357756 287026 357768
rect 306374 357756 306380 357768
rect 306432 357756 306438 357808
rect 162118 357688 162124 357740
rect 162176 357728 162182 357740
rect 247678 357728 247684 357740
rect 162176 357700 247684 357728
rect 162176 357688 162182 357700
rect 247678 357688 247684 357700
rect 247736 357728 247742 357740
rect 248138 357728 248144 357740
rect 247736 357700 248144 357728
rect 247736 357688 247742 357700
rect 248138 357688 248144 357700
rect 248196 357728 248202 357740
rect 262858 357728 262864 357740
rect 248196 357700 262864 357728
rect 248196 357688 248202 357700
rect 262858 357688 262864 357700
rect 262916 357688 262922 357740
rect 265342 357688 265348 357740
rect 265400 357728 265406 357740
rect 265618 357728 265624 357740
rect 265400 357700 265624 357728
rect 265400 357688 265406 357700
rect 265618 357688 265624 357700
rect 265676 357728 265682 357740
rect 300302 357728 300308 357740
rect 265676 357700 300308 357728
rect 265676 357688 265682 357700
rect 300302 357688 300308 357700
rect 300360 357688 300366 357740
rect 170490 357620 170496 357672
rect 170548 357660 170554 357672
rect 283650 357660 283656 357672
rect 170548 357632 283656 357660
rect 170548 357620 170554 357632
rect 283650 357620 283656 357632
rect 283708 357660 283714 357672
rect 287330 357660 287336 357672
rect 283708 357632 287336 357660
rect 283708 357620 283714 357632
rect 287330 357620 287336 357632
rect 287388 357620 287394 357672
rect 91738 357552 91744 357604
rect 91796 357592 91802 357604
rect 212442 357592 212448 357604
rect 91796 357564 212448 357592
rect 91796 357552 91802 357564
rect 212442 357552 212448 357564
rect 212500 357552 212506 357604
rect 231118 357552 231124 357604
rect 231176 357592 231182 357604
rect 293218 357592 293224 357604
rect 231176 357564 293224 357592
rect 231176 357552 231182 357564
rect 293218 357552 293224 357564
rect 293276 357552 293282 357604
rect 169110 357484 169116 357536
rect 169168 357524 169174 357536
rect 202874 357524 202880 357536
rect 169168 357496 202880 357524
rect 169168 357484 169174 357496
rect 202874 357484 202880 357496
rect 202932 357524 202938 357536
rect 307754 357524 307760 357536
rect 202932 357496 307760 357524
rect 202932 357484 202938 357496
rect 307754 357484 307760 357496
rect 307812 357484 307818 357536
rect 43990 357416 43996 357468
rect 44048 357456 44054 357468
rect 243906 357456 243912 357468
rect 44048 357428 243912 357456
rect 44048 357416 44054 357428
rect 243906 357416 243912 357428
rect 243964 357416 243970 357468
rect 251082 357416 251088 357468
rect 251140 357456 251146 357468
rect 253934 357456 253940 357468
rect 251140 357428 253940 357456
rect 251140 357416 251146 357428
rect 253934 357416 253940 357428
rect 253992 357416 253998 357468
rect 256694 357416 256700 357468
rect 256752 357456 256758 357468
rect 304534 357456 304540 357468
rect 256752 357428 304540 357456
rect 256752 357416 256758 357428
rect 304534 357416 304540 357428
rect 304592 357416 304598 357468
rect 212442 357348 212448 357400
rect 212500 357388 212506 357400
rect 261570 357388 261576 357400
rect 212500 357360 261576 357388
rect 212500 357348 212506 357360
rect 261570 357348 261576 357360
rect 261628 357388 261634 357400
rect 262122 357388 262128 357400
rect 261628 357360 262128 357388
rect 261628 357348 261634 357360
rect 262122 357348 262128 357360
rect 262180 357348 262186 357400
rect 273714 357348 273720 357400
rect 273772 357388 273778 357400
rect 274542 357388 274548 357400
rect 273772 357360 274548 357388
rect 273772 357348 273778 357360
rect 274542 357348 274548 357360
rect 274600 357348 274606 357400
rect 117958 356736 117964 356788
rect 118016 356776 118022 356788
rect 212350 356776 212356 356788
rect 118016 356748 212356 356776
rect 118016 356736 118022 356748
rect 212350 356736 212356 356748
rect 212408 356736 212414 356788
rect 262122 356736 262128 356788
rect 262180 356776 262186 356788
rect 297450 356776 297456 356788
rect 262180 356748 297456 356776
rect 262180 356736 262186 356748
rect 297450 356736 297456 356748
rect 297508 356736 297514 356788
rect 109678 356668 109684 356720
rect 109736 356708 109742 356720
rect 251082 356708 251088 356720
rect 109736 356680 251088 356708
rect 109736 356668 109742 356680
rect 251082 356668 251088 356680
rect 251140 356668 251146 356720
rect 262858 356668 262864 356720
rect 262916 356708 262922 356720
rect 429838 356708 429844 356720
rect 262916 356680 429844 356708
rect 262916 356668 262922 356680
rect 429838 356668 429844 356680
rect 429896 356668 429902 356720
rect 171134 356260 171140 356312
rect 171192 356300 171198 356312
rect 199654 356300 199660 356312
rect 171192 356272 199660 356300
rect 171192 356260 171198 356272
rect 199654 356260 199660 356272
rect 199712 356260 199718 356312
rect 262766 356260 262772 356312
rect 262824 356300 262830 356312
rect 351178 356300 351184 356312
rect 262824 356272 351184 356300
rect 262824 356260 262830 356272
rect 351178 356260 351184 356272
rect 351236 356260 351242 356312
rect 154482 356192 154488 356244
rect 154540 356232 154546 356244
rect 186774 356232 186780 356244
rect 154540 356204 186780 356232
rect 154540 356192 154546 356204
rect 186774 356192 186780 356204
rect 186832 356192 186838 356244
rect 193398 356192 193404 356244
rect 193456 356232 193462 356244
rect 297634 356232 297640 356244
rect 193456 356204 297640 356232
rect 193456 356192 193462 356204
rect 297634 356192 297640 356204
rect 297692 356192 297698 356244
rect 134610 356124 134616 356176
rect 134668 356164 134674 356176
rect 266354 356164 266360 356176
rect 134668 356136 266360 356164
rect 134668 356124 134674 356136
rect 266354 356124 266360 356136
rect 266412 356164 266418 356176
rect 266814 356164 266820 356176
rect 266412 356136 266820 356164
rect 266412 356124 266418 356136
rect 266814 356124 266820 356136
rect 266872 356164 266878 356176
rect 270402 356164 270408 356176
rect 266872 356136 270408 356164
rect 266872 356124 266878 356136
rect 270402 356124 270408 356136
rect 270460 356124 270466 356176
rect 273714 356124 273720 356176
rect 273772 356164 273778 356176
rect 298738 356164 298744 356176
rect 273772 356136 298744 356164
rect 273772 356124 273778 356136
rect 298738 356124 298744 356136
rect 298796 356124 298802 356176
rect 170582 356056 170588 356108
rect 170640 356096 170646 356108
rect 326430 356096 326436 356108
rect 170640 356068 326436 356096
rect 170640 356056 170646 356068
rect 326430 356056 326436 356068
rect 326488 356056 326494 356108
rect 270402 355988 270408 356040
rect 270460 356028 270466 356040
rect 417418 356028 417424 356040
rect 270460 356000 417424 356028
rect 270460 355988 270466 356000
rect 417418 355988 417424 356000
rect 417476 355988 417482 356040
rect 164142 355444 164148 355496
rect 164200 355484 164206 355496
rect 191098 355484 191104 355496
rect 164200 355456 191104 355484
rect 164200 355444 164206 355456
rect 191098 355444 191104 355456
rect 191156 355444 191162 355496
rect 49418 355376 49424 355428
rect 49476 355416 49482 355428
rect 166994 355416 167000 355428
rect 49476 355388 167000 355416
rect 49476 355376 49482 355388
rect 166994 355376 167000 355388
rect 167052 355376 167058 355428
rect 173802 355376 173808 355428
rect 173860 355416 173866 355428
rect 189718 355416 189724 355428
rect 173860 355388 189724 355416
rect 173860 355376 173866 355388
rect 189718 355376 189724 355388
rect 189776 355376 189782 355428
rect 254394 355376 254400 355428
rect 254452 355416 254458 355428
rect 425698 355416 425704 355428
rect 254452 355388 425704 355416
rect 254452 355376 254458 355388
rect 425698 355376 425704 355388
rect 425756 355376 425762 355428
rect 112530 355308 112536 355360
rect 112588 355348 112594 355360
rect 289170 355348 289176 355360
rect 112588 355320 289176 355348
rect 112588 355308 112594 355320
rect 289170 355308 289176 355320
rect 289228 355348 289234 355360
rect 295518 355348 295524 355360
rect 289228 355320 295524 355348
rect 289228 355308 289234 355320
rect 295518 355308 295524 355320
rect 295576 355308 295582 355360
rect 424318 355308 424324 355360
rect 424376 355348 424382 355360
rect 450538 355348 450544 355360
rect 424376 355320 450544 355348
rect 424376 355308 424382 355320
rect 450538 355308 450544 355320
rect 450596 355308 450602 355360
rect 292298 354900 292304 354952
rect 292356 354940 292362 354952
rect 292574 354940 292580 354952
rect 292356 354912 292580 354940
rect 292356 354900 292362 354912
rect 292574 354900 292580 354912
rect 292632 354900 292638 354952
rect 179414 354832 179420 354884
rect 179472 354872 179478 354884
rect 219434 354872 219440 354884
rect 179472 354844 219440 354872
rect 179472 354832 179478 354844
rect 219434 354832 219440 354844
rect 219492 354872 219498 354884
rect 220446 354872 220452 354884
rect 219492 354844 220452 354872
rect 219492 354832 219498 354844
rect 220446 354832 220452 354844
rect 220504 354872 220510 354884
rect 301498 354872 301504 354884
rect 220504 354844 301504 354872
rect 220504 354832 220510 354844
rect 301498 354832 301504 354844
rect 301556 354832 301562 354884
rect 174538 354764 174544 354816
rect 174596 354804 174602 354816
rect 279050 354804 279056 354816
rect 174596 354776 279056 354804
rect 174596 354764 174602 354776
rect 279050 354764 279056 354776
rect 279108 354764 279114 354816
rect 284018 354764 284024 354816
rect 284076 354804 284082 354816
rect 302878 354804 302884 354816
rect 284076 354776 302884 354804
rect 284076 354764 284082 354776
rect 302878 354764 302884 354776
rect 302936 354764 302942 354816
rect 166994 354696 167000 354748
rect 167052 354736 167058 354748
rect 209866 354736 209872 354748
rect 167052 354708 209872 354736
rect 167052 354696 167058 354708
rect 209866 354696 209872 354708
rect 209924 354696 209930 354748
rect 271138 354696 271144 354748
rect 271196 354736 271202 354748
rect 385034 354736 385040 354748
rect 271196 354708 385040 354736
rect 271196 354696 271202 354708
rect 385034 354696 385040 354708
rect 385092 354696 385098 354748
rect 292482 354492 292488 354544
rect 292540 354532 292546 354544
rect 293310 354532 293316 354544
rect 292540 354504 293316 354532
rect 292540 354492 292546 354504
rect 293310 354492 293316 354504
rect 293368 354492 293374 354544
rect 295426 354424 295432 354476
rect 295484 354464 295490 354476
rect 295610 354464 295616 354476
rect 295484 354436 295616 354464
rect 295484 354424 295490 354436
rect 295610 354424 295616 354436
rect 295668 354424 295674 354476
rect 53742 353948 53748 354000
rect 53800 353988 53806 354000
rect 179414 353988 179420 354000
rect 53800 353960 179420 353988
rect 53800 353948 53806 353960
rect 179414 353948 179420 353960
rect 179472 353948 179478 354000
rect 295426 353268 295432 353320
rect 295484 353308 295490 353320
rect 346302 353308 346308 353320
rect 295484 353280 346308 353308
rect 295484 353268 295490 353280
rect 346302 353268 346308 353280
rect 346360 353268 346366 353320
rect 43898 353200 43904 353252
rect 43956 353240 43962 353252
rect 171134 353240 171140 353252
rect 43956 353212 171140 353240
rect 43956 353200 43962 353212
rect 171134 353200 171140 353212
rect 171192 353200 171198 353252
rect 54938 352520 54944 352572
rect 54996 352560 55002 352572
rect 68278 352560 68284 352572
rect 54996 352532 68284 352560
rect 54996 352520 55002 352532
rect 68278 352520 68284 352532
rect 68336 352520 68342 352572
rect 295426 352520 295432 352572
rect 295484 352560 295490 352572
rect 297910 352560 297916 352572
rect 295484 352532 297916 352560
rect 295484 352520 295490 352532
rect 297910 352520 297916 352532
rect 297968 352560 297974 352572
rect 297968 352532 335354 352560
rect 297968 352520 297974 352532
rect 335326 352492 335354 352532
rect 346302 352520 346308 352572
rect 346360 352560 346366 352572
rect 442166 352560 442172 352572
rect 346360 352532 442172 352560
rect 346360 352520 346366 352532
rect 442166 352520 442172 352532
rect 442224 352520 442230 352572
rect 345658 352492 345664 352504
rect 335326 352464 345664 352492
rect 345658 352452 345664 352464
rect 345716 352452 345722 352504
rect 437382 351908 437388 351960
rect 437440 351948 437446 351960
rect 580166 351948 580172 351960
rect 437440 351920 580172 351948
rect 437440 351908 437446 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 442166 351840 442172 351892
rect 442224 351880 442230 351892
rect 442902 351880 442908 351892
rect 442224 351852 442908 351880
rect 442224 351840 442230 351852
rect 442902 351840 442908 351852
rect 442960 351880 442966 351892
rect 548058 351880 548064 351892
rect 442960 351852 548064 351880
rect 442960 351840 442966 351852
rect 548058 351840 548064 351852
rect 548116 351840 548122 351892
rect 293218 351160 293224 351212
rect 293276 351200 293282 351212
rect 438854 351200 438860 351212
rect 293276 351172 438860 351200
rect 293276 351160 293282 351172
rect 438854 351160 438860 351172
rect 438912 351160 438918 351212
rect 295426 350480 295432 350532
rect 295484 350520 295490 350532
rect 302326 350520 302332 350532
rect 295484 350492 302332 350520
rect 295484 350480 295490 350492
rect 302326 350480 302332 350492
rect 302384 350520 302390 350532
rect 302970 350520 302976 350532
rect 302384 350492 302976 350520
rect 302384 350480 302390 350492
rect 302970 350480 302976 350492
rect 303028 350480 303034 350532
rect 438854 350480 438860 350532
rect 438912 350520 438918 350532
rect 440142 350520 440148 350532
rect 438912 350492 440148 350520
rect 438912 350480 438918 350492
rect 440142 350480 440148 350492
rect 440200 350520 440206 350532
rect 547874 350520 547880 350532
rect 440200 350492 547880 350520
rect 440200 350480 440206 350492
rect 547874 350480 547880 350492
rect 547932 350480 547938 350532
rect 45278 349800 45284 349852
rect 45336 349840 45342 349852
rect 171778 349840 171784 349852
rect 45336 349812 171784 349840
rect 45336 349800 45342 349812
rect 171778 349800 171784 349812
rect 171836 349800 171842 349852
rect 302326 349800 302332 349852
rect 302384 349840 302390 349852
rect 325142 349840 325148 349852
rect 302384 349812 325148 349840
rect 302384 349800 302390 349812
rect 325142 349800 325148 349812
rect 325200 349800 325206 349852
rect 63218 348372 63224 348424
rect 63276 348412 63282 348424
rect 133138 348412 133144 348424
rect 63276 348384 133144 348412
rect 63276 348372 63282 348384
rect 133138 348372 133144 348384
rect 133196 348372 133202 348424
rect 429102 348372 429108 348424
rect 429160 348412 429166 348424
rect 574738 348412 574744 348424
rect 429160 348384 574744 348412
rect 429160 348372 429166 348384
rect 574738 348372 574744 348384
rect 574796 348372 574802 348424
rect 132586 347760 132592 347812
rect 132644 347800 132650 347812
rect 133138 347800 133144 347812
rect 132644 347772 133144 347800
rect 132644 347760 132650 347772
rect 133138 347760 133144 347772
rect 133196 347800 133202 347812
rect 176654 347800 176660 347812
rect 133196 347772 176660 347800
rect 133196 347760 133202 347772
rect 176654 347760 176660 347772
rect 176712 347760 176718 347812
rect 49418 347012 49424 347064
rect 49476 347052 49482 347064
rect 179230 347052 179236 347064
rect 49476 347024 179236 347052
rect 49476 347012 49482 347024
rect 179230 347012 179236 347024
rect 179288 347012 179294 347064
rect 295426 347012 295432 347064
rect 295484 347052 295490 347064
rect 295794 347052 295800 347064
rect 295484 347024 295800 347052
rect 295484 347012 295490 347024
rect 295794 347012 295800 347024
rect 295852 347052 295858 347064
rect 300762 347052 300768 347064
rect 295852 347024 300768 347052
rect 295852 347012 295858 347024
rect 300762 347012 300768 347024
rect 300820 347052 300826 347064
rect 311250 347052 311256 347064
rect 300820 347024 311256 347052
rect 300820 347012 300826 347024
rect 311250 347012 311256 347024
rect 311308 347012 311314 347064
rect 355318 347012 355324 347064
rect 355376 347052 355382 347064
rect 437474 347052 437480 347064
rect 355376 347024 437480 347052
rect 355376 347012 355382 347024
rect 437474 347012 437480 347024
rect 437532 347012 437538 347064
rect 3326 345652 3332 345704
rect 3384 345692 3390 345704
rect 44818 345692 44824 345704
rect 3384 345664 44824 345692
rect 3384 345652 3390 345664
rect 44818 345652 44824 345664
rect 44876 345692 44882 345704
rect 118510 345692 118516 345704
rect 44876 345664 118516 345692
rect 44876 345652 44882 345664
rect 118510 345652 118516 345664
rect 118568 345652 118574 345704
rect 130470 345652 130476 345704
rect 130528 345692 130534 345704
rect 173710 345692 173716 345704
rect 130528 345664 173716 345692
rect 130528 345652 130534 345664
rect 173710 345652 173716 345664
rect 173768 345692 173774 345704
rect 176654 345692 176660 345704
rect 173768 345664 176660 345692
rect 173768 345652 173774 345664
rect 176654 345652 176660 345664
rect 176712 345652 176718 345704
rect 295610 345652 295616 345704
rect 295668 345692 295674 345704
rect 318610 345692 318616 345704
rect 295668 345664 318616 345692
rect 295668 345652 295674 345664
rect 318610 345652 318616 345664
rect 318668 345692 318674 345704
rect 534166 345692 534172 345704
rect 318668 345664 534172 345692
rect 318668 345652 318674 345664
rect 534166 345652 534172 345664
rect 534224 345652 534230 345704
rect 118510 344972 118516 345024
rect 118568 345012 118574 345024
rect 178678 345012 178684 345024
rect 118568 344984 178684 345012
rect 118568 344972 118574 344984
rect 178678 344972 178684 344984
rect 178736 344972 178742 345024
rect 295426 342864 295432 342916
rect 295484 342904 295490 342916
rect 296806 342904 296812 342916
rect 295484 342876 296812 342904
rect 295484 342864 295490 342876
rect 296806 342864 296812 342876
rect 296864 342904 296870 342916
rect 299934 342904 299940 342916
rect 296864 342876 299940 342904
rect 296864 342864 296870 342876
rect 299934 342864 299940 342876
rect 299992 342864 299998 342916
rect 359458 342184 359464 342236
rect 359516 342224 359522 342236
rect 502978 342224 502984 342236
rect 359516 342196 502984 342224
rect 359516 342184 359522 342196
rect 502978 342184 502984 342196
rect 503036 342184 503042 342236
rect 359458 341572 359464 341624
rect 359516 341612 359522 341624
rect 360010 341612 360016 341624
rect 359516 341584 360016 341612
rect 359516 341572 359522 341584
rect 360010 341572 360016 341584
rect 360068 341572 360074 341624
rect 78582 341504 78588 341556
rect 78640 341544 78646 341556
rect 132494 341544 132500 341556
rect 78640 341516 132500 341544
rect 78640 341504 78646 341516
rect 132494 341504 132500 341516
rect 132552 341504 132558 341556
rect 174998 340824 175004 340876
rect 175056 340864 175062 340876
rect 176654 340864 176660 340876
rect 175056 340836 176660 340864
rect 175056 340824 175062 340836
rect 176654 340824 176660 340836
rect 176712 340824 176718 340876
rect 295426 340824 295432 340876
rect 295484 340864 295490 340876
rect 311802 340864 311808 340876
rect 295484 340836 311808 340864
rect 295484 340824 295490 340836
rect 311802 340824 311808 340836
rect 311860 340824 311866 340876
rect 68646 340144 68652 340196
rect 68704 340184 68710 340196
rect 175918 340184 175924 340196
rect 68704 340156 175924 340184
rect 68704 340144 68710 340156
rect 175918 340144 175924 340156
rect 175976 340144 175982 340196
rect 311802 340144 311808 340196
rect 311860 340184 311866 340196
rect 344278 340184 344284 340196
rect 311860 340156 344284 340184
rect 311860 340144 311866 340156
rect 344278 340144 344284 340156
rect 344336 340144 344342 340196
rect 362218 340144 362224 340196
rect 362276 340184 362282 340196
rect 528554 340184 528560 340196
rect 362276 340156 528560 340184
rect 362276 340144 362282 340156
rect 528554 340144 528560 340156
rect 528612 340144 528618 340196
rect 295426 339396 295432 339448
rect 295484 339436 295490 339448
rect 301038 339436 301044 339448
rect 295484 339408 301044 339436
rect 295484 339396 295490 339408
rect 301038 339396 301044 339408
rect 301096 339436 301102 339448
rect 301314 339436 301320 339448
rect 301096 339408 301320 339436
rect 301096 339396 301102 339408
rect 301314 339396 301320 339408
rect 301372 339396 301378 339448
rect 301314 338784 301320 338836
rect 301372 338824 301378 338836
rect 325234 338824 325240 338836
rect 301372 338796 325240 338824
rect 301372 338784 301378 338796
rect 325234 338784 325240 338796
rect 325292 338784 325298 338836
rect 295978 338716 295984 338768
rect 296036 338756 296042 338768
rect 538398 338756 538404 338768
rect 296036 338728 538404 338756
rect 296036 338716 296042 338728
rect 538398 338716 538404 338728
rect 538456 338716 538462 338768
rect 175090 338104 175096 338156
rect 175148 338144 175154 338156
rect 176654 338144 176660 338156
rect 175148 338116 176660 338144
rect 175148 338104 175154 338116
rect 176654 338104 176660 338116
rect 176712 338104 176718 338156
rect 49510 337356 49516 337408
rect 49568 337396 49574 337408
rect 122926 337396 122932 337408
rect 49568 337368 122932 337396
rect 49568 337356 49574 337368
rect 122926 337356 122932 337368
rect 122984 337396 122990 337408
rect 174998 337396 175004 337408
rect 122984 337368 175004 337396
rect 122984 337356 122990 337368
rect 174998 337356 175004 337368
rect 175056 337356 175062 337408
rect 299934 335996 299940 336048
rect 299992 336036 299998 336048
rect 401594 336036 401600 336048
rect 299992 336008 401600 336036
rect 299992 335996 299998 336008
rect 401594 335996 401600 336008
rect 401652 335996 401658 336048
rect 371878 334636 371884 334688
rect 371936 334676 371942 334688
rect 396074 334676 396080 334688
rect 371936 334648 396080 334676
rect 371936 334636 371942 334648
rect 396074 334636 396080 334648
rect 396132 334636 396138 334688
rect 477954 334636 477960 334688
rect 478012 334676 478018 334688
rect 552014 334676 552020 334688
rect 478012 334648 552020 334676
rect 478012 334636 478018 334648
rect 552014 334636 552020 334648
rect 552072 334636 552078 334688
rect 175182 334568 175188 334620
rect 175240 334608 175246 334620
rect 176654 334608 176660 334620
rect 175240 334580 176660 334608
rect 175240 334568 175246 334580
rect 176654 334568 176660 334580
rect 176712 334568 176718 334620
rect 295702 334568 295708 334620
rect 295760 334608 295766 334620
rect 365254 334608 365260 334620
rect 295760 334580 365260 334608
rect 295760 334568 295766 334580
rect 365254 334568 365260 334580
rect 365312 334568 365318 334620
rect 379238 334568 379244 334620
rect 379296 334608 379302 334620
rect 512638 334608 512644 334620
rect 379296 334580 512644 334608
rect 379296 334568 379302 334580
rect 512638 334568 512644 334580
rect 512696 334568 512702 334620
rect 401594 333956 401600 334008
rect 401652 333996 401658 334008
rect 477494 333996 477500 334008
rect 401652 333968 477500 333996
rect 401652 333956 401658 333968
rect 477494 333956 477500 333968
rect 477552 333996 477558 334008
rect 477954 333996 477960 334008
rect 477552 333968 477960 333996
rect 477552 333956 477558 333968
rect 477954 333956 477960 333968
rect 478012 333956 478018 334008
rect 169754 333888 169760 333940
rect 169812 333928 169818 333940
rect 170950 333928 170956 333940
rect 169812 333900 170956 333928
rect 169812 333888 169818 333900
rect 170950 333888 170956 333900
rect 171008 333928 171014 333940
rect 176654 333928 176660 333940
rect 171008 333900 176660 333928
rect 171008 333888 171014 333900
rect 176654 333888 176660 333900
rect 176712 333888 176718 333940
rect 130654 333276 130660 333328
rect 130712 333316 130718 333328
rect 169754 333316 169760 333328
rect 130712 333288 169760 333316
rect 130712 333276 130718 333288
rect 169754 333276 169760 333288
rect 169812 333276 169818 333328
rect 295426 333276 295432 333328
rect 295484 333316 295490 333328
rect 353938 333316 353944 333328
rect 295484 333288 353944 333316
rect 295484 333276 295490 333288
rect 353938 333276 353944 333288
rect 353996 333276 354002 333328
rect 66898 333208 66904 333260
rect 66956 333248 66962 333260
rect 149054 333248 149060 333260
rect 66956 333220 149060 333248
rect 66956 333208 66962 333220
rect 149054 333208 149060 333220
rect 149112 333208 149118 333260
rect 304442 333208 304448 333260
rect 304500 333248 304506 333260
rect 513374 333248 513380 333260
rect 304500 333220 513380 333248
rect 304500 333208 304506 333220
rect 513374 333208 513380 333220
rect 513432 333208 513438 333260
rect 106918 331848 106924 331900
rect 106976 331888 106982 331900
rect 175182 331888 175188 331900
rect 106976 331860 175188 331888
rect 106976 331848 106982 331860
rect 175182 331848 175188 331860
rect 175240 331848 175246 331900
rect 355410 331848 355416 331900
rect 355468 331888 355474 331900
rect 441614 331888 441620 331900
rect 355468 331860 441620 331888
rect 355468 331848 355474 331860
rect 441614 331848 441620 331860
rect 441672 331848 441678 331900
rect 293862 331236 293868 331288
rect 293920 331276 293926 331288
rect 337378 331276 337384 331288
rect 293920 331248 337384 331276
rect 293920 331236 293926 331248
rect 337378 331236 337384 331248
rect 337436 331236 337442 331288
rect 295426 330488 295432 330540
rect 295484 330528 295490 330540
rect 300946 330528 300952 330540
rect 295484 330500 300952 330528
rect 295484 330488 295490 330500
rect 300946 330488 300952 330500
rect 301004 330528 301010 330540
rect 301314 330528 301320 330540
rect 301004 330500 301320 330528
rect 301004 330488 301010 330500
rect 301314 330488 301320 330500
rect 301372 330488 301378 330540
rect 58986 329060 58992 329112
rect 59044 329100 59050 329112
rect 74626 329100 74632 329112
rect 59044 329072 74632 329100
rect 59044 329060 59050 329072
rect 74626 329060 74632 329072
rect 74684 329100 74690 329112
rect 75270 329100 75276 329112
rect 74684 329072 75276 329100
rect 74684 329060 74690 329072
rect 75270 329060 75276 329072
rect 75328 329060 75334 329112
rect 301314 329060 301320 329112
rect 301372 329100 301378 329112
rect 440234 329100 440240 329112
rect 301372 329072 440240 329100
rect 301372 329060 301378 329072
rect 440234 329060 440240 329072
rect 440292 329060 440298 329112
rect 75270 328448 75276 328500
rect 75328 328488 75334 328500
rect 134518 328488 134524 328500
rect 75328 328460 134524 328488
rect 75328 328448 75334 328460
rect 134518 328448 134524 328460
rect 134576 328448 134582 328500
rect 440234 328380 440240 328432
rect 440292 328420 440298 328432
rect 440878 328420 440884 328432
rect 440292 328392 440884 328420
rect 440292 328380 440298 328392
rect 440878 328380 440884 328392
rect 440936 328420 440942 328432
rect 543734 328420 543740 328432
rect 440936 328392 543740 328420
rect 440936 328380 440942 328392
rect 543734 328380 543740 328392
rect 543792 328380 543798 328432
rect 295518 327700 295524 327752
rect 295576 327740 295582 327752
rect 310422 327740 310428 327752
rect 295576 327712 310428 327740
rect 295576 327700 295582 327712
rect 310422 327700 310428 327712
rect 310480 327700 310486 327752
rect 293126 327020 293132 327072
rect 293184 327060 293190 327072
rect 310330 327060 310336 327072
rect 293184 327032 310336 327060
rect 293184 327020 293190 327032
rect 310330 327020 310336 327032
rect 310388 327020 310394 327072
rect 310330 326408 310336 326460
rect 310388 326448 310394 326460
rect 348418 326448 348424 326460
rect 310388 326420 348424 326448
rect 310388 326408 310394 326420
rect 348418 326408 348424 326420
rect 348476 326408 348482 326460
rect 296622 326340 296628 326392
rect 296680 326380 296686 326392
rect 537110 326380 537116 326392
rect 296680 326352 537116 326380
rect 296680 326340 296686 326352
rect 537110 326340 537116 326352
rect 537168 326340 537174 326392
rect 173250 325660 173256 325712
rect 173308 325700 173314 325712
rect 176654 325700 176660 325712
rect 173308 325672 176660 325700
rect 173308 325660 173314 325672
rect 176654 325660 176660 325672
rect 176712 325660 176718 325712
rect 310330 324912 310336 324964
rect 310388 324952 310394 324964
rect 391198 324952 391204 324964
rect 310388 324924 391204 324952
rect 310388 324912 310394 324924
rect 391198 324912 391204 324924
rect 391256 324912 391262 324964
rect 337930 323552 337936 323604
rect 337988 323592 337994 323604
rect 458174 323592 458180 323604
rect 337988 323564 458180 323592
rect 337988 323552 337994 323564
rect 458174 323552 458180 323564
rect 458232 323552 458238 323604
rect 294322 322940 294328 322992
rect 294380 322980 294386 322992
rect 337930 322980 337936 322992
rect 294380 322952 337936 322980
rect 294380 322940 294386 322952
rect 337930 322940 337936 322952
rect 337988 322940 337994 322992
rect 81526 322872 81532 322924
rect 81584 322912 81590 322924
rect 82814 322912 82820 322924
rect 81584 322884 82820 322912
rect 81584 322872 81590 322884
rect 82814 322872 82820 322884
rect 82872 322912 82878 322924
rect 146294 322912 146300 322924
rect 82872 322884 146300 322912
rect 82872 322872 82878 322884
rect 146294 322872 146300 322884
rect 146352 322872 146358 322924
rect 300210 322192 300216 322244
rect 300268 322232 300274 322244
rect 369854 322232 369860 322244
rect 300268 322204 369860 322232
rect 300268 322192 300274 322204
rect 369854 322192 369860 322204
rect 369912 322192 369918 322244
rect 370498 322192 370504 322244
rect 370556 322232 370562 322244
rect 434714 322232 434720 322244
rect 370556 322204 434720 322232
rect 370556 322192 370562 322204
rect 434714 322192 434720 322204
rect 434772 322192 434778 322244
rect 438762 322192 438768 322244
rect 438820 322232 438826 322244
rect 509234 322232 509240 322244
rect 438820 322204 509240 322232
rect 438820 322192 438826 322204
rect 509234 322192 509240 322204
rect 509292 322192 509298 322244
rect 413278 321648 413284 321700
rect 413336 321688 413342 321700
rect 420178 321688 420184 321700
rect 413336 321660 420184 321688
rect 413336 321648 413342 321660
rect 420178 321648 420184 321660
rect 420236 321648 420242 321700
rect 175182 321580 175188 321632
rect 175240 321620 175246 321632
rect 177574 321620 177580 321632
rect 175240 321592 177580 321620
rect 175240 321580 175246 321592
rect 177574 321580 177580 321592
rect 177632 321620 177638 321632
rect 177758 321620 177764 321632
rect 177632 321592 177764 321620
rect 177632 321580 177638 321592
rect 177758 321580 177764 321592
rect 177816 321580 177822 321632
rect 295334 321512 295340 321564
rect 295392 321552 295398 321564
rect 305730 321552 305736 321564
rect 295392 321524 305736 321552
rect 295392 321512 295398 321524
rect 305730 321512 305736 321524
rect 305788 321552 305794 321564
rect 306282 321552 306288 321564
rect 305788 321524 306288 321552
rect 305788 321512 305794 321524
rect 306282 321512 306288 321524
rect 306340 321512 306346 321564
rect 310422 321512 310428 321564
rect 310480 321552 310486 321564
rect 393958 321552 393964 321564
rect 310480 321524 393964 321552
rect 310480 321512 310486 321524
rect 393958 321512 393964 321524
rect 394016 321512 394022 321564
rect 305730 320832 305736 320884
rect 305788 320872 305794 320884
rect 319622 320872 319628 320884
rect 305788 320844 319628 320872
rect 305788 320832 305794 320844
rect 319622 320832 319628 320844
rect 319680 320832 319686 320884
rect 359458 320832 359464 320884
rect 359516 320872 359522 320884
rect 448514 320872 448520 320884
rect 359516 320844 448520 320872
rect 359516 320832 359522 320844
rect 448514 320832 448520 320844
rect 448572 320832 448578 320884
rect 3142 320084 3148 320136
rect 3200 320124 3206 320136
rect 59262 320124 59268 320136
rect 3200 320096 59268 320124
rect 3200 320084 3206 320096
rect 59262 320084 59268 320096
rect 59320 320084 59326 320136
rect 367738 319472 367744 319524
rect 367796 319512 367802 319524
rect 394694 319512 394700 319524
rect 367796 319484 394700 319512
rect 367796 319472 367802 319484
rect 394694 319472 394700 319484
rect 394752 319472 394758 319524
rect 59262 319404 59268 319456
rect 59320 319444 59326 319456
rect 87598 319444 87604 319456
rect 59320 319416 87604 319444
rect 59320 319404 59326 319416
rect 87598 319404 87604 319416
rect 87656 319404 87662 319456
rect 313366 319404 313372 319456
rect 313424 319444 313430 319456
rect 314562 319444 314568 319456
rect 313424 319416 314568 319444
rect 313424 319404 313430 319416
rect 314562 319404 314568 319416
rect 314620 319444 314626 319456
rect 325050 319444 325056 319456
rect 314620 319416 325056 319444
rect 314620 319404 314626 319416
rect 325050 319404 325056 319416
rect 325108 319404 325114 319456
rect 379514 319404 379520 319456
rect 379572 319444 379578 319456
rect 483014 319444 483020 319456
rect 379572 319416 483020 319444
rect 379572 319404 379578 319416
rect 483014 319404 483020 319416
rect 483072 319404 483078 319456
rect 295334 318792 295340 318844
rect 295392 318832 295398 318844
rect 313366 318832 313372 318844
rect 295392 318804 313372 318832
rect 295392 318792 295398 318804
rect 313366 318792 313372 318804
rect 313424 318792 313430 318844
rect 447134 318792 447140 318844
rect 447192 318832 447198 318844
rect 466454 318832 466460 318844
rect 447192 318804 466460 318832
rect 447192 318792 447198 318804
rect 466454 318792 466460 318804
rect 466512 318792 466518 318844
rect 81434 318724 81440 318776
rect 81492 318764 81498 318776
rect 106274 318764 106280 318776
rect 81492 318736 106280 318764
rect 81492 318724 81498 318736
rect 106274 318724 106280 318736
rect 106332 318764 106338 318776
rect 106918 318764 106924 318776
rect 106332 318736 106924 318764
rect 106332 318724 106338 318736
rect 106918 318724 106924 318736
rect 106976 318724 106982 318776
rect 33042 318044 33048 318096
rect 33100 318084 33106 318096
rect 136726 318084 136732 318096
rect 33100 318056 136732 318084
rect 33100 318044 33106 318056
rect 136726 318044 136732 318056
rect 136784 318044 136790 318096
rect 147582 318044 147588 318096
rect 147640 318084 147646 318096
rect 173250 318084 173256 318096
rect 147640 318056 173256 318084
rect 147640 318044 147646 318056
rect 173250 318044 173256 318056
rect 173308 318044 173314 318096
rect 379146 318044 379152 318096
rect 379204 318084 379210 318096
rect 447134 318084 447140 318096
rect 379204 318056 447140 318084
rect 379204 318044 379210 318056
rect 447134 318044 447140 318056
rect 447192 318044 447198 318096
rect 136726 317432 136732 317484
rect 136784 317472 136790 317484
rect 147582 317472 147588 317484
rect 136784 317444 147588 317472
rect 136784 317432 136790 317444
rect 147582 317432 147588 317444
rect 147640 317432 147646 317484
rect 177942 317364 177948 317416
rect 178000 317404 178006 317416
rect 179138 317404 179144 317416
rect 178000 317376 179144 317404
rect 178000 317364 178006 317376
rect 179138 317364 179144 317376
rect 179196 317364 179202 317416
rect 345842 316820 345848 316872
rect 345900 316860 345906 316872
rect 377398 316860 377404 316872
rect 345900 316832 377404 316860
rect 345900 316820 345906 316832
rect 377398 316820 377404 316832
rect 377456 316820 377462 316872
rect 304534 316752 304540 316804
rect 304592 316792 304598 316804
rect 362954 316792 362960 316804
rect 304592 316764 362960 316792
rect 304592 316752 304598 316764
rect 362954 316752 362960 316764
rect 363012 316752 363018 316804
rect 59170 316684 59176 316736
rect 59228 316724 59234 316736
rect 105538 316724 105544 316736
rect 59228 316696 105544 316724
rect 59228 316684 59234 316696
rect 105538 316684 105544 316696
rect 105596 316684 105602 316736
rect 295334 316684 295340 316736
rect 295392 316724 295398 316736
rect 299290 316724 299296 316736
rect 295392 316696 299296 316724
rect 295392 316684 295398 316696
rect 299290 316684 299296 316696
rect 299348 316684 299354 316736
rect 338022 316684 338028 316736
rect 338080 316724 338086 316736
rect 443086 316724 443092 316736
rect 338080 316696 443092 316724
rect 338080 316684 338086 316696
rect 443086 316684 443092 316696
rect 443144 316684 443150 316736
rect 362954 316004 362960 316056
rect 363012 316044 363018 316056
rect 364242 316044 364248 316056
rect 363012 316016 364248 316044
rect 363012 316004 363018 316016
rect 364242 316004 364248 316016
rect 364300 316044 364306 316056
rect 415578 316044 415584 316056
rect 364300 316016 415584 316044
rect 364300 316004 364306 316016
rect 415578 316004 415584 316016
rect 415636 316004 415642 316056
rect 299290 315936 299296 315988
rect 299348 315976 299354 315988
rect 304994 315976 305000 315988
rect 299348 315948 305000 315976
rect 299348 315936 299354 315948
rect 304994 315936 305000 315948
rect 305052 315936 305058 315988
rect 49602 315256 49608 315308
rect 49660 315296 49666 315308
rect 59262 315296 59268 315308
rect 49660 315268 59268 315296
rect 49660 315256 49666 315268
rect 59262 315256 59268 315268
rect 59320 315256 59326 315308
rect 87598 315256 87604 315308
rect 87656 315296 87662 315308
rect 116762 315296 116768 315308
rect 87656 315268 116768 315296
rect 87656 315256 87662 315268
rect 116762 315256 116768 315268
rect 116820 315256 116826 315308
rect 304994 315256 305000 315308
rect 305052 315296 305058 315308
rect 373258 315296 373264 315308
rect 305052 315268 373264 315296
rect 305052 315256 305058 315268
rect 373258 315256 373264 315268
rect 373316 315256 373322 315308
rect 452562 315256 452568 315308
rect 452620 315296 452626 315308
rect 556798 315296 556804 315308
rect 452620 315268 556804 315296
rect 452620 315256 452626 315268
rect 556798 315256 556804 315268
rect 556856 315256 556862 315308
rect 59262 314644 59268 314696
rect 59320 314684 59326 314696
rect 157242 314684 157248 314696
rect 59320 314656 157248 314684
rect 59320 314644 59326 314656
rect 157242 314644 157248 314656
rect 157300 314684 157306 314696
rect 179322 314684 179328 314696
rect 157300 314656 179328 314684
rect 157300 314644 157306 314656
rect 179322 314644 179328 314656
rect 179380 314644 179386 314696
rect 451274 314684 451280 314696
rect 387720 314656 451280 314684
rect 295334 314576 295340 314628
rect 295392 314616 295398 314628
rect 317598 314616 317604 314628
rect 295392 314588 317604 314616
rect 295392 314576 295398 314588
rect 317598 314576 317604 314588
rect 317656 314616 317662 314628
rect 318518 314616 318524 314628
rect 317656 314588 318524 314616
rect 317656 314576 317662 314588
rect 318518 314576 318524 314588
rect 318576 314576 318582 314628
rect 320818 314576 320824 314628
rect 320876 314616 320882 314628
rect 386506 314616 386512 314628
rect 320876 314588 386512 314616
rect 320876 314576 320882 314588
rect 386506 314576 386512 314588
rect 386564 314616 386570 314628
rect 387720 314616 387748 314656
rect 451274 314644 451280 314656
rect 451332 314684 451338 314696
rect 452562 314684 452568 314696
rect 451332 314656 452568 314684
rect 451332 314644 451338 314656
rect 452562 314644 452568 314656
rect 452620 314644 452626 314696
rect 386564 314588 387748 314616
rect 386564 314576 386570 314588
rect 34422 313896 34428 313948
rect 34480 313936 34486 313948
rect 124214 313936 124220 313948
rect 34480 313908 124220 313936
rect 34480 313896 34486 313908
rect 124214 313896 124220 313908
rect 124272 313896 124278 313948
rect 296070 313896 296076 313948
rect 296128 313936 296134 313948
rect 306466 313936 306472 313948
rect 296128 313908 306472 313936
rect 296128 313896 296134 313908
rect 306466 313896 306472 313908
rect 306524 313896 306530 313948
rect 318518 313896 318524 313948
rect 318576 313936 318582 313948
rect 386322 313936 386328 313948
rect 318576 313908 386328 313936
rect 318576 313896 318582 313908
rect 386322 313896 386328 313908
rect 386380 313896 386386 313948
rect 385678 313420 385684 313472
rect 385736 313460 385742 313472
rect 389174 313460 389180 313472
rect 385736 313432 389180 313460
rect 385736 313420 385742 313432
rect 389174 313420 389180 313432
rect 389232 313420 389238 313472
rect 57790 313216 57796 313268
rect 57848 313256 57854 313268
rect 109034 313256 109040 313268
rect 57848 313228 109040 313256
rect 57848 313216 57854 313228
rect 109034 313216 109040 313228
rect 109092 313216 109098 313268
rect 109034 312604 109040 312656
rect 109092 312644 109098 312656
rect 109678 312644 109684 312656
rect 109092 312616 109684 312644
rect 109092 312604 109098 312616
rect 109678 312604 109684 312616
rect 109736 312604 109742 312656
rect 420178 312604 420184 312656
rect 420236 312644 420242 312656
rect 440970 312644 440976 312656
rect 420236 312616 440976 312644
rect 420236 312604 420242 312616
rect 440970 312604 440976 312616
rect 441028 312604 441034 312656
rect 170674 312536 170680 312588
rect 170732 312576 170738 312588
rect 171042 312576 171048 312588
rect 170732 312548 171048 312576
rect 170732 312536 170738 312548
rect 171042 312536 171048 312548
rect 171100 312576 171106 312588
rect 176654 312576 176660 312588
rect 171100 312548 176660 312576
rect 171100 312536 171106 312548
rect 176654 312536 176660 312548
rect 176712 312536 176718 312588
rect 295334 312536 295340 312588
rect 295392 312576 295398 312588
rect 304994 312576 305000 312588
rect 295392 312548 305000 312576
rect 295392 312536 295398 312548
rect 304994 312536 305000 312548
rect 305052 312536 305058 312588
rect 360838 312536 360844 312588
rect 360896 312576 360902 312588
rect 430574 312576 430580 312588
rect 360896 312548 430580 312576
rect 360896 312536 360902 312548
rect 430574 312536 430580 312548
rect 430632 312536 430638 312588
rect 450538 312536 450544 312588
rect 450596 312576 450602 312588
rect 458174 312576 458180 312588
rect 450596 312548 458180 312576
rect 450596 312536 450602 312548
rect 458174 312536 458180 312548
rect 458232 312536 458238 312588
rect 304994 311856 305000 311908
rect 305052 311896 305058 311908
rect 372614 311896 372620 311908
rect 305052 311868 372620 311896
rect 305052 311856 305058 311868
rect 372614 311856 372620 311868
rect 372672 311856 372678 311908
rect 458174 311856 458180 311908
rect 458232 311896 458238 311908
rect 579982 311896 579988 311908
rect 458232 311868 579988 311896
rect 458232 311856 458238 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 457438 311788 457444 311840
rect 457496 311828 457502 311840
rect 460934 311828 460940 311840
rect 457496 311800 460940 311828
rect 457496 311788 457502 311800
rect 460934 311788 460940 311800
rect 460992 311788 460998 311840
rect 79318 311176 79324 311228
rect 79376 311216 79382 311228
rect 157978 311216 157984 311228
rect 79376 311188 157984 311216
rect 79376 311176 79382 311188
rect 157978 311176 157984 311188
rect 158036 311176 158042 311228
rect 43806 311108 43812 311160
rect 43864 311148 43870 311160
rect 132494 311148 132500 311160
rect 43864 311120 132500 311148
rect 43864 311108 43870 311120
rect 132494 311108 132500 311120
rect 132552 311108 132558 311160
rect 85574 310972 85580 311024
rect 85632 311012 85638 311024
rect 86218 311012 86224 311024
rect 85632 310984 86224 311012
rect 85632 310972 85638 310984
rect 86218 310972 86224 310984
rect 86276 310972 86282 311024
rect 86218 310496 86224 310548
rect 86276 310536 86282 310548
rect 170398 310536 170404 310548
rect 86276 310508 170404 310536
rect 86276 310496 86282 310508
rect 170398 310496 170404 310508
rect 170456 310496 170462 310548
rect 295334 310428 295340 310480
rect 295392 310468 295398 310480
rect 307846 310468 307852 310480
rect 295392 310440 307852 310468
rect 295392 310428 295398 310440
rect 307846 310428 307852 310440
rect 307904 310468 307910 310480
rect 308950 310468 308956 310480
rect 307904 310440 308956 310468
rect 307904 310428 307910 310440
rect 308950 310428 308956 310440
rect 309008 310428 309014 310480
rect 173342 310224 173348 310276
rect 173400 310264 173406 310276
rect 173802 310264 173808 310276
rect 173400 310236 173808 310264
rect 173400 310224 173406 310236
rect 173802 310224 173808 310236
rect 173860 310264 173866 310276
rect 176654 310264 176660 310276
rect 173860 310236 176660 310264
rect 173860 310224 173866 310236
rect 176654 310224 176660 310236
rect 176712 310224 176718 310276
rect 386322 309884 386328 309936
rect 386380 309924 386386 309936
rect 395338 309924 395344 309936
rect 386380 309896 395344 309924
rect 386380 309884 386386 309896
rect 395338 309884 395344 309896
rect 395396 309884 395402 309936
rect 308950 309816 308956 309868
rect 309008 309856 309014 309868
rect 360286 309856 360292 309868
rect 309008 309828 360292 309856
rect 309008 309816 309014 309828
rect 360286 309816 360292 309828
rect 360344 309816 360350 309868
rect 372614 309816 372620 309868
rect 372672 309856 372678 309868
rect 391198 309856 391204 309868
rect 372672 309828 391204 309856
rect 372672 309816 372678 309828
rect 391198 309816 391204 309828
rect 391256 309816 391262 309868
rect 41230 309748 41236 309800
rect 41288 309788 41294 309800
rect 68278 309788 68284 309800
rect 41288 309760 68284 309788
rect 41288 309748 41294 309760
rect 68278 309748 68284 309760
rect 68336 309748 68342 309800
rect 326430 309748 326436 309800
rect 326488 309788 326494 309800
rect 419534 309788 419540 309800
rect 326488 309760 419540 309788
rect 326488 309748 326494 309760
rect 419534 309748 419540 309760
rect 419592 309748 419598 309800
rect 360286 309136 360292 309188
rect 360344 309176 360350 309188
rect 361482 309176 361488 309188
rect 360344 309148 361488 309176
rect 360344 309136 360350 309148
rect 361482 309136 361488 309148
rect 361540 309176 361546 309188
rect 384298 309176 384304 309188
rect 361540 309148 384304 309176
rect 361540 309136 361546 309148
rect 384298 309136 384304 309148
rect 384356 309136 384362 309188
rect 419534 309068 419540 309120
rect 419592 309108 419598 309120
rect 420178 309108 420184 309120
rect 419592 309080 420184 309108
rect 419592 309068 419598 309080
rect 420178 309068 420184 309080
rect 420236 309108 420242 309120
rect 436922 309108 436928 309120
rect 420236 309080 436928 309108
rect 420236 309068 420242 309080
rect 436922 309068 436928 309080
rect 436980 309108 436986 309120
rect 437382 309108 437388 309120
rect 436980 309080 437388 309108
rect 436980 309068 436986 309080
rect 437382 309068 437388 309080
rect 437440 309068 437446 309120
rect 39758 308456 39764 308508
rect 39816 308496 39822 308508
rect 69014 308496 69020 308508
rect 39816 308468 69020 308496
rect 39816 308456 39822 308468
rect 69014 308456 69020 308468
rect 69072 308456 69078 308508
rect 93762 308456 93768 308508
rect 93820 308496 93826 308508
rect 114554 308496 114560 308508
rect 93820 308468 114560 308496
rect 93820 308456 93826 308468
rect 114554 308456 114560 308468
rect 114612 308456 114618 308508
rect 436922 308456 436928 308508
rect 436980 308496 436986 308508
rect 465074 308496 465080 308508
rect 436980 308468 465080 308496
rect 436980 308456 436986 308468
rect 465074 308456 465080 308468
rect 465132 308456 465138 308508
rect 48038 308388 48044 308440
rect 48096 308428 48102 308440
rect 131850 308428 131856 308440
rect 48096 308400 131856 308428
rect 48096 308388 48102 308400
rect 131850 308388 131856 308400
rect 131908 308388 131914 308440
rect 458358 308388 458364 308440
rect 458416 308428 458422 308440
rect 575474 308428 575480 308440
rect 458416 308400 575480 308428
rect 458416 308388 458422 308400
rect 575474 308388 575480 308400
rect 575532 308388 575538 308440
rect 73062 307776 73068 307828
rect 73120 307816 73126 307828
rect 75914 307816 75920 307828
rect 73120 307788 75920 307816
rect 73120 307776 73126 307788
rect 75914 307776 75920 307788
rect 75972 307776 75978 307828
rect 295334 307776 295340 307828
rect 295392 307816 295398 307828
rect 303614 307816 303620 307828
rect 295392 307788 303620 307816
rect 295392 307776 295398 307788
rect 303614 307776 303620 307788
rect 303672 307816 303678 307828
rect 399478 307816 399484 307828
rect 303672 307788 399484 307816
rect 303672 307776 303678 307788
rect 399478 307776 399484 307788
rect 399536 307776 399542 307828
rect 434162 307776 434168 307828
rect 434220 307816 434226 307828
rect 458358 307816 458364 307828
rect 434220 307788 458364 307816
rect 434220 307776 434226 307788
rect 458358 307776 458364 307788
rect 458416 307776 458422 307828
rect 88426 307300 88432 307352
rect 88484 307340 88490 307352
rect 89714 307340 89720 307352
rect 88484 307312 89720 307340
rect 88484 307300 88490 307312
rect 89714 307300 89720 307312
rect 89772 307300 89778 307352
rect 379606 307164 379612 307216
rect 379664 307204 379670 307216
rect 386414 307204 386420 307216
rect 379664 307176 386420 307204
rect 379664 307164 379670 307176
rect 386414 307164 386420 307176
rect 386472 307164 386478 307216
rect 377490 307096 377496 307148
rect 377548 307136 377554 307148
rect 398834 307136 398840 307148
rect 377548 307108 398840 307136
rect 377548 307096 377554 307108
rect 398834 307096 398840 307108
rect 398892 307096 398898 307148
rect 300302 307028 300308 307080
rect 300360 307068 300366 307080
rect 441706 307068 441712 307080
rect 300360 307040 441712 307068
rect 300360 307028 300366 307040
rect 441706 307028 441712 307040
rect 441764 307028 441770 307080
rect 89714 306960 89720 307012
rect 89772 307000 89778 307012
rect 90358 307000 90364 307012
rect 89772 306972 90364 307000
rect 89772 306960 89778 306972
rect 90358 306960 90364 306972
rect 90416 306960 90422 307012
rect 80054 306688 80060 306740
rect 80112 306728 80118 306740
rect 83458 306728 83464 306740
rect 80112 306700 83464 306728
rect 80112 306688 80118 306700
rect 83458 306688 83464 306700
rect 83516 306688 83522 306740
rect 113266 306484 113272 306536
rect 113324 306524 113330 306536
rect 113818 306524 113824 306536
rect 113324 306496 113824 306524
rect 113324 306484 113330 306496
rect 113818 306484 113824 306496
rect 113876 306524 113882 306536
rect 159450 306524 159456 306536
rect 113876 306496 159456 306524
rect 113876 306484 113882 306496
rect 159450 306484 159456 306496
rect 159508 306484 159514 306536
rect 102134 306416 102140 306468
rect 102192 306456 102198 306468
rect 160922 306456 160928 306468
rect 102192 306428 160928 306456
rect 102192 306416 102198 306428
rect 160922 306416 160928 306428
rect 160980 306416 160986 306468
rect 90358 306348 90364 306400
rect 90416 306388 90422 306400
rect 152458 306388 152464 306400
rect 90416 306360 152464 306388
rect 90416 306348 90422 306360
rect 152458 306348 152464 306360
rect 152516 306348 152522 306400
rect 391198 306348 391204 306400
rect 391256 306388 391262 306400
rect 469214 306388 469220 306400
rect 391256 306360 469220 306388
rect 391256 306348 391262 306360
rect 469214 306348 469220 306360
rect 469272 306348 469278 306400
rect 172330 306076 172336 306128
rect 172388 306116 172394 306128
rect 176654 306116 176660 306128
rect 172388 306088 176660 306116
rect 172388 306076 172394 306088
rect 176654 306076 176660 306088
rect 176712 306076 176718 306128
rect 76650 305668 76656 305720
rect 76708 305708 76714 305720
rect 112530 305708 112536 305720
rect 76708 305680 112536 305708
rect 76708 305668 76714 305680
rect 112530 305668 112536 305680
rect 112588 305668 112594 305720
rect 121362 305668 121368 305720
rect 121420 305708 121426 305720
rect 172330 305708 172336 305720
rect 121420 305680 172336 305708
rect 121420 305668 121426 305680
rect 172330 305668 172336 305680
rect 172388 305668 172394 305720
rect 45370 305600 45376 305652
rect 45428 305640 45434 305652
rect 127066 305640 127072 305652
rect 45428 305612 127072 305640
rect 45428 305600 45434 305612
rect 127066 305600 127072 305612
rect 127124 305600 127130 305652
rect 410518 305600 410524 305652
rect 410576 305640 410582 305652
rect 448606 305640 448612 305652
rect 410576 305612 448612 305640
rect 410576 305600 410582 305612
rect 448606 305600 448612 305612
rect 448664 305600 448670 305652
rect 294046 305328 294052 305380
rect 294104 305368 294110 305380
rect 295334 305368 295340 305380
rect 294104 305340 295340 305368
rect 294104 305328 294110 305340
rect 295334 305328 295340 305340
rect 295392 305328 295398 305380
rect 88334 305056 88340 305108
rect 88392 305096 88398 305108
rect 88978 305096 88984 305108
rect 88392 305068 88984 305096
rect 88392 305056 88398 305068
rect 88978 305056 88984 305068
rect 89036 305096 89042 305108
rect 136082 305096 136088 305108
rect 89036 305068 136088 305096
rect 89036 305056 89042 305068
rect 136082 305056 136088 305068
rect 136140 305056 136146 305108
rect 404998 305056 405004 305108
rect 405056 305096 405062 305108
rect 455414 305096 455420 305108
rect 405056 305068 455420 305096
rect 405056 305056 405062 305068
rect 455414 305056 455420 305068
rect 455472 305056 455478 305108
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 120258 305028 120264 305040
rect 3292 305000 120264 305028
rect 3292 304988 3298 305000
rect 120258 304988 120264 305000
rect 120316 305028 120322 305040
rect 121362 305028 121368 305040
rect 120316 305000 121368 305028
rect 120316 304988 120322 305000
rect 121362 304988 121368 305000
rect 121420 304988 121426 305040
rect 409598 304988 409604 305040
rect 409656 305028 409662 305040
rect 463694 305028 463700 305040
rect 409656 305000 463700 305028
rect 409656 304988 409662 305000
rect 463694 304988 463700 305000
rect 463752 304988 463758 305040
rect 134518 304376 134524 304428
rect 134576 304416 134582 304428
rect 173250 304416 173256 304428
rect 134576 304388 173256 304416
rect 134576 304376 134582 304388
rect 173250 304376 173256 304388
rect 173308 304376 173314 304428
rect 114738 304308 114744 304360
rect 114796 304348 114802 304360
rect 173342 304348 173348 304360
rect 114796 304320 173348 304348
rect 114796 304308 114802 304320
rect 173342 304308 173348 304320
rect 173400 304308 173406 304360
rect 104986 304240 104992 304292
rect 105044 304280 105050 304292
rect 167730 304280 167736 304292
rect 105044 304252 167736 304280
rect 105044 304240 105050 304252
rect 167730 304240 167736 304252
rect 167788 304240 167794 304292
rect 295334 304240 295340 304292
rect 295392 304280 295398 304292
rect 441614 304280 441620 304292
rect 295392 304252 441620 304280
rect 295392 304240 295398 304252
rect 441614 304240 441620 304252
rect 441672 304240 441678 304292
rect 103514 303900 103520 303952
rect 103572 303940 103578 303952
rect 104986 303940 104992 303952
rect 103572 303912 104992 303940
rect 103572 303900 103578 303912
rect 104986 303900 104992 303912
rect 105044 303900 105050 303952
rect 429838 303900 429844 303952
rect 429896 303940 429902 303952
rect 430298 303940 430304 303952
rect 429896 303912 430304 303940
rect 429896 303900 429902 303912
rect 430298 303900 430304 303912
rect 430356 303940 430362 303952
rect 447134 303940 447140 303952
rect 430356 303912 447140 303940
rect 430356 303900 430362 303912
rect 447134 303900 447140 303912
rect 447192 303900 447198 303952
rect 98546 303832 98552 303884
rect 98604 303872 98610 303884
rect 98730 303872 98736 303884
rect 98604 303844 98736 303872
rect 98604 303832 98610 303844
rect 98730 303832 98736 303844
rect 98788 303872 98794 303884
rect 128998 303872 129004 303884
rect 98788 303844 129004 303872
rect 98788 303832 98794 303844
rect 128998 303832 129004 303844
rect 129056 303832 129062 303884
rect 406378 303832 406384 303884
rect 406436 303872 406442 303884
rect 442994 303872 443000 303884
rect 406436 303844 443000 303872
rect 406436 303832 406442 303844
rect 442994 303832 443000 303844
rect 443052 303832 443058 303884
rect 81434 303764 81440 303816
rect 81492 303804 81498 303816
rect 138658 303804 138664 303816
rect 81492 303776 138664 303804
rect 81492 303764 81498 303776
rect 138658 303764 138664 303776
rect 138716 303764 138722 303816
rect 417602 303764 417608 303816
rect 417660 303804 417666 303816
rect 458174 303804 458180 303816
rect 417660 303776 458180 303804
rect 417660 303764 417666 303776
rect 458174 303764 458180 303776
rect 458232 303764 458238 303816
rect 70486 303696 70492 303748
rect 70544 303736 70550 303748
rect 71038 303736 71044 303748
rect 70544 303708 71044 303736
rect 70544 303696 70550 303708
rect 71038 303696 71044 303708
rect 71096 303736 71102 303748
rect 153838 303736 153844 303748
rect 71096 303708 153844 303736
rect 71096 303696 71102 303708
rect 153838 303696 153844 303708
rect 153896 303696 153902 303748
rect 373718 303696 373724 303748
rect 373776 303736 373782 303748
rect 380894 303736 380900 303748
rect 373776 303708 380900 303736
rect 373776 303696 373782 303708
rect 380894 303696 380900 303708
rect 380952 303696 380958 303748
rect 399478 303696 399484 303748
rect 399536 303736 399542 303748
rect 444374 303736 444380 303748
rect 399536 303708 444380 303736
rect 399536 303696 399542 303708
rect 444374 303696 444380 303708
rect 444432 303696 444438 303748
rect 22738 303628 22744 303680
rect 22796 303668 22802 303680
rect 117866 303668 117872 303680
rect 22796 303640 117872 303668
rect 22796 303628 22802 303640
rect 117866 303628 117872 303640
rect 117924 303628 117930 303680
rect 362862 303628 362868 303680
rect 362920 303668 362926 303680
rect 389174 303668 389180 303680
rect 362920 303640 389180 303668
rect 362920 303628 362926 303640
rect 389174 303628 389180 303640
rect 389232 303628 389238 303680
rect 395338 303628 395344 303680
rect 395396 303668 395402 303680
rect 471974 303668 471980 303680
rect 395396 303640 471980 303668
rect 395396 303628 395402 303640
rect 471974 303628 471980 303640
rect 472032 303628 472038 303680
rect 295334 303560 295340 303612
rect 295392 303600 295398 303612
rect 300854 303600 300860 303612
rect 295392 303572 300860 303600
rect 295392 303560 295398 303572
rect 300854 303560 300860 303572
rect 300912 303560 300918 303612
rect 398098 303560 398104 303612
rect 398156 303600 398162 303612
rect 404998 303600 405004 303612
rect 398156 303572 405004 303600
rect 398156 303560 398162 303572
rect 404998 303560 405004 303572
rect 405056 303560 405062 303612
rect 111794 303016 111800 303068
rect 111852 303056 111858 303068
rect 128354 303056 128360 303068
rect 111852 303028 128360 303056
rect 111852 303016 111858 303028
rect 128354 303016 128360 303028
rect 128412 303016 128418 303068
rect 46842 302948 46848 303000
rect 46900 302988 46906 303000
rect 68738 302988 68744 303000
rect 46900 302960 68744 302988
rect 46900 302948 46906 302960
rect 68738 302948 68744 302960
rect 68796 302988 68802 303000
rect 102134 302988 102140 303000
rect 68796 302960 102140 302988
rect 68796 302948 68802 302960
rect 102134 302948 102140 302960
rect 102192 302948 102198 303000
rect 106182 302948 106188 303000
rect 106240 302988 106246 303000
rect 122834 302988 122840 303000
rect 106240 302960 122840 302988
rect 106240 302948 106246 302960
rect 122834 302948 122840 302960
rect 122892 302948 122898 303000
rect 300854 302948 300860 303000
rect 300912 302988 300918 303000
rect 356790 302988 356796 303000
rect 300912 302960 356796 302988
rect 300912 302948 300918 302960
rect 356790 302948 356796 302960
rect 356848 302948 356854 303000
rect 35710 302880 35716 302932
rect 35768 302920 35774 302932
rect 126422 302920 126428 302932
rect 35768 302892 126428 302920
rect 35768 302880 35774 302892
rect 126422 302880 126428 302892
rect 126480 302880 126486 302932
rect 297542 302880 297548 302932
rect 297600 302920 297606 302932
rect 304350 302920 304356 302932
rect 297600 302892 304356 302920
rect 297600 302880 297606 302892
rect 304350 302880 304356 302892
rect 304408 302920 304414 302932
rect 374730 302920 374736 302932
rect 304408 302892 374736 302920
rect 304408 302880 304414 302892
rect 374730 302880 374736 302892
rect 374788 302880 374794 302932
rect 403618 302540 403624 302592
rect 403676 302580 403682 302592
rect 459646 302580 459652 302592
rect 403676 302552 459652 302580
rect 403676 302540 403682 302552
rect 459646 302540 459652 302552
rect 459704 302540 459710 302592
rect 425882 302472 425888 302524
rect 425940 302512 425946 302524
rect 446398 302512 446404 302524
rect 425940 302484 446404 302512
rect 425940 302472 425946 302484
rect 446398 302472 446404 302484
rect 446456 302472 446462 302524
rect 428366 302404 428372 302456
rect 428424 302444 428430 302456
rect 429102 302444 429108 302456
rect 428424 302416 429108 302444
rect 428424 302404 428430 302416
rect 429102 302404 429108 302416
rect 429160 302444 429166 302456
rect 451366 302444 451372 302456
rect 429160 302416 451372 302444
rect 429160 302404 429166 302416
rect 451366 302404 451372 302416
rect 451424 302404 451430 302456
rect 360102 302336 360108 302388
rect 360160 302376 360166 302388
rect 385034 302376 385040 302388
rect 360160 302348 385040 302376
rect 360160 302336 360166 302348
rect 385034 302336 385040 302348
rect 385092 302376 385098 302388
rect 385770 302376 385776 302388
rect 385092 302348 385776 302376
rect 385092 302336 385098 302348
rect 385770 302336 385776 302348
rect 385828 302336 385834 302388
rect 440142 302336 440148 302388
rect 440200 302376 440206 302388
rect 470686 302376 470692 302388
rect 440200 302348 470692 302376
rect 440200 302336 440206 302348
rect 470686 302336 470692 302348
rect 470744 302336 470750 302388
rect 88426 302268 88432 302320
rect 88484 302308 88490 302320
rect 157978 302308 157984 302320
rect 88484 302280 157984 302308
rect 88484 302268 88490 302280
rect 157978 302268 157984 302280
rect 158036 302268 158042 302320
rect 376202 302268 376208 302320
rect 376260 302308 376266 302320
rect 423858 302308 423864 302320
rect 376260 302280 423864 302308
rect 376260 302268 376266 302280
rect 423858 302268 423864 302280
rect 423916 302308 423922 302320
rect 456794 302308 456800 302320
rect 423916 302280 456800 302308
rect 423916 302268 423922 302280
rect 456794 302268 456800 302280
rect 456852 302268 456858 302320
rect 90266 302200 90272 302252
rect 90324 302240 90330 302252
rect 162210 302240 162216 302252
rect 90324 302212 162216 302240
rect 90324 302200 90330 302212
rect 162210 302200 162216 302212
rect 162268 302200 162274 302252
rect 374730 302200 374736 302252
rect 374788 302240 374794 302252
rect 375282 302240 375288 302252
rect 374788 302212 375288 302240
rect 374788 302200 374794 302212
rect 375282 302200 375288 302212
rect 375340 302240 375346 302252
rect 407666 302240 407672 302252
rect 375340 302212 407672 302240
rect 375340 302200 375346 302212
rect 407666 302200 407672 302212
rect 407724 302200 407730 302252
rect 103606 301588 103612 301640
rect 103664 301628 103670 301640
rect 130654 301628 130660 301640
rect 103664 301600 130660 301628
rect 103664 301588 103670 301600
rect 130654 301588 130660 301600
rect 130712 301588 130718 301640
rect 107654 301520 107660 301572
rect 107712 301560 107718 301572
rect 139302 301560 139308 301572
rect 107712 301532 139308 301560
rect 107712 301520 107718 301532
rect 139302 301520 139308 301532
rect 139360 301560 139366 301572
rect 144270 301560 144276 301572
rect 139360 301532 144276 301560
rect 139360 301520 139366 301532
rect 144270 301520 144276 301532
rect 144328 301520 144334 301572
rect 129182 301452 129188 301504
rect 129240 301492 129246 301504
rect 162302 301492 162308 301504
rect 129240 301464 162308 301492
rect 129240 301452 129246 301464
rect 162302 301452 162308 301464
rect 162360 301452 162366 301504
rect 418798 301452 418804 301504
rect 418856 301492 418862 301504
rect 448514 301492 448520 301504
rect 418856 301464 448520 301492
rect 418856 301452 418862 301464
rect 448514 301452 448520 301464
rect 448572 301452 448578 301504
rect 74534 300976 74540 301028
rect 74592 301016 74598 301028
rect 149790 301016 149796 301028
rect 74592 300988 149796 301016
rect 74592 300976 74598 300988
rect 149790 300976 149796 300988
rect 149848 300976 149854 301028
rect 393590 300976 393596 301028
rect 393648 301016 393654 301028
rect 393958 301016 393964 301028
rect 393648 300988 393964 301016
rect 393648 300976 393654 300988
rect 393958 300976 393964 300988
rect 394016 301016 394022 301028
rect 446490 301016 446496 301028
rect 394016 300988 446496 301016
rect 394016 300976 394022 300988
rect 446490 300976 446496 300988
rect 446548 300976 446554 301028
rect 79226 300908 79232 300960
rect 79284 300948 79290 300960
rect 164970 300948 164976 300960
rect 79284 300920 164976 300948
rect 79284 300908 79290 300920
rect 164970 300908 164976 300920
rect 165028 300908 165034 300960
rect 376110 300908 376116 300960
rect 376168 300948 376174 300960
rect 409598 300948 409604 300960
rect 376168 300920 409604 300948
rect 376168 300908 376174 300920
rect 409598 300908 409604 300920
rect 409656 300908 409662 300960
rect 412358 300908 412364 300960
rect 412416 300948 412422 300960
rect 484394 300948 484400 300960
rect 412416 300920 484400 300948
rect 412416 300908 412422 300920
rect 484394 300908 484400 300920
rect 484452 300908 484458 300960
rect 59078 300840 59084 300892
rect 59136 300880 59142 300892
rect 59136 300852 155816 300880
rect 59136 300840 59142 300852
rect 155788 300824 155816 300852
rect 295334 300840 295340 300892
rect 295392 300880 295398 300892
rect 300302 300880 300308 300892
rect 295392 300852 300308 300880
rect 295392 300840 295398 300852
rect 300302 300840 300308 300852
rect 300360 300840 300366 300892
rect 301590 300840 301596 300892
rect 301648 300880 301654 300892
rect 436002 300880 436008 300892
rect 301648 300852 436008 300880
rect 301648 300840 301654 300852
rect 436002 300840 436008 300852
rect 436060 300840 436066 300892
rect 438486 300840 438492 300892
rect 438544 300880 438550 300892
rect 449894 300880 449900 300892
rect 438544 300852 449900 300880
rect 438544 300840 438550 300852
rect 449894 300840 449900 300852
rect 449952 300840 449958 300892
rect 155770 300772 155776 300824
rect 155828 300812 155834 300824
rect 159358 300812 159364 300824
rect 155828 300784 159364 300812
rect 155828 300772 155834 300784
rect 159358 300772 159364 300784
rect 159416 300772 159422 300824
rect 421006 300772 421012 300824
rect 421064 300812 421070 300824
rect 421834 300812 421840 300824
rect 421064 300784 421840 300812
rect 421064 300772 421070 300784
rect 421834 300772 421840 300784
rect 421892 300772 421898 300824
rect 116578 300228 116584 300280
rect 116636 300268 116642 300280
rect 129734 300268 129740 300280
rect 116636 300240 129740 300268
rect 116636 300228 116642 300240
rect 129734 300228 129740 300240
rect 129792 300228 129798 300280
rect 91094 300160 91100 300212
rect 91152 300200 91158 300212
rect 170674 300200 170680 300212
rect 91152 300172 170680 300200
rect 91152 300160 91158 300172
rect 170674 300160 170680 300172
rect 170732 300160 170738 300212
rect 39850 300092 39856 300144
rect 39908 300132 39914 300144
rect 127158 300132 127164 300144
rect 39908 300104 127164 300132
rect 39908 300092 39914 300104
rect 127158 300092 127164 300104
rect 127216 300092 127222 300144
rect 101490 299616 101496 299668
rect 101548 299656 101554 299668
rect 137278 299656 137284 299668
rect 101548 299628 137284 299656
rect 101548 299616 101554 299628
rect 137278 299616 137284 299628
rect 137336 299616 137342 299668
rect 416498 299616 416504 299668
rect 416556 299656 416562 299668
rect 438854 299656 438860 299668
rect 416556 299628 438860 299656
rect 416556 299616 416562 299628
rect 438854 299616 438860 299628
rect 438912 299616 438918 299668
rect 86954 299548 86960 299600
rect 87012 299588 87018 299600
rect 142798 299588 142804 299600
rect 87012 299560 142804 299588
rect 87012 299548 87018 299560
rect 142798 299548 142804 299560
rect 142856 299548 142862 299600
rect 358078 299548 358084 299600
rect 358136 299588 358142 299600
rect 414014 299588 414020 299600
rect 358136 299560 414020 299588
rect 358136 299548 358142 299560
rect 414014 299548 414020 299560
rect 414072 299548 414078 299600
rect 422018 299548 422024 299600
rect 422076 299588 422082 299600
rect 454126 299588 454132 299600
rect 422076 299560 454132 299588
rect 422076 299548 422082 299560
rect 454126 299548 454132 299560
rect 454184 299548 454190 299600
rect 67450 299480 67456 299532
rect 67508 299520 67514 299532
rect 152550 299520 152556 299532
rect 67508 299492 152556 299520
rect 67508 299480 67514 299492
rect 152550 299480 152556 299492
rect 152608 299480 152614 299532
rect 293218 299480 293224 299532
rect 293276 299520 293282 299532
rect 411806 299520 411812 299532
rect 293276 299492 411812 299520
rect 293276 299480 293282 299492
rect 411806 299480 411812 299492
rect 411864 299480 411870 299532
rect 414474 299480 414480 299532
rect 414532 299520 414538 299532
rect 476206 299520 476212 299532
rect 414532 299492 476212 299520
rect 414532 299480 414538 299492
rect 476206 299480 476212 299492
rect 476264 299480 476270 299532
rect 105538 299412 105544 299464
rect 105596 299452 105602 299464
rect 106090 299452 106096 299464
rect 105596 299424 106096 299452
rect 105596 299412 105602 299424
rect 106090 299412 106096 299424
rect 106148 299412 106154 299464
rect 167086 299412 167092 299464
rect 167144 299452 167150 299464
rect 168190 299452 168196 299464
rect 167144 299424 168196 299452
rect 167144 299412 167150 299424
rect 168190 299412 168196 299424
rect 168248 299452 168254 299464
rect 176654 299452 176660 299464
rect 168248 299424 176660 299452
rect 168248 299412 168254 299424
rect 176654 299412 176660 299424
rect 176712 299412 176718 299464
rect 438854 299412 438860 299464
rect 438912 299452 438918 299464
rect 553486 299452 553492 299464
rect 438912 299424 553492 299452
rect 438912 299412 438918 299424
rect 553486 299412 553492 299424
rect 553544 299452 553550 299464
rect 579614 299452 579620 299464
rect 553544 299424 579620 299452
rect 553544 299412 553550 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 108666 299344 108672 299396
rect 108724 299384 108730 299396
rect 111794 299384 111800 299396
rect 108724 299356 111800 299384
rect 108724 299344 108730 299356
rect 111794 299344 111800 299356
rect 111852 299344 111858 299396
rect 53558 298732 53564 298784
rect 53616 298772 53622 298784
rect 167086 298772 167092 298784
rect 53616 298744 167092 298772
rect 53616 298732 53622 298744
rect 167086 298732 167092 298744
rect 167144 298732 167150 298784
rect 112898 298392 112904 298444
rect 112956 298432 112962 298444
rect 149698 298432 149704 298444
rect 112956 298404 149704 298432
rect 112956 298392 112962 298404
rect 149698 298392 149704 298404
rect 149756 298392 149762 298444
rect 106090 298324 106096 298376
rect 106148 298364 106154 298376
rect 145650 298364 145656 298376
rect 106148 298336 145656 298364
rect 106148 298324 106154 298336
rect 145650 298324 145656 298336
rect 145708 298324 145714 298376
rect 84194 298256 84200 298308
rect 84252 298296 84258 298308
rect 141510 298296 141516 298308
rect 84252 298268 141516 298296
rect 84252 298256 84258 298268
rect 141510 298256 141516 298268
rect 141568 298256 141574 298308
rect 68462 298188 68468 298240
rect 68520 298228 68526 298240
rect 160830 298228 160836 298240
rect 68520 298200 160836 298228
rect 68520 298188 68526 298200
rect 160830 298188 160836 298200
rect 160888 298188 160894 298240
rect 72970 298120 72976 298172
rect 73028 298160 73034 298172
rect 170582 298160 170588 298172
rect 73028 298132 170588 298160
rect 73028 298120 73034 298132
rect 170582 298120 170588 298132
rect 170640 298120 170646 298172
rect 52454 298052 52460 298104
rect 52512 298092 52518 298104
rect 53650 298092 53656 298104
rect 52512 298064 53656 298092
rect 52512 298052 52518 298064
rect 53650 298052 53656 298064
rect 53708 298092 53714 298104
rect 101398 298092 101404 298104
rect 53708 298064 101404 298092
rect 53708 298052 53714 298064
rect 101398 298052 101404 298064
rect 101456 298052 101462 298104
rect 44818 297372 44824 297424
rect 44876 297412 44882 297424
rect 52454 297412 52460 297424
rect 44876 297384 52460 297412
rect 44876 297372 44882 297384
rect 52454 297372 52460 297384
rect 52512 297372 52518 297424
rect 314010 297372 314016 297424
rect 314068 297412 314074 297424
rect 369762 297412 369768 297424
rect 314068 297384 369768 297412
rect 314068 297372 314074 297384
rect 369762 297372 369768 297384
rect 369820 297372 369826 297424
rect 102870 297032 102876 297084
rect 102928 297072 102934 297084
rect 134518 297072 134524 297084
rect 102928 297044 134524 297072
rect 102928 297032 102934 297044
rect 134518 297032 134524 297044
rect 134576 297032 134582 297084
rect 93210 296964 93216 297016
rect 93268 297004 93274 297016
rect 124858 297004 124864 297016
rect 93268 296976 124864 297004
rect 93268 296964 93274 296976
rect 124858 296964 124864 296976
rect 124916 296964 124922 297016
rect 83550 296896 83556 296948
rect 83608 296936 83614 296948
rect 144362 296936 144368 296948
rect 83608 296908 144368 296936
rect 83608 296896 83614 296908
rect 144362 296896 144368 296908
rect 144420 296896 144426 296948
rect 172330 296896 172336 296948
rect 172388 296936 172394 296948
rect 176654 296936 176660 296948
rect 172388 296908 176660 296936
rect 172388 296896 172394 296908
rect 176654 296896 176660 296908
rect 176712 296896 176718 296948
rect 442810 296896 442816 296948
rect 442868 296936 442874 296948
rect 444558 296936 444564 296948
rect 442868 296908 444564 296936
rect 442868 296896 442874 296908
rect 444558 296896 444564 296908
rect 444616 296896 444622 296948
rect 93854 296828 93860 296880
rect 93912 296868 93918 296880
rect 159358 296868 159364 296880
rect 93912 296840 159364 296868
rect 93912 296828 93918 296840
rect 159358 296828 159364 296840
rect 159416 296828 159422 296880
rect 95142 296760 95148 296812
rect 95200 296800 95206 296812
rect 102778 296800 102784 296812
rect 95200 296772 102784 296800
rect 95200 296760 95206 296772
rect 102778 296760 102784 296772
rect 102836 296800 102842 296812
rect 172330 296800 172336 296812
rect 102836 296772 172336 296800
rect 102836 296760 102842 296772
rect 172330 296760 172336 296772
rect 172388 296760 172394 296812
rect 50706 296692 50712 296744
rect 50764 296732 50770 296744
rect 158162 296732 158168 296744
rect 50764 296704 158168 296732
rect 50764 296692 50770 296704
rect 158162 296692 158168 296704
rect 158220 296692 158226 296744
rect 369762 296692 369768 296744
rect 369820 296732 369826 296744
rect 376938 296732 376944 296744
rect 369820 296704 376944 296732
rect 369820 296692 369826 296704
rect 376938 296692 376944 296704
rect 376996 296692 377002 296744
rect 60458 296012 60464 296064
rect 60516 296052 60522 296064
rect 84838 296052 84844 296064
rect 60516 296024 84844 296052
rect 60516 296012 60522 296024
rect 84838 296012 84844 296024
rect 84896 296012 84902 296064
rect 67358 295944 67364 295996
rect 67416 295984 67422 295996
rect 169110 295984 169116 295996
rect 67416 295956 169116 295984
rect 67416 295944 67422 295956
rect 169110 295944 169116 295956
rect 169168 295944 169174 295996
rect 113818 295604 113824 295656
rect 113876 295644 113882 295656
rect 123570 295644 123576 295656
rect 113876 295616 123576 295644
rect 113876 295604 113882 295616
rect 123570 295604 123576 295616
rect 123628 295604 123634 295656
rect 118510 295536 118516 295588
rect 118568 295576 118574 295588
rect 119614 295576 119620 295588
rect 118568 295548 119620 295576
rect 118568 295536 118574 295548
rect 119614 295536 119620 295548
rect 119672 295536 119678 295588
rect 82906 295468 82912 295520
rect 82964 295508 82970 295520
rect 134702 295508 134708 295520
rect 82964 295480 134708 295508
rect 82964 295468 82970 295480
rect 134702 295468 134708 295480
rect 134760 295468 134766 295520
rect 100938 295400 100944 295452
rect 100996 295440 101002 295452
rect 155218 295440 155224 295452
rect 100996 295412 155224 295440
rect 100996 295400 101002 295412
rect 155218 295400 155224 295412
rect 155276 295400 155282 295452
rect 69014 295332 69020 295384
rect 69072 295372 69078 295384
rect 71774 295372 71780 295384
rect 69072 295344 71780 295372
rect 69072 295332 69078 295344
rect 71774 295332 71780 295344
rect 71832 295332 71838 295384
rect 94498 295332 94504 295384
rect 94556 295372 94562 295384
rect 95050 295372 95056 295384
rect 94556 295344 95056 295372
rect 94556 295332 94562 295344
rect 95050 295332 95056 295344
rect 95108 295372 95114 295384
rect 148502 295372 148508 295384
rect 95108 295344 148508 295372
rect 95108 295332 95114 295344
rect 148502 295332 148508 295344
rect 148560 295332 148566 295384
rect 295334 295332 295340 295384
rect 295392 295372 295398 295384
rect 309870 295372 309876 295384
rect 295392 295344 309876 295372
rect 295392 295332 295398 295344
rect 309870 295332 309876 295344
rect 309928 295372 309934 295384
rect 310330 295372 310336 295384
rect 309928 295344 310336 295372
rect 309928 295332 309934 295344
rect 310330 295332 310336 295344
rect 310388 295332 310394 295384
rect 46566 295264 46572 295316
rect 46624 295304 46630 295316
rect 72970 295304 72976 295316
rect 46624 295276 72976 295304
rect 46624 295264 46630 295276
rect 72970 295264 72976 295276
rect 73028 295304 73034 295316
rect 73890 295304 73896 295316
rect 73028 295276 73896 295304
rect 73028 295264 73034 295276
rect 73890 295264 73896 295276
rect 73948 295264 73954 295316
rect 297634 295264 297640 295316
rect 297692 295304 297698 295316
rect 379146 295304 379152 295316
rect 297692 295276 379152 295304
rect 297692 295264 297698 295276
rect 379146 295264 379152 295276
rect 379204 295264 379210 295316
rect 310330 295196 310336 295248
rect 310388 295236 310394 295248
rect 319438 295236 319444 295248
rect 310388 295208 319444 295236
rect 310388 295196 310394 295208
rect 319438 295196 319444 295208
rect 319496 295196 319502 295248
rect 73246 294924 73252 294976
rect 73304 294964 73310 294976
rect 74626 294964 74632 294976
rect 73304 294936 74632 294964
rect 73304 294924 73310 294936
rect 74626 294924 74632 294936
rect 74684 294924 74690 294976
rect 73798 294788 73804 294840
rect 73856 294828 73862 294840
rect 84838 294828 84844 294840
rect 73856 294800 84844 294828
rect 73856 294788 73862 294800
rect 84838 294788 84844 294800
rect 84896 294788 84902 294840
rect 70026 294652 70032 294704
rect 70084 294692 70090 294704
rect 101490 294692 101496 294704
rect 70084 294664 101496 294692
rect 70084 294652 70090 294664
rect 101490 294652 101496 294664
rect 101548 294652 101554 294704
rect 9582 294584 9588 294636
rect 9640 294624 9646 294636
rect 72602 294624 72608 294636
rect 9640 294596 72608 294624
rect 9640 294584 9646 294596
rect 72602 294584 72608 294596
rect 72660 294584 72666 294636
rect 95786 294584 95792 294636
rect 95844 294624 95850 294636
rect 168282 294624 168288 294636
rect 95844 294596 168288 294624
rect 95844 294584 95850 294596
rect 168282 294584 168288 294596
rect 168340 294584 168346 294636
rect 442810 294584 442816 294636
rect 442868 294624 442874 294636
rect 452746 294624 452752 294636
rect 442868 294596 452752 294624
rect 442868 294584 442874 294596
rect 452746 294584 452752 294596
rect 452804 294584 452810 294636
rect 75178 294244 75184 294296
rect 75236 294284 75242 294296
rect 141418 294284 141424 294296
rect 75236 294256 141424 294284
rect 75236 294244 75242 294256
rect 141418 294244 141424 294256
rect 141476 294244 141482 294296
rect 85482 294176 85488 294228
rect 85540 294216 85546 294228
rect 91738 294216 91744 294228
rect 85540 294188 91744 294216
rect 85540 294176 85546 294188
rect 91738 294176 91744 294188
rect 91796 294176 91802 294228
rect 91922 294176 91928 294228
rect 91980 294216 91986 294228
rect 133138 294216 133144 294228
rect 91980 294188 133144 294216
rect 91980 294176 91986 294188
rect 133138 294176 133144 294188
rect 133196 294176 133202 294228
rect 62758 294108 62764 294160
rect 62816 294148 62822 294160
rect 96614 294148 96620 294160
rect 62816 294120 96620 294148
rect 62816 294108 62822 294120
rect 96614 294108 96620 294120
rect 96672 294108 96678 294160
rect 102226 294108 102232 294160
rect 102284 294148 102290 294160
rect 151170 294148 151176 294160
rect 102284 294120 151176 294148
rect 102284 294108 102290 294120
rect 151170 294108 151176 294120
rect 151228 294108 151234 294160
rect 78398 294040 78404 294092
rect 78456 294080 78462 294092
rect 129090 294080 129096 294092
rect 78456 294052 129096 294080
rect 78456 294040 78462 294052
rect 129090 294040 129096 294052
rect 129148 294040 129154 294092
rect 70394 293972 70400 294024
rect 70452 294012 70458 294024
rect 71038 294012 71044 294024
rect 70452 293984 71044 294012
rect 70452 293972 70458 293984
rect 71038 293972 71044 293984
rect 71096 293972 71102 294024
rect 76466 293972 76472 294024
rect 76524 294012 76530 294024
rect 77938 294012 77944 294024
rect 76524 293984 77944 294012
rect 76524 293972 76530 293984
rect 77938 293972 77944 293984
rect 77996 293972 78002 294024
rect 81434 293972 81440 294024
rect 81492 294012 81498 294024
rect 81894 294012 81900 294024
rect 81492 293984 81900 294012
rect 81492 293972 81498 293984
rect 81894 293972 81900 293984
rect 81952 293972 81958 294024
rect 88334 293972 88340 294024
rect 88392 294012 88398 294024
rect 89070 294012 89076 294024
rect 88392 293984 89076 294012
rect 88392 293972 88398 293984
rect 89070 293972 89076 293984
rect 89128 293972 89134 294024
rect 103606 293972 103612 294024
rect 103664 294012 103670 294024
rect 104526 294012 104532 294024
rect 103664 293984 104532 294012
rect 103664 293972 103670 293984
rect 104526 293972 104532 293984
rect 104584 293972 104590 294024
rect 109034 293972 109040 294024
rect 109092 294012 109098 294024
rect 109678 294012 109684 294024
rect 109092 293984 109684 294012
rect 109092 293972 109098 293984
rect 109678 293972 109684 293984
rect 109736 293972 109742 294024
rect 111886 293972 111892 294024
rect 111944 294012 111950 294024
rect 111944 293984 114508 294012
rect 111944 293972 111950 293984
rect 114480 293944 114508 293984
rect 114554 293972 114560 294024
rect 114612 294012 114618 294024
rect 115382 294012 115388 294024
rect 114612 293984 115388 294012
rect 114612 293972 114618 293984
rect 115382 293972 115388 293984
rect 115440 293972 115446 294024
rect 120350 294012 120356 294024
rect 115492 293984 120356 294012
rect 115492 293944 115520 293984
rect 120350 293972 120356 293984
rect 120408 293972 120414 294024
rect 173342 293972 173348 294024
rect 173400 294012 173406 294024
rect 176654 294012 176660 294024
rect 173400 293984 176660 294012
rect 173400 293972 173406 293984
rect 176654 293972 176660 293984
rect 176712 293972 176718 294024
rect 114480 293916 115520 293944
rect 79042 293496 79048 293548
rect 79100 293536 79106 293548
rect 79318 293536 79324 293548
rect 79100 293508 79324 293536
rect 79100 293496 79106 293508
rect 79318 293496 79324 293508
rect 79376 293496 79382 293548
rect 98362 293496 98368 293548
rect 98420 293536 98426 293548
rect 98638 293536 98644 293548
rect 98420 293508 98644 293536
rect 98420 293496 98426 293508
rect 98638 293496 98644 293508
rect 98696 293496 98702 293548
rect 296714 293224 296720 293276
rect 296772 293264 296778 293276
rect 307018 293264 307024 293276
rect 296772 293236 307024 293264
rect 296772 293224 296778 293236
rect 307018 293224 307024 293236
rect 307076 293224 307082 293276
rect 116394 292884 116400 292936
rect 116452 292924 116458 292936
rect 116762 292924 116768 292936
rect 116452 292896 116768 292924
rect 116452 292884 116458 292896
rect 116762 292884 116768 292896
rect 116820 292924 116826 292936
rect 123662 292924 123668 292936
rect 116820 292896 123668 292924
rect 116820 292884 116826 292896
rect 123662 292884 123668 292896
rect 123720 292884 123726 292936
rect 99650 292816 99656 292868
rect 99708 292856 99714 292868
rect 131758 292856 131764 292868
rect 99708 292828 131764 292856
rect 99708 292816 99714 292828
rect 131758 292816 131764 292828
rect 131816 292816 131822 292868
rect 58710 292748 58716 292800
rect 58768 292788 58774 292800
rect 92566 292788 92572 292800
rect 58768 292760 92572 292788
rect 58768 292748 58774 292760
rect 92566 292748 92572 292760
rect 92624 292748 92630 292800
rect 105446 292748 105452 292800
rect 105504 292788 105510 292800
rect 106182 292788 106188 292800
rect 105504 292760 106188 292788
rect 105504 292748 105510 292760
rect 106182 292748 106188 292760
rect 106240 292788 106246 292800
rect 152642 292788 152648 292800
rect 106240 292760 152648 292788
rect 106240 292748 106246 292760
rect 152642 292748 152648 292760
rect 152700 292748 152706 292800
rect 88058 292680 88064 292732
rect 88116 292720 88122 292732
rect 136174 292720 136180 292732
rect 88116 292692 136180 292720
rect 88116 292680 88122 292692
rect 136174 292680 136180 292692
rect 136232 292680 136238 292732
rect 57238 292612 57244 292664
rect 57296 292652 57302 292664
rect 79042 292652 79048 292664
rect 57296 292624 79048 292652
rect 57296 292612 57302 292624
rect 79042 292612 79048 292624
rect 79100 292612 79106 292664
rect 80974 292612 80980 292664
rect 81032 292652 81038 292664
rect 138750 292652 138756 292664
rect 81032 292624 138756 292652
rect 81032 292612 81038 292624
rect 138750 292612 138756 292624
rect 138808 292612 138814 292664
rect 4062 292544 4068 292596
rect 4120 292584 4126 292596
rect 95970 292584 95976 292596
rect 4120 292556 95976 292584
rect 4120 292544 4126 292556
rect 95970 292544 95976 292556
rect 96028 292544 96034 292596
rect 98362 292544 98368 292596
rect 98420 292584 98426 292596
rect 178678 292584 178684 292596
rect 98420 292556 178684 292584
rect 98420 292544 98426 292556
rect 178678 292544 178684 292556
rect 178736 292544 178742 292596
rect 295334 292476 295340 292528
rect 295392 292516 295398 292528
rect 305086 292516 305092 292528
rect 295392 292488 305092 292516
rect 295392 292476 295398 292488
rect 305086 292476 305092 292488
rect 305144 292516 305150 292528
rect 305546 292516 305552 292528
rect 305144 292488 305552 292516
rect 305144 292476 305150 292488
rect 305546 292476 305552 292488
rect 305604 292476 305610 292528
rect 86402 291864 86408 291916
rect 86460 291904 86466 291916
rect 86460 291876 93854 291904
rect 86460 291864 86466 291876
rect 3234 291796 3240 291848
rect 3292 291836 3298 291848
rect 17218 291836 17224 291848
rect 3292 291808 17224 291836
rect 3292 291796 3298 291808
rect 17218 291796 17224 291808
rect 17276 291796 17282 291848
rect 68462 291796 68468 291848
rect 68520 291836 68526 291848
rect 68646 291836 68652 291848
rect 68520 291808 68652 291836
rect 68520 291796 68526 291808
rect 68646 291796 68652 291808
rect 68704 291796 68710 291848
rect 93826 291224 93854 291876
rect 110782 291864 110788 291916
rect 110840 291864 110846 291916
rect 122558 291864 122564 291916
rect 122616 291904 122622 291916
rect 122742 291904 122748 291916
rect 122616 291876 122748 291904
rect 122616 291864 122622 291876
rect 122742 291864 122748 291876
rect 122800 291864 122806 291916
rect 110800 291292 110828 291864
rect 120350 291796 120356 291848
rect 120408 291836 120414 291848
rect 141602 291836 141608 291848
rect 120408 291808 141608 291836
rect 120408 291796 120414 291808
rect 141602 291796 141608 291808
rect 141660 291796 141666 291848
rect 151354 291292 151360 291304
rect 110800 291264 151360 291292
rect 151354 291252 151360 291264
rect 151412 291252 151418 291304
rect 147030 291224 147036 291236
rect 93826 291196 147036 291224
rect 147030 291184 147036 291196
rect 147088 291184 147094 291236
rect 163682 291116 163688 291168
rect 163740 291156 163746 291168
rect 164142 291156 164148 291168
rect 163740 291128 164148 291156
rect 163740 291116 163746 291128
rect 164142 291116 164148 291128
rect 164200 291116 164206 291168
rect 294046 291116 294052 291168
rect 294104 291156 294110 291168
rect 343726 291156 343732 291168
rect 294104 291128 343732 291156
rect 294104 291116 294110 291128
rect 343726 291116 343732 291128
rect 343784 291116 343790 291168
rect 13078 290436 13084 290488
rect 13136 290476 13142 290488
rect 39942 290476 39948 290488
rect 13136 290448 39948 290476
rect 13136 290436 13142 290448
rect 39942 290436 39948 290448
rect 40000 290476 40006 290488
rect 49602 290476 49608 290488
rect 40000 290448 49608 290476
rect 40000 290436 40006 290448
rect 49602 290436 49608 290448
rect 49660 290436 49666 290488
rect 126330 290436 126336 290488
rect 126388 290476 126394 290488
rect 148318 290476 148324 290488
rect 126388 290448 148324 290476
rect 126388 290436 126394 290448
rect 148318 290436 148324 290448
rect 148376 290436 148382 290488
rect 163682 290436 163688 290488
rect 163740 290476 163746 290488
rect 176654 290476 176660 290488
rect 163740 290448 176660 290476
rect 163740 290436 163746 290448
rect 176654 290436 176660 290448
rect 176712 290436 176718 290488
rect 343726 290436 343732 290488
rect 343784 290476 343790 290488
rect 365162 290476 365168 290488
rect 343784 290448 365168 290476
rect 343784 290436 343790 290448
rect 365162 290436 365168 290448
rect 365220 290436 365226 290488
rect 373258 290436 373264 290488
rect 373316 290476 373322 290488
rect 373810 290476 373816 290488
rect 373316 290448 373816 290476
rect 373316 290436 373322 290448
rect 373810 290436 373816 290448
rect 373868 290476 373874 290488
rect 376938 290476 376944 290488
rect 373868 290448 376944 290476
rect 373868 290436 373874 290448
rect 376938 290436 376944 290448
rect 376996 290436 377002 290488
rect 49602 289892 49608 289944
rect 49660 289932 49666 289944
rect 67726 289932 67732 289944
rect 49660 289904 67732 289932
rect 49660 289892 49666 289904
rect 67726 289892 67732 289904
rect 67784 289892 67790 289944
rect 121546 289892 121552 289944
rect 121604 289932 121610 289944
rect 140130 289932 140136 289944
rect 121604 289904 140136 289932
rect 121604 289892 121610 289904
rect 140130 289892 140136 289904
rect 140188 289892 140194 289944
rect 43806 289824 43812 289876
rect 43864 289864 43870 289876
rect 67634 289864 67640 289876
rect 43864 289836 67640 289864
rect 43864 289824 43870 289836
rect 67634 289824 67640 289836
rect 67692 289824 67698 289876
rect 121638 289824 121644 289876
rect 121696 289864 121702 289876
rect 167638 289864 167644 289876
rect 121696 289836 167644 289864
rect 121696 289824 121702 289836
rect 167638 289824 167644 289836
rect 167696 289824 167702 289876
rect 295334 289824 295340 289876
rect 295392 289864 295398 289876
rect 295392 289836 306374 289864
rect 295392 289824 295398 289836
rect 306346 289808 306374 289836
rect 440326 289824 440332 289876
rect 440384 289864 440390 289876
rect 449986 289864 449992 289876
rect 440384 289836 449992 289864
rect 440384 289824 440390 289836
rect 449986 289824 449992 289836
rect 450044 289824 450050 289876
rect 121546 289756 121552 289808
rect 121604 289796 121610 289808
rect 145558 289796 145564 289808
rect 121604 289768 145564 289796
rect 121604 289756 121610 289768
rect 145558 289756 145564 289768
rect 145616 289756 145622 289808
rect 306282 289756 306288 289808
rect 306340 289796 306374 289808
rect 307754 289796 307760 289808
rect 306340 289768 307760 289796
rect 306340 289756 306346 289768
rect 307754 289756 307760 289768
rect 307812 289756 307818 289808
rect 377950 289756 377956 289808
rect 378008 289796 378014 289808
rect 378778 289796 378784 289808
rect 378008 289768 378784 289796
rect 378008 289756 378014 289768
rect 378778 289756 378784 289768
rect 378836 289756 378842 289808
rect 121638 289688 121644 289740
rect 121696 289728 121702 289740
rect 133874 289728 133880 289740
rect 121696 289700 133880 289728
rect 121696 289688 121702 289700
rect 133874 289688 133880 289700
rect 133932 289728 133938 289740
rect 135162 289728 135168 289740
rect 133932 289700 135168 289728
rect 133932 289688 133938 289700
rect 135162 289688 135168 289700
rect 135220 289688 135226 289740
rect 300302 289688 300308 289740
rect 300360 289728 300366 289740
rect 311894 289728 311900 289740
rect 300360 289700 311900 289728
rect 300360 289688 300366 289700
rect 311894 289688 311900 289700
rect 311952 289688 311958 289740
rect 43898 289076 43904 289128
rect 43956 289116 43962 289128
rect 64874 289116 64880 289128
rect 43956 289088 64880 289116
rect 43956 289076 43962 289088
rect 64874 289076 64880 289088
rect 64932 289116 64938 289128
rect 67726 289116 67732 289128
rect 64932 289088 67732 289116
rect 64932 289076 64938 289088
rect 67726 289076 67732 289088
rect 67784 289076 67790 289128
rect 311894 289076 311900 289128
rect 311952 289116 311958 289128
rect 312538 289116 312544 289128
rect 311952 289088 312544 289116
rect 311952 289076 311958 289088
rect 312538 289076 312544 289088
rect 312596 289116 312602 289128
rect 367002 289116 367008 289128
rect 312596 289088 367008 289116
rect 312596 289076 312602 289088
rect 367002 289076 367008 289088
rect 367060 289076 367066 289128
rect 64598 288396 64604 288448
rect 64656 288436 64662 288448
rect 67634 288436 67640 288448
rect 64656 288408 67640 288436
rect 64656 288396 64662 288408
rect 67634 288396 67640 288408
rect 67692 288396 67698 288448
rect 367002 288396 367008 288448
rect 367060 288436 367066 288448
rect 376938 288436 376944 288448
rect 367060 288408 376944 288436
rect 367060 288396 367066 288408
rect 376938 288396 376944 288408
rect 376996 288396 377002 288448
rect 121546 288328 121552 288380
rect 121604 288368 121610 288380
rect 174538 288368 174544 288380
rect 121604 288340 174544 288368
rect 121604 288328 121610 288340
rect 174538 288328 174544 288340
rect 174596 288328 174602 288380
rect 170582 288260 170588 288312
rect 170640 288300 170646 288312
rect 176654 288300 176660 288312
rect 170640 288272 176660 288300
rect 170640 288260 170646 288272
rect 176654 288260 176660 288272
rect 176712 288260 176718 288312
rect 48038 287036 48044 287088
rect 48096 287076 48102 287088
rect 67634 287076 67640 287088
rect 48096 287048 67640 287076
rect 48096 287036 48102 287048
rect 67634 287036 67640 287048
rect 67692 287036 67698 287088
rect 296162 287036 296168 287088
rect 296220 287076 296226 287088
rect 342898 287076 342904 287088
rect 296220 287048 342904 287076
rect 296220 287036 296226 287048
rect 342898 287036 342904 287048
rect 342956 287036 342962 287088
rect 441522 287036 441528 287088
rect 441580 287076 441586 287088
rect 447778 287076 447784 287088
rect 441580 287048 447784 287076
rect 441580 287036 441586 287048
rect 447778 287036 447784 287048
rect 447836 287036 447842 287088
rect 138842 286356 138848 286408
rect 138900 286396 138906 286408
rect 142154 286396 142160 286408
rect 138900 286368 142160 286396
rect 138900 286356 138906 286368
rect 142154 286356 142160 286368
rect 142212 286396 142218 286408
rect 157150 286396 157156 286408
rect 142212 286368 157156 286396
rect 142212 286356 142218 286368
rect 157150 286356 157156 286368
rect 157208 286396 157214 286408
rect 173342 286396 173348 286408
rect 157208 286368 173348 286396
rect 157208 286356 157214 286368
rect 173342 286356 173348 286368
rect 173400 286356 173406 286408
rect 121730 286288 121736 286340
rect 121788 286328 121794 286340
rect 124306 286328 124312 286340
rect 121788 286300 124312 286328
rect 121788 286288 121794 286300
rect 124306 286288 124312 286300
rect 124364 286328 124370 286340
rect 163590 286328 163596 286340
rect 124364 286300 163596 286328
rect 124364 286288 124370 286300
rect 163590 286288 163596 286300
rect 163648 286288 163654 286340
rect 325234 286288 325240 286340
rect 325292 286328 325298 286340
rect 369854 286328 369860 286340
rect 325292 286300 369860 286328
rect 325292 286288 325298 286300
rect 369854 286288 369860 286300
rect 369912 286288 369918 286340
rect 50982 285676 50988 285728
rect 51040 285716 51046 285728
rect 67726 285716 67732 285728
rect 51040 285688 67732 285716
rect 51040 285676 51046 285688
rect 67726 285676 67732 285688
rect 67784 285676 67790 285728
rect 369854 285676 369860 285728
rect 369912 285716 369918 285728
rect 371142 285716 371148 285728
rect 369912 285688 371148 285716
rect 369912 285676 369918 285688
rect 371142 285676 371148 285688
rect 371200 285716 371206 285728
rect 376938 285716 376944 285728
rect 371200 285688 376944 285716
rect 371200 285676 371206 285688
rect 376938 285676 376944 285688
rect 376996 285676 377002 285728
rect 445018 285676 445024 285728
rect 445076 285716 445082 285728
rect 480346 285716 480352 285728
rect 445076 285688 480352 285716
rect 445076 285676 445082 285688
rect 480346 285676 480352 285688
rect 480404 285676 480410 285728
rect 121454 285608 121460 285660
rect 121512 285648 121518 285660
rect 125594 285648 125600 285660
rect 121512 285620 125600 285648
rect 121512 285608 121518 285620
rect 125594 285608 125600 285620
rect 125652 285608 125658 285660
rect 442166 285608 442172 285660
rect 442224 285648 442230 285660
rect 445036 285648 445064 285676
rect 442224 285620 445064 285648
rect 442224 285608 442230 285620
rect 122466 284928 122472 284980
rect 122524 284968 122530 284980
rect 169110 284968 169116 284980
rect 122524 284940 169116 284968
rect 122524 284928 122530 284940
rect 169110 284928 169116 284940
rect 169168 284928 169174 284980
rect 41230 284316 41236 284368
rect 41288 284356 41294 284368
rect 67634 284356 67640 284368
rect 41288 284328 67640 284356
rect 41288 284316 41294 284328
rect 67634 284316 67640 284328
rect 67692 284316 67698 284368
rect 160830 284316 160836 284368
rect 160888 284356 160894 284368
rect 162762 284356 162768 284368
rect 160888 284328 162768 284356
rect 160888 284316 160894 284328
rect 162762 284316 162768 284328
rect 162820 284356 162826 284368
rect 174630 284356 174636 284368
rect 162820 284328 174636 284356
rect 162820 284316 162826 284328
rect 174630 284316 174636 284328
rect 174688 284316 174694 284368
rect 50706 284248 50712 284300
rect 50764 284288 50770 284300
rect 67726 284288 67732 284300
rect 50764 284260 67732 284288
rect 50764 284248 50770 284260
rect 67726 284248 67732 284260
rect 67784 284248 67790 284300
rect 122742 284248 122748 284300
rect 122800 284288 122806 284300
rect 124214 284288 124220 284300
rect 122800 284260 124220 284288
rect 122800 284248 122806 284260
rect 124214 284248 124220 284260
rect 124272 284248 124278 284300
rect 158622 284248 158628 284300
rect 158680 284288 158686 284300
rect 176654 284288 176660 284300
rect 158680 284260 176660 284288
rect 158680 284248 158686 284260
rect 176654 284248 176660 284260
rect 176712 284248 176718 284300
rect 121454 283568 121460 283620
rect 121512 283608 121518 283620
rect 173158 283608 173164 283620
rect 121512 283580 173164 283608
rect 121512 283568 121518 283580
rect 173158 283568 173164 283580
rect 173216 283608 173222 283620
rect 173342 283608 173348 283620
rect 173216 283580 173348 283608
rect 173216 283568 173222 283580
rect 173342 283568 173348 283580
rect 173400 283568 173406 283620
rect 298738 283568 298744 283620
rect 298796 283608 298802 283620
rect 377306 283608 377312 283620
rect 298796 283580 377312 283608
rect 298796 283568 298802 283580
rect 377306 283568 377312 283580
rect 377364 283608 377370 283620
rect 377858 283608 377864 283620
rect 377364 283580 377864 283608
rect 377364 283568 377370 283580
rect 377858 283568 377864 283580
rect 377916 283568 377922 283620
rect 294782 282888 294788 282940
rect 294840 282928 294846 282940
rect 310514 282928 310520 282940
rect 294840 282900 310520 282928
rect 294840 282888 294846 282900
rect 310514 282888 310520 282900
rect 310572 282928 310578 282940
rect 376018 282928 376024 282940
rect 310572 282900 376024 282928
rect 310572 282888 310578 282900
rect 376018 282888 376024 282900
rect 376076 282888 376082 282940
rect 166258 282820 166264 282872
rect 166316 282860 166322 282872
rect 176654 282860 176660 282872
rect 166316 282832 176660 282860
rect 166316 282820 166322 282832
rect 176654 282820 176660 282832
rect 176712 282820 176718 282872
rect 442718 281800 442724 281852
rect 442776 281840 442782 281852
rect 450078 281840 450084 281852
rect 442776 281812 450084 281840
rect 442776 281800 442782 281812
rect 450078 281800 450084 281812
rect 450136 281800 450142 281852
rect 121546 281596 121552 281648
rect 121604 281636 121610 281648
rect 148318 281636 148324 281648
rect 121604 281608 148324 281636
rect 121604 281596 121610 281608
rect 148318 281596 148324 281608
rect 148376 281596 148382 281648
rect 311710 281596 311716 281648
rect 311768 281636 311774 281648
rect 313366 281636 313372 281648
rect 311768 281608 313372 281636
rect 311768 281596 311774 281608
rect 313366 281596 313372 281608
rect 313424 281636 313430 281648
rect 354582 281636 354588 281648
rect 313424 281608 354588 281636
rect 313424 281596 313430 281608
rect 354582 281596 354588 281608
rect 354640 281636 354646 281648
rect 354640 281596 354674 281636
rect 121454 281528 121460 281580
rect 121512 281568 121518 281580
rect 158070 281568 158076 281580
rect 121512 281540 158076 281568
rect 121512 281528 121518 281540
rect 158070 281528 158076 281540
rect 158128 281528 158134 281580
rect 295334 281528 295340 281580
rect 295392 281568 295398 281580
rect 298278 281568 298284 281580
rect 295392 281540 298284 281568
rect 295392 281528 295398 281540
rect 298278 281528 298284 281540
rect 298336 281568 298342 281580
rect 349890 281568 349896 281580
rect 298336 281540 349896 281568
rect 298336 281528 298342 281540
rect 349890 281528 349896 281540
rect 349948 281528 349954 281580
rect 354646 281568 354674 281596
rect 376938 281568 376944 281580
rect 354646 281540 376944 281568
rect 376938 281528 376944 281540
rect 376996 281528 377002 281580
rect 360010 280848 360016 280900
rect 360068 280888 360074 280900
rect 371234 280888 371240 280900
rect 360068 280860 371240 280888
rect 360068 280848 360074 280860
rect 371234 280848 371240 280860
rect 371292 280848 371298 280900
rect 56318 280780 56324 280832
rect 56376 280820 56382 280832
rect 67634 280820 67640 280832
rect 56376 280792 67640 280820
rect 56376 280780 56382 280792
rect 67634 280780 67640 280792
rect 67692 280780 67698 280832
rect 125134 280780 125140 280832
rect 125192 280820 125198 280832
rect 163682 280820 163688 280832
rect 125192 280792 163688 280820
rect 125192 280780 125198 280792
rect 163682 280780 163688 280792
rect 163740 280780 163746 280832
rect 300302 280780 300308 280832
rect 300360 280820 300366 280832
rect 376202 280820 376208 280832
rect 300360 280792 376208 280820
rect 300360 280780 300366 280792
rect 376202 280780 376208 280792
rect 376260 280780 376266 280832
rect 476114 280780 476120 280832
rect 476172 280820 476178 280832
rect 496078 280820 496084 280832
rect 476172 280792 496084 280820
rect 476172 280780 476178 280792
rect 496078 280780 496084 280792
rect 496136 280780 496142 280832
rect 52178 280168 52184 280220
rect 52236 280208 52242 280220
rect 67634 280208 67640 280220
rect 52236 280180 67640 280208
rect 52236 280168 52242 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121454 280168 121460 280220
rect 121512 280208 121518 280220
rect 134794 280208 134800 280220
rect 121512 280180 134800 280208
rect 121512 280168 121518 280180
rect 134794 280168 134800 280180
rect 134852 280168 134858 280220
rect 371234 280168 371240 280220
rect 371292 280208 371298 280220
rect 372522 280208 372528 280220
rect 371292 280180 372528 280208
rect 371292 280168 371298 280180
rect 372522 280168 372528 280180
rect 372580 280208 372586 280220
rect 376938 280208 376944 280220
rect 372580 280180 376944 280208
rect 372580 280168 372586 280180
rect 376938 280168 376944 280180
rect 376996 280168 377002 280220
rect 442810 280168 442816 280220
rect 442868 280208 442874 280220
rect 476114 280208 476120 280220
rect 442868 280180 476120 280208
rect 442868 280168 442874 280180
rect 476114 280168 476120 280180
rect 476172 280168 476178 280220
rect 174630 280100 174636 280152
rect 174688 280140 174694 280152
rect 176654 280140 176660 280152
rect 174688 280112 176660 280140
rect 174688 280100 174694 280112
rect 176654 280100 176660 280112
rect 176712 280100 176718 280152
rect 31018 279420 31024 279472
rect 31076 279460 31082 279472
rect 67450 279460 67456 279472
rect 31076 279432 67456 279460
rect 31076 279420 31082 279432
rect 67450 279420 67456 279432
rect 67508 279460 67514 279472
rect 67634 279460 67640 279472
rect 67508 279432 67640 279460
rect 67508 279420 67514 279432
rect 67634 279420 67640 279432
rect 67692 279420 67698 279472
rect 122650 279420 122656 279472
rect 122708 279460 122714 279472
rect 160830 279460 160836 279472
rect 122708 279432 160836 279460
rect 122708 279420 122714 279432
rect 160830 279420 160836 279432
rect 160888 279420 160894 279472
rect 296530 279420 296536 279472
rect 296588 279460 296594 279472
rect 351270 279460 351276 279472
rect 296588 279432 351276 279460
rect 296588 279420 296594 279432
rect 351270 279420 351276 279432
rect 351328 279420 351334 279472
rect 39942 278740 39948 278792
rect 40000 278780 40006 278792
rect 58618 278780 58624 278792
rect 40000 278752 58624 278780
rect 40000 278740 40006 278752
rect 58618 278740 58624 278752
rect 58676 278780 58682 278792
rect 58676 278752 59308 278780
rect 58676 278740 58682 278752
rect 59280 278712 59308 278752
rect 121454 278740 121460 278792
rect 121512 278780 121518 278792
rect 145558 278780 145564 278792
rect 121512 278752 145564 278780
rect 121512 278740 121518 278752
rect 145558 278740 145564 278752
rect 145616 278740 145622 278792
rect 67634 278712 67640 278724
rect 59280 278684 67640 278712
rect 67634 278672 67640 278684
rect 67692 278672 67698 278724
rect 121546 278672 121552 278724
rect 121604 278712 121610 278724
rect 132402 278712 132408 278724
rect 121604 278684 132408 278712
rect 121604 278672 121610 278684
rect 132402 278672 132408 278684
rect 132460 278672 132466 278724
rect 152642 278128 152648 278180
rect 152700 278168 152706 278180
rect 166718 278168 166724 278180
rect 152700 278140 166724 278168
rect 152700 278128 152706 278140
rect 166718 278128 166724 278140
rect 166776 278128 166782 278180
rect 132402 278060 132408 278112
rect 132460 278100 132466 278112
rect 164878 278100 164884 278112
rect 132460 278072 164884 278100
rect 132460 278060 132466 278072
rect 164878 278060 164884 278072
rect 164936 278060 164942 278112
rect 122742 277992 122748 278044
rect 122800 278032 122806 278044
rect 169202 278032 169208 278044
rect 122800 278004 169208 278032
rect 122800 277992 122806 278004
rect 169202 277992 169208 278004
rect 169260 277992 169266 278044
rect 305730 277992 305736 278044
rect 305788 278032 305794 278044
rect 371970 278032 371976 278044
rect 305788 278004 371976 278032
rect 305788 277992 305794 278004
rect 371970 277992 371976 278004
rect 372028 277992 372034 278044
rect 375190 277584 375196 277636
rect 375248 277624 375254 277636
rect 376754 277624 376760 277636
rect 375248 277596 376760 277624
rect 375248 277584 375254 277596
rect 376754 277584 376760 277596
rect 376812 277584 376818 277636
rect 53650 277380 53656 277432
rect 53708 277420 53714 277432
rect 67634 277420 67640 277432
rect 53708 277392 67640 277420
rect 53708 277380 53714 277392
rect 67634 277380 67640 277392
rect 67692 277380 67698 277432
rect 126422 277420 126428 277432
rect 125566 277392 126428 277420
rect 121454 277312 121460 277364
rect 121512 277352 121518 277364
rect 125566 277352 125594 277392
rect 126422 277380 126428 277392
rect 126480 277420 126486 277432
rect 142890 277420 142896 277432
rect 126480 277392 142896 277420
rect 126480 277380 126486 277392
rect 142890 277380 142896 277392
rect 142948 277380 142954 277432
rect 166718 277380 166724 277432
rect 166776 277420 166782 277432
rect 176654 277420 176660 277432
rect 166776 277392 176660 277420
rect 166776 277380 166782 277392
rect 176654 277380 176660 277392
rect 176712 277380 176718 277432
rect 373902 277380 373908 277432
rect 373960 277420 373966 277432
rect 375190 277420 375196 277432
rect 373960 277392 375196 277420
rect 373960 277380 373966 277392
rect 375190 277380 375196 277392
rect 375248 277380 375254 277432
rect 442626 277380 442632 277432
rect 442684 277420 442690 277432
rect 467926 277420 467932 277432
rect 442684 277392 467932 277420
rect 442684 277380 442690 277392
rect 467926 277380 467932 277392
rect 467984 277380 467990 277432
rect 121512 277324 125594 277352
rect 121512 277312 121518 277324
rect 299566 276740 299572 276752
rect 296686 276712 299572 276740
rect 56410 276632 56416 276684
rect 56468 276672 56474 276684
rect 67634 276672 67640 276684
rect 56468 276644 67640 276672
rect 56468 276632 56474 276644
rect 67634 276632 67640 276644
rect 67692 276632 67698 276684
rect 293034 276632 293040 276684
rect 293092 276672 293098 276684
rect 296686 276672 296714 276712
rect 299566 276700 299572 276712
rect 299624 276740 299630 276752
rect 300302 276740 300308 276752
rect 299624 276712 300308 276740
rect 299624 276700 299630 276712
rect 300302 276700 300308 276712
rect 300360 276700 300366 276752
rect 293092 276644 296714 276672
rect 293092 276632 293098 276644
rect 308490 276632 308496 276684
rect 308548 276672 308554 276684
rect 355502 276672 355508 276684
rect 308548 276644 355508 276672
rect 308548 276632 308554 276644
rect 355502 276632 355508 276644
rect 355560 276632 355566 276684
rect 46842 276020 46848 276072
rect 46900 276060 46906 276072
rect 67726 276060 67732 276072
rect 46900 276032 67732 276060
rect 46900 276020 46906 276032
rect 67726 276020 67732 276032
rect 67784 276020 67790 276072
rect 121454 276020 121460 276072
rect 121512 276060 121518 276072
rect 166258 276060 166264 276072
rect 121512 276032 166264 276060
rect 121512 276020 121518 276032
rect 166258 276020 166264 276032
rect 166316 276020 166322 276072
rect 371970 276020 371976 276072
rect 372028 276060 372034 276072
rect 377766 276060 377772 276072
rect 372028 276032 377772 276060
rect 372028 276020 372034 276032
rect 377766 276020 377772 276032
rect 377824 276020 377830 276072
rect 54846 275952 54852 276004
rect 54904 275992 54910 276004
rect 55122 275992 55128 276004
rect 54904 275964 55128 275992
rect 54904 275952 54910 275964
rect 55122 275952 55128 275964
rect 55180 275992 55186 276004
rect 67634 275992 67640 276004
rect 55180 275964 67640 275992
rect 55180 275952 55186 275964
rect 67634 275952 67640 275964
rect 67692 275952 67698 276004
rect 123662 275272 123668 275324
rect 123720 275312 123726 275324
rect 160094 275312 160100 275324
rect 123720 275284 160100 275312
rect 123720 275272 123726 275284
rect 160094 275272 160100 275284
rect 160152 275272 160158 275324
rect 301314 275272 301320 275324
rect 301372 275312 301378 275324
rect 376110 275312 376116 275324
rect 301372 275284 376116 275312
rect 301372 275272 301378 275284
rect 376110 275272 376116 275284
rect 376168 275272 376174 275324
rect 121454 274728 121460 274780
rect 121512 274768 121518 274780
rect 144454 274768 144460 274780
rect 121512 274740 144460 274768
rect 121512 274728 121518 274740
rect 144454 274728 144460 274740
rect 144512 274728 144518 274780
rect 160094 274728 160100 274780
rect 160152 274768 160158 274780
rect 161290 274768 161296 274780
rect 160152 274740 161296 274768
rect 160152 274728 160158 274740
rect 161290 274728 161296 274740
rect 161348 274768 161354 274780
rect 176654 274768 176660 274780
rect 161348 274740 176660 274768
rect 161348 274728 161354 274740
rect 176654 274728 176660 274740
rect 176712 274728 176718 274780
rect 121546 274660 121552 274712
rect 121604 274700 121610 274712
rect 170582 274700 170588 274712
rect 121604 274672 170588 274700
rect 121604 274660 121610 274672
rect 170582 274660 170588 274672
rect 170640 274660 170646 274712
rect 295334 274660 295340 274712
rect 295392 274700 295398 274712
rect 300854 274700 300860 274712
rect 295392 274672 300860 274700
rect 295392 274660 295398 274672
rect 300854 274660 300860 274672
rect 300912 274700 300918 274712
rect 301314 274700 301320 274712
rect 300912 274672 301320 274700
rect 300912 274660 300918 274672
rect 301314 274660 301320 274672
rect 301372 274660 301378 274712
rect 121454 274592 121460 274644
rect 121512 274632 121518 274644
rect 170490 274632 170496 274644
rect 121512 274604 170496 274632
rect 121512 274592 121518 274604
rect 170490 274592 170496 274604
rect 170548 274592 170554 274644
rect 41322 273912 41328 273964
rect 41380 273952 41386 273964
rect 56502 273952 56508 273964
rect 41380 273924 56508 273952
rect 41380 273912 41386 273924
rect 56502 273912 56508 273924
rect 56560 273912 56566 273964
rect 306282 273912 306288 273964
rect 306340 273952 306346 273964
rect 359642 273952 359648 273964
rect 306340 273924 359648 273952
rect 306340 273912 306346 273924
rect 359642 273912 359648 273924
rect 359700 273912 359706 273964
rect 463602 273912 463608 273964
rect 463660 273952 463666 273964
rect 531958 273952 531964 273964
rect 463660 273924 531964 273952
rect 463660 273912 463666 273924
rect 531958 273912 531964 273924
rect 532016 273912 532022 273964
rect 121454 273368 121460 273420
rect 121512 273408 121518 273420
rect 123478 273408 123484 273420
rect 121512 273380 123484 273408
rect 121512 273368 121518 273380
rect 123478 273368 123484 273380
rect 123536 273368 123542 273420
rect 66162 273300 66168 273352
rect 66220 273340 66226 273352
rect 67818 273340 67824 273352
rect 66220 273312 67824 273340
rect 66220 273300 66226 273312
rect 67818 273300 67824 273312
rect 67876 273300 67882 273352
rect 56226 273232 56232 273284
rect 56284 273272 56290 273284
rect 56502 273272 56508 273284
rect 56284 273244 56508 273272
rect 56284 273232 56290 273244
rect 56502 273232 56508 273244
rect 56560 273272 56566 273284
rect 67634 273272 67640 273284
rect 56560 273244 67640 273272
rect 56560 273232 56566 273244
rect 67634 273232 67640 273244
rect 67692 273232 67698 273284
rect 359642 273232 359648 273284
rect 359700 273272 359706 273284
rect 360010 273272 360016 273284
rect 359700 273244 360016 273272
rect 359700 273232 359706 273244
rect 360010 273232 360016 273244
rect 360068 273272 360074 273284
rect 377766 273272 377772 273284
rect 360068 273244 377772 273272
rect 360068 273232 360074 273244
rect 377766 273232 377772 273244
rect 377824 273232 377830 273284
rect 442718 273232 442724 273284
rect 442776 273272 442782 273284
rect 462314 273272 462320 273284
rect 442776 273244 462320 273272
rect 442776 273232 442782 273244
rect 462314 273232 462320 273244
rect 462372 273272 462378 273284
rect 463602 273272 463608 273284
rect 462372 273244 463608 273272
rect 462372 273232 462378 273244
rect 463602 273232 463608 273244
rect 463660 273232 463666 273284
rect 121454 272552 121460 272604
rect 121512 272592 121518 272604
rect 121638 272592 121644 272604
rect 121512 272564 121644 272592
rect 121512 272552 121518 272564
rect 121638 272552 121644 272564
rect 121696 272592 121702 272604
rect 143074 272592 143080 272604
rect 121696 272564 143080 272592
rect 121696 272552 121702 272564
rect 143074 272552 143080 272564
rect 143132 272552 143138 272604
rect 120810 272484 120816 272536
rect 120868 272524 120874 272536
rect 130562 272524 130568 272536
rect 120868 272496 130568 272524
rect 120868 272484 120874 272496
rect 130562 272484 130568 272496
rect 130620 272524 130626 272536
rect 158714 272524 158720 272536
rect 130620 272496 158720 272524
rect 130620 272484 130626 272496
rect 158714 272484 158720 272496
rect 158772 272484 158778 272536
rect 442810 272076 442816 272128
rect 442868 272116 442874 272128
rect 448606 272116 448612 272128
rect 442868 272088 448612 272116
rect 442868 272076 442874 272088
rect 448606 272076 448612 272088
rect 448664 272076 448670 272128
rect 66070 271872 66076 271924
rect 66128 271912 66134 271924
rect 67634 271912 67640 271924
rect 66128 271884 67640 271912
rect 66128 271872 66134 271884
rect 67634 271872 67640 271884
rect 67692 271872 67698 271924
rect 158714 271872 158720 271924
rect 158772 271912 158778 271924
rect 160002 271912 160008 271924
rect 158772 271884 160008 271912
rect 158772 271872 158778 271884
rect 160002 271872 160008 271884
rect 160060 271912 160066 271924
rect 176654 271912 176660 271924
rect 160060 271884 176660 271912
rect 160060 271872 160066 271884
rect 176654 271872 176660 271884
rect 176712 271872 176718 271924
rect 295334 271872 295340 271924
rect 295392 271912 295398 271924
rect 301682 271912 301688 271924
rect 295392 271884 301688 271912
rect 295392 271872 295398 271884
rect 301682 271872 301688 271884
rect 301740 271872 301746 271924
rect 176286 271804 176292 271856
rect 176344 271844 176350 271856
rect 179690 271844 179696 271856
rect 176344 271816 179696 271844
rect 176344 271804 176350 271816
rect 179690 271804 179696 271816
rect 179748 271804 179754 271856
rect 296530 271804 296536 271856
rect 296588 271844 296594 271856
rect 298094 271844 298100 271856
rect 296588 271816 298100 271844
rect 296588 271804 296594 271816
rect 298094 271804 298100 271816
rect 298152 271804 298158 271856
rect 64782 270580 64788 270632
rect 64840 270620 64846 270632
rect 67726 270620 67732 270632
rect 64840 270592 67732 270620
rect 64840 270580 64846 270592
rect 67726 270580 67732 270592
rect 67784 270580 67790 270632
rect 41322 270512 41328 270564
rect 41380 270552 41386 270564
rect 54478 270552 54484 270564
rect 41380 270524 54484 270552
rect 41380 270512 41386 270524
rect 54478 270512 54484 270524
rect 54536 270552 54542 270564
rect 54536 270524 55214 270552
rect 54536 270512 54542 270524
rect 55186 270484 55214 270524
rect 59170 270512 59176 270564
rect 59228 270552 59234 270564
rect 67634 270552 67640 270564
rect 59228 270524 67640 270552
rect 59228 270512 59234 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 121454 270512 121460 270564
rect 121512 270552 121518 270564
rect 152734 270552 152740 270564
rect 121512 270524 152740 270552
rect 121512 270512 121518 270524
rect 152734 270512 152740 270524
rect 152792 270512 152798 270564
rect 67726 270484 67732 270496
rect 55186 270456 67732 270484
rect 67726 270444 67732 270456
rect 67784 270444 67790 270496
rect 165522 269764 165528 269816
rect 165580 269804 165586 269816
rect 177298 269804 177304 269816
rect 165580 269776 177304 269804
rect 165580 269764 165586 269776
rect 177298 269764 177304 269776
rect 177356 269764 177362 269816
rect 121454 269152 121460 269204
rect 121512 269192 121518 269204
rect 130562 269192 130568 269204
rect 121512 269164 130568 269192
rect 121512 269152 121518 269164
rect 130562 269152 130568 269164
rect 130620 269152 130626 269204
rect 61838 269084 61844 269136
rect 61896 269124 61902 269136
rect 67634 269124 67640 269136
rect 61896 269096 67640 269124
rect 61896 269084 61902 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121546 269084 121552 269136
rect 121604 269124 121610 269136
rect 151262 269124 151268 269136
rect 121604 269096 151268 269124
rect 121604 269084 121610 269096
rect 151262 269084 151268 269096
rect 151320 269084 151326 269136
rect 442258 269084 442264 269136
rect 442316 269124 442322 269136
rect 448790 269124 448796 269136
rect 442316 269096 448796 269124
rect 442316 269084 442322 269096
rect 448790 269084 448796 269096
rect 448848 269084 448854 269136
rect 121454 269016 121460 269068
rect 121512 269056 121518 269068
rect 160738 269056 160744 269068
rect 121512 269028 160744 269056
rect 121512 269016 121518 269028
rect 160738 269016 160744 269028
rect 160796 269016 160802 269068
rect 126882 268948 126888 269000
rect 126940 268988 126946 269000
rect 130378 268988 130384 269000
rect 126940 268960 130384 268988
rect 126940 268948 126946 268960
rect 130378 268948 130384 268960
rect 130436 268948 130442 269000
rect 121362 268336 121368 268388
rect 121420 268376 121426 268388
rect 163682 268376 163688 268388
rect 121420 268348 163688 268376
rect 121420 268336 121426 268348
rect 163682 268336 163688 268348
rect 163740 268336 163746 268388
rect 294230 268336 294236 268388
rect 294288 268376 294294 268388
rect 299382 268376 299388 268388
rect 294288 268348 299388 268376
rect 294288 268336 294294 268348
rect 299382 268336 299388 268348
rect 299440 268376 299446 268388
rect 356698 268376 356704 268388
rect 299440 268348 356704 268376
rect 299440 268336 299446 268348
rect 356698 268336 356704 268348
rect 356756 268336 356762 268388
rect 35710 267792 35716 267844
rect 35768 267832 35774 267844
rect 67634 267832 67640 267844
rect 35768 267804 67640 267832
rect 35768 267792 35774 267804
rect 67634 267792 67640 267804
rect 67692 267792 67698 267844
rect 8202 267764 8208 267776
rect 6932 267736 8208 267764
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 6932 267696 6960 267736
rect 8202 267724 8208 267736
rect 8260 267764 8266 267776
rect 48958 267764 48964 267776
rect 8260 267736 48964 267764
rect 8260 267724 8266 267736
rect 48958 267724 48964 267736
rect 49016 267724 49022 267776
rect 53466 267724 53472 267776
rect 53524 267764 53530 267776
rect 67726 267764 67732 267776
rect 53524 267736 67732 267764
rect 53524 267724 53530 267736
rect 67726 267724 67732 267736
rect 67784 267724 67790 267776
rect 121454 267724 121460 267776
rect 121512 267764 121518 267776
rect 126882 267764 126888 267776
rect 121512 267736 126888 267764
rect 121512 267724 121518 267736
rect 126882 267724 126888 267736
rect 126940 267724 126946 267776
rect 161382 267724 161388 267776
rect 161440 267764 161446 267776
rect 176654 267764 176660 267776
rect 161440 267736 176660 267764
rect 161440 267724 161446 267736
rect 176654 267724 176660 267736
rect 176712 267724 176718 267776
rect 3568 267668 6960 267696
rect 3568 267656 3574 267668
rect 45278 267656 45284 267708
rect 45336 267696 45342 267708
rect 67634 267696 67640 267708
rect 45336 267668 67640 267696
rect 45336 267656 45342 267668
rect 67634 267656 67640 267668
rect 67692 267656 67698 267708
rect 301498 267656 301504 267708
rect 301556 267696 301562 267708
rect 379238 267696 379244 267708
rect 301556 267668 379244 267696
rect 301556 267656 301562 267668
rect 379238 267656 379244 267668
rect 379296 267656 379302 267708
rect 59078 267588 59084 267640
rect 59136 267628 59142 267640
rect 67726 267628 67732 267640
rect 59136 267600 67732 267628
rect 59136 267588 59142 267600
rect 67726 267588 67732 267600
rect 67784 267588 67790 267640
rect 125042 267044 125048 267096
rect 125100 267084 125106 267096
rect 169018 267084 169024 267096
rect 125100 267056 169024 267084
rect 125100 267044 125106 267056
rect 169018 267044 169024 267056
rect 169076 267044 169082 267096
rect 122466 266976 122472 267028
rect 122524 267016 122530 267028
rect 169294 267016 169300 267028
rect 122524 266988 169300 267016
rect 122524 266976 122530 266988
rect 169294 266976 169300 266988
rect 169352 266976 169358 267028
rect 442810 266364 442816 266416
rect 442868 266404 442874 266416
rect 460198 266404 460204 266416
rect 442868 266376 460204 266404
rect 442868 266364 442874 266376
rect 460198 266364 460204 266376
rect 460256 266404 460262 266416
rect 460256 266376 460934 266404
rect 460256 266364 460262 266376
rect 49418 266296 49424 266348
rect 49476 266336 49482 266348
rect 67634 266336 67640 266348
rect 49476 266308 67640 266336
rect 49476 266296 49482 266308
rect 67634 266296 67640 266308
rect 67692 266296 67698 266348
rect 152550 266296 152556 266348
rect 152608 266336 152614 266348
rect 176654 266336 176660 266348
rect 152608 266308 176660 266336
rect 152608 266296 152614 266308
rect 176654 266296 176660 266308
rect 176712 266296 176718 266348
rect 460906 266336 460934 266376
rect 542354 266336 542360 266348
rect 460906 266308 542360 266336
rect 542354 266296 542360 266308
rect 542412 266296 542418 266348
rect 133322 265684 133328 265736
rect 133380 265724 133386 265736
rect 163498 265724 163504 265736
rect 133380 265696 163504 265724
rect 133380 265684 133386 265696
rect 163498 265684 163504 265696
rect 163556 265684 163562 265736
rect 121454 265616 121460 265668
rect 121512 265656 121518 265668
rect 125502 265656 125508 265668
rect 121512 265628 125508 265656
rect 121512 265616 121518 265628
rect 125502 265616 125508 265628
rect 125560 265656 125566 265668
rect 174538 265656 174544 265668
rect 125560 265628 174544 265656
rect 125560 265616 125566 265628
rect 174538 265616 174544 265628
rect 174596 265616 174602 265668
rect 442350 265072 442356 265124
rect 442408 265112 442414 265124
rect 444650 265112 444656 265124
rect 442408 265084 444656 265112
rect 442408 265072 442414 265084
rect 444650 265072 444656 265084
rect 444708 265072 444714 265124
rect 364150 264936 364156 264988
rect 364208 264976 364214 264988
rect 376938 264976 376944 264988
rect 364208 264948 376944 264976
rect 364208 264936 364214 264948
rect 376938 264936 376944 264948
rect 376996 264936 377002 264988
rect 49510 263644 49516 263696
rect 49568 263684 49574 263696
rect 67634 263684 67640 263696
rect 49568 263656 67640 263684
rect 49568 263644 49574 263656
rect 67634 263644 67640 263656
rect 67692 263644 67698 263696
rect 8938 263576 8944 263628
rect 8996 263616 9002 263628
rect 54846 263616 54852 263628
rect 8996 263588 54852 263616
rect 8996 263576 9002 263588
rect 54846 263576 54852 263588
rect 54904 263616 54910 263628
rect 67726 263616 67732 263628
rect 54904 263588 67732 263616
rect 54904 263576 54910 263588
rect 67726 263576 67732 263588
rect 67784 263576 67790 263628
rect 121454 263576 121460 263628
rect 121512 263616 121518 263628
rect 171870 263616 171876 263628
rect 121512 263588 171876 263616
rect 121512 263576 121518 263588
rect 171870 263576 171876 263588
rect 171928 263576 171934 263628
rect 376570 263576 376576 263628
rect 376628 263616 376634 263628
rect 377490 263616 377496 263628
rect 376628 263588 377496 263616
rect 376628 263576 376634 263588
rect 377490 263576 377496 263588
rect 377548 263576 377554 263628
rect 121546 263508 121552 263560
rect 121604 263548 121610 263560
rect 132494 263548 132500 263560
rect 121604 263520 132500 263548
rect 121604 263508 121610 263520
rect 132494 263508 132500 263520
rect 132552 263548 132558 263560
rect 133782 263548 133788 263560
rect 132552 263520 133788 263548
rect 132552 263508 132558 263520
rect 133782 263508 133788 263520
rect 133840 263508 133846 263560
rect 296346 263508 296352 263560
rect 296404 263548 296410 263560
rect 345750 263548 345756 263560
rect 296404 263520 345756 263548
rect 296404 263508 296410 263520
rect 345750 263508 345756 263520
rect 345808 263508 345814 263560
rect 353938 263508 353944 263560
rect 353996 263548 354002 263560
rect 377306 263548 377312 263560
rect 353996 263520 377312 263548
rect 353996 263508 354002 263520
rect 377306 263508 377312 263520
rect 377364 263508 377370 263560
rect 121454 262828 121460 262880
rect 121512 262868 121518 262880
rect 153194 262868 153200 262880
rect 121512 262840 153200 262868
rect 121512 262828 121518 262840
rect 153194 262828 153200 262840
rect 153252 262868 153258 262880
rect 153930 262868 153936 262880
rect 153252 262840 153936 262868
rect 153252 262828 153258 262840
rect 153930 262828 153936 262840
rect 153988 262828 153994 262880
rect 60366 262284 60372 262336
rect 60424 262324 60430 262336
rect 67726 262324 67732 262336
rect 60424 262296 67732 262324
rect 60424 262284 60430 262296
rect 67726 262284 67732 262296
rect 67784 262284 67790 262336
rect 55122 262216 55128 262268
rect 55180 262256 55186 262268
rect 67634 262256 67640 262268
rect 55180 262228 67640 262256
rect 55180 262216 55186 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 442718 262216 442724 262268
rect 442776 262256 442782 262268
rect 467098 262256 467104 262268
rect 442776 262228 467104 262256
rect 442776 262216 442782 262228
rect 467098 262216 467104 262228
rect 467156 262216 467162 262268
rect 60550 262148 60556 262200
rect 60608 262188 60614 262200
rect 67726 262188 67732 262200
rect 60608 262160 67732 262188
rect 60608 262148 60614 262160
rect 67726 262148 67732 262160
rect 67784 262148 67790 262200
rect 121454 262148 121460 262200
rect 121512 262188 121518 262200
rect 171134 262188 171140 262200
rect 121512 262160 171140 262188
rect 121512 262148 121518 262160
rect 171134 262148 171140 262160
rect 171192 262148 171198 262200
rect 302878 262148 302884 262200
rect 302936 262188 302942 262200
rect 303706 262188 303712 262200
rect 302936 262160 303712 262188
rect 302936 262148 302942 262160
rect 303706 262148 303712 262160
rect 303764 262148 303770 262200
rect 61930 262080 61936 262132
rect 61988 262120 61994 262132
rect 67634 262120 67640 262132
rect 61988 262092 67640 262120
rect 61988 262080 61994 262092
rect 67634 262080 67640 262092
rect 67692 262080 67698 262132
rect 158162 261468 158168 261520
rect 158220 261508 158226 261520
rect 158622 261508 158628 261520
rect 158220 261480 158628 261508
rect 158220 261468 158226 261480
rect 158622 261468 158628 261480
rect 158680 261508 158686 261520
rect 176654 261508 176660 261520
rect 158680 261480 176660 261508
rect 158680 261468 158686 261480
rect 176654 261468 176660 261480
rect 176712 261468 176718 261520
rect 442810 261468 442816 261520
rect 442868 261508 442874 261520
rect 570598 261508 570604 261520
rect 442868 261480 570604 261508
rect 442868 261468 442874 261480
rect 570598 261468 570604 261480
rect 570656 261468 570662 261520
rect 295334 261128 295340 261180
rect 295392 261168 295398 261180
rect 299382 261168 299388 261180
rect 295392 261140 299388 261168
rect 295392 261128 295398 261140
rect 299382 261128 299388 261140
rect 299440 261168 299446 261180
rect 304442 261168 304448 261180
rect 299440 261140 304448 261168
rect 299440 261128 299446 261140
rect 304442 261128 304448 261140
rect 304500 261128 304506 261180
rect 303706 260856 303712 260908
rect 303764 260896 303770 260908
rect 379330 260896 379336 260908
rect 303764 260868 379336 260896
rect 303764 260856 303770 260868
rect 379330 260856 379336 260868
rect 379388 260856 379394 260908
rect 21358 260788 21364 260840
rect 21416 260828 21422 260840
rect 67634 260828 67640 260840
rect 21416 260800 67640 260828
rect 21416 260788 21422 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 121454 260788 121460 260840
rect 121512 260828 121518 260840
rect 127158 260828 127164 260840
rect 121512 260800 127164 260828
rect 121512 260788 121518 260800
rect 127158 260788 127164 260800
rect 127216 260828 127222 260840
rect 127434 260828 127440 260840
rect 127216 260800 127440 260828
rect 127216 260788 127222 260800
rect 127434 260788 127440 260800
rect 127492 260788 127498 260840
rect 63310 260720 63316 260772
rect 63368 260760 63374 260772
rect 67726 260760 67732 260772
rect 63368 260732 67732 260760
rect 63368 260720 63374 260732
rect 67726 260720 67732 260732
rect 67784 260720 67790 260772
rect 127434 260176 127440 260228
rect 127492 260216 127498 260228
rect 149974 260216 149980 260228
rect 127492 260188 149980 260216
rect 127492 260176 127498 260188
rect 149974 260176 149980 260188
rect 150032 260176 150038 260228
rect 121638 260108 121644 260160
rect 121696 260148 121702 260160
rect 167822 260148 167828 260160
rect 121696 260120 167828 260148
rect 121696 260108 121702 260120
rect 167822 260108 167828 260120
rect 167880 260108 167886 260160
rect 121454 259428 121460 259480
rect 121512 259468 121518 259480
rect 131942 259468 131948 259480
rect 121512 259440 131948 259468
rect 121512 259428 121518 259440
rect 131942 259428 131948 259440
rect 132000 259428 132006 259480
rect 293862 259360 293868 259412
rect 293920 259400 293926 259412
rect 308398 259400 308404 259412
rect 293920 259372 308404 259400
rect 293920 259360 293926 259372
rect 308398 259360 308404 259372
rect 308456 259360 308462 259412
rect 365254 259360 365260 259412
rect 365312 259400 365318 259412
rect 371050 259400 371056 259412
rect 365312 259372 371056 259400
rect 365312 259360 365318 259372
rect 371050 259360 371056 259372
rect 371108 259360 371114 259412
rect 440234 259360 440240 259412
rect 440292 259400 440298 259412
rect 454034 259400 454040 259412
rect 440292 259372 454040 259400
rect 440292 259360 440298 259372
rect 454034 259360 454040 259372
rect 454092 259360 454098 259412
rect 446490 259292 446496 259344
rect 446548 259332 446554 259344
rect 448606 259332 448612 259344
rect 446548 259304 448612 259332
rect 446548 259292 446554 259304
rect 448606 259292 448612 259304
rect 448664 259292 448670 259344
rect 3970 258680 3976 258732
rect 4028 258720 4034 258732
rect 62850 258720 62856 258732
rect 4028 258692 62856 258720
rect 4028 258680 4034 258692
rect 62850 258680 62856 258692
rect 62908 258680 62914 258732
rect 57790 258068 57796 258120
rect 57848 258108 57854 258120
rect 67726 258108 67732 258120
rect 57848 258080 67732 258108
rect 57848 258068 57854 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 121454 258068 121460 258120
rect 121512 258108 121518 258120
rect 156690 258108 156696 258120
rect 121512 258080 156696 258108
rect 121512 258068 121518 258080
rect 156690 258068 156696 258080
rect 156748 258068 156754 258120
rect 371050 258068 371056 258120
rect 371108 258108 371114 258120
rect 376938 258108 376944 258120
rect 371108 258080 376944 258108
rect 371108 258068 371114 258080
rect 376938 258068 376944 258080
rect 376996 258068 377002 258120
rect 448606 258068 448612 258120
rect 448664 258108 448670 258120
rect 580166 258108 580172 258120
rect 448664 258080 580172 258108
rect 448664 258068 448670 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 53742 258000 53748 258052
rect 53800 258040 53806 258052
rect 67634 258040 67640 258052
rect 53800 258012 67640 258040
rect 53800 258000 53806 258012
rect 67634 258000 67640 258012
rect 67692 258000 67698 258052
rect 18598 257320 18604 257372
rect 18656 257360 18662 257372
rect 53742 257360 53748 257372
rect 18656 257332 53748 257360
rect 18656 257320 18662 257332
rect 53742 257320 53748 257332
rect 53800 257320 53806 257372
rect 121454 256776 121460 256828
rect 121512 256816 121518 256828
rect 150066 256816 150072 256828
rect 121512 256788 150072 256816
rect 121512 256776 121518 256788
rect 150066 256776 150072 256788
rect 150124 256776 150130 256828
rect 121546 256708 121552 256760
rect 121604 256748 121610 256760
rect 162302 256748 162308 256760
rect 121604 256720 162308 256748
rect 121604 256708 121610 256720
rect 162302 256708 162308 256720
rect 162360 256708 162366 256760
rect 176654 256748 176660 256760
rect 174924 256720 176660 256748
rect 140590 256640 140596 256692
rect 140648 256680 140654 256692
rect 174924 256680 174952 256720
rect 176654 256708 176660 256720
rect 176712 256708 176718 256760
rect 295334 256708 295340 256760
rect 295392 256748 295398 256760
rect 302326 256748 302332 256760
rect 295392 256720 302332 256748
rect 295392 256708 295398 256720
rect 302326 256708 302332 256720
rect 302384 256748 302390 256760
rect 379882 256748 379888 256760
rect 302384 256720 379888 256748
rect 302384 256708 302390 256720
rect 379882 256708 379888 256720
rect 379940 256708 379946 256760
rect 440510 256708 440516 256760
rect 440568 256748 440574 256760
rect 446490 256748 446496 256760
rect 440568 256720 446496 256748
rect 440568 256708 440574 256720
rect 446490 256708 446496 256720
rect 446548 256708 446554 256760
rect 140648 256652 174952 256680
rect 140648 256640 140654 256652
rect 121454 256096 121460 256148
rect 121512 256136 121518 256148
rect 127066 256136 127072 256148
rect 121512 256108 127072 256136
rect 121512 256096 121518 256108
rect 127066 256096 127072 256108
rect 127124 256096 127130 256148
rect 122190 256028 122196 256080
rect 122248 256068 122254 256080
rect 130378 256068 130384 256080
rect 122248 256040 130384 256068
rect 122248 256028 122254 256040
rect 130378 256028 130384 256040
rect 130436 256028 130442 256080
rect 63402 255960 63408 256012
rect 63460 256000 63466 256012
rect 67634 256000 67640 256012
rect 63460 255972 67640 256000
rect 63460 255960 63466 255972
rect 67634 255960 67640 255972
rect 67692 255960 67698 256012
rect 122466 255960 122472 256012
rect 122524 256000 122530 256012
rect 155310 256000 155316 256012
rect 122524 255972 155316 256000
rect 122524 255960 122530 255972
rect 155310 255960 155316 255972
rect 155368 255960 155374 256012
rect 318610 255960 318616 256012
rect 318668 256000 318674 256012
rect 377306 256000 377312 256012
rect 318668 255972 377312 256000
rect 318668 255960 318674 255972
rect 377306 255960 377312 255972
rect 377364 255960 377370 256012
rect 127066 255348 127072 255400
rect 127124 255388 127130 255400
rect 127618 255388 127624 255400
rect 127124 255360 127624 255388
rect 127124 255348 127130 255360
rect 127618 255348 127624 255360
rect 127676 255348 127682 255400
rect 60550 255280 60556 255332
rect 60608 255320 60614 255332
rect 67726 255320 67732 255332
rect 60608 255292 67732 255320
rect 60608 255280 60614 255292
rect 67726 255280 67732 255292
rect 67784 255280 67790 255332
rect 121454 255280 121460 255332
rect 121512 255320 121518 255332
rect 152642 255320 152648 255332
rect 121512 255292 152648 255320
rect 121512 255280 121518 255292
rect 152642 255280 152648 255292
rect 152700 255280 152706 255332
rect 166626 255212 166632 255264
rect 166684 255252 166690 255264
rect 176654 255252 176660 255264
rect 166684 255224 176660 255252
rect 166684 255212 166690 255224
rect 176654 255212 176660 255224
rect 176712 255212 176718 255264
rect 295334 254532 295340 254584
rect 295392 254572 295398 254584
rect 300118 254572 300124 254584
rect 295392 254544 300124 254572
rect 295392 254532 295398 254544
rect 300118 254532 300124 254544
rect 300176 254572 300182 254584
rect 300762 254572 300768 254584
rect 300176 254544 300768 254572
rect 300176 254532 300182 254544
rect 300762 254532 300768 254544
rect 300820 254532 300826 254584
rect 61654 253988 61660 254040
rect 61712 254028 61718 254040
rect 67634 254028 67640 254040
rect 61712 254000 67640 254028
rect 61712 253988 61718 254000
rect 67634 253988 67640 254000
rect 67692 253988 67698 254040
rect 123662 253988 123668 254040
rect 123720 254028 123726 254040
rect 164142 254028 164148 254040
rect 123720 254000 164148 254028
rect 123720 253988 123726 254000
rect 164142 253988 164148 254000
rect 164200 254028 164206 254040
rect 166626 254028 166632 254040
rect 164200 254000 166632 254028
rect 164200 253988 164206 254000
rect 166626 253988 166632 254000
rect 166684 253988 166690 254040
rect 61930 253920 61936 253972
rect 61988 253960 61994 253972
rect 67726 253960 67732 253972
rect 61988 253932 67732 253960
rect 61988 253920 61994 253932
rect 67726 253920 67732 253932
rect 67784 253920 67790 253972
rect 121454 253920 121460 253972
rect 121512 253960 121518 253972
rect 173158 253960 173164 253972
rect 121512 253932 173164 253960
rect 121512 253920 121518 253932
rect 173158 253920 173164 253932
rect 173216 253920 173222 253972
rect 36814 253852 36820 253904
rect 36872 253892 36878 253904
rect 36998 253892 37004 253904
rect 36872 253864 37004 253892
rect 36872 253852 36878 253864
rect 36998 253852 37004 253864
rect 37056 253892 37062 253904
rect 67634 253892 67640 253904
rect 37056 253864 67640 253892
rect 37056 253852 37062 253864
rect 67634 253852 67640 253864
rect 67692 253852 67698 253904
rect 121546 253852 121552 253904
rect 121604 253892 121610 253904
rect 140038 253892 140044 253904
rect 121604 253864 140044 253892
rect 121604 253852 121610 253864
rect 140038 253852 140044 253864
rect 140096 253852 140102 253904
rect 4798 253172 4804 253224
rect 4856 253212 4862 253224
rect 36814 253212 36820 253224
rect 4856 253184 36820 253212
rect 4856 253172 4862 253184
rect 36814 253172 36820 253184
rect 36872 253172 36878 253224
rect 300762 253172 300768 253224
rect 300820 253212 300826 253224
rect 373258 253212 373264 253224
rect 300820 253184 373264 253212
rect 300820 253172 300826 253184
rect 373258 253172 373264 253184
rect 373316 253172 373322 253224
rect 64506 252560 64512 252612
rect 64564 252600 64570 252612
rect 66898 252600 66904 252612
rect 64564 252572 66904 252600
rect 64564 252560 64570 252572
rect 66898 252560 66904 252572
rect 66956 252600 66962 252612
rect 67542 252600 67548 252612
rect 66956 252572 67548 252600
rect 66956 252560 66962 252572
rect 67542 252560 67548 252572
rect 67600 252560 67606 252612
rect 121454 252560 121460 252612
rect 121512 252600 121518 252612
rect 158162 252600 158168 252612
rect 121512 252572 158168 252600
rect 121512 252560 121518 252572
rect 158162 252560 158168 252572
rect 158220 252560 158226 252612
rect 62022 252492 62028 252544
rect 62080 252532 62086 252544
rect 67634 252532 67640 252544
rect 62080 252504 67640 252532
rect 62080 252492 62086 252504
rect 67634 252492 67640 252504
rect 67692 252492 67698 252544
rect 296622 251880 296628 251932
rect 296680 251920 296686 251932
rect 311158 251920 311164 251932
rect 296680 251892 311164 251920
rect 296680 251880 296686 251892
rect 311158 251880 311164 251892
rect 311216 251880 311222 251932
rect 56410 251812 56416 251864
rect 56468 251852 56474 251864
rect 68278 251852 68284 251864
rect 56468 251824 68284 251852
rect 56468 251812 56474 251824
rect 68278 251812 68284 251824
rect 68336 251812 68342 251864
rect 297450 251812 297456 251864
rect 297508 251852 297514 251864
rect 368290 251852 368296 251864
rect 297508 251824 368296 251852
rect 297508 251812 297514 251824
rect 368290 251812 368296 251824
rect 368348 251812 368354 251864
rect 442902 251812 442908 251864
rect 442960 251852 442966 251864
rect 448514 251852 448520 251864
rect 442960 251824 448520 251852
rect 442960 251812 442966 251824
rect 448514 251812 448520 251824
rect 448572 251852 448578 251864
rect 462406 251852 462412 251864
rect 448572 251824 462412 251852
rect 448572 251812 448578 251824
rect 462406 251812 462412 251824
rect 462464 251812 462470 251864
rect 295334 251744 295340 251796
rect 295392 251784 295398 251796
rect 297358 251784 297364 251796
rect 295392 251756 297364 251784
rect 295392 251744 295398 251756
rect 297358 251744 297364 251756
rect 297416 251744 297422 251796
rect 121546 251268 121552 251320
rect 121604 251308 121610 251320
rect 159542 251308 159548 251320
rect 121604 251280 159548 251308
rect 121604 251268 121610 251280
rect 159542 251268 159548 251280
rect 159600 251268 159606 251320
rect 121454 251200 121460 251252
rect 121512 251240 121518 251252
rect 170674 251240 170680 251252
rect 121512 251212 170680 251240
rect 121512 251200 121518 251212
rect 170674 251200 170680 251212
rect 170732 251200 170738 251252
rect 368290 251200 368296 251252
rect 368348 251240 368354 251252
rect 376938 251240 376944 251252
rect 368348 251212 376944 251240
rect 368348 251200 368354 251212
rect 376938 251200 376944 251212
rect 376996 251200 377002 251252
rect 442718 251200 442724 251252
rect 442776 251240 442782 251252
rect 460934 251240 460940 251252
rect 442776 251212 460940 251240
rect 442776 251200 442782 251212
rect 460934 251200 460940 251212
rect 460992 251200 460998 251252
rect 120626 251132 120632 251184
rect 120684 251172 120690 251184
rect 132586 251172 132592 251184
rect 120684 251144 132592 251172
rect 120684 251132 120690 251144
rect 132586 251132 132592 251144
rect 132644 251132 132650 251184
rect 295334 250452 295340 250504
rect 295392 250492 295398 250504
rect 296622 250492 296628 250504
rect 295392 250464 296628 250492
rect 295392 250452 295398 250464
rect 296622 250452 296628 250464
rect 296680 250492 296686 250504
rect 300118 250492 300124 250504
rect 296680 250464 300124 250492
rect 296680 250452 296686 250464
rect 300118 250452 300124 250464
rect 300176 250452 300182 250504
rect 57698 249840 57704 249892
rect 57756 249880 57762 249892
rect 67634 249880 67640 249892
rect 57756 249852 67640 249880
rect 57756 249840 57762 249852
rect 67634 249840 67640 249852
rect 67692 249840 67698 249892
rect 121454 249772 121460 249824
rect 121512 249812 121518 249824
rect 133230 249812 133236 249824
rect 121512 249784 133236 249812
rect 121512 249772 121518 249784
rect 133230 249772 133236 249784
rect 133288 249772 133294 249824
rect 52270 249704 52276 249756
rect 52328 249744 52334 249756
rect 67634 249744 67640 249756
rect 52328 249716 67640 249744
rect 52328 249704 52334 249716
rect 67634 249704 67640 249716
rect 67692 249704 67698 249756
rect 121546 249704 121552 249756
rect 121604 249744 121610 249756
rect 129734 249744 129740 249756
rect 121604 249716 129740 249744
rect 121604 249704 121610 249716
rect 129734 249704 129740 249716
rect 129792 249704 129798 249756
rect 121454 249636 121460 249688
rect 121512 249676 121518 249688
rect 129182 249676 129188 249688
rect 121512 249648 129188 249676
rect 121512 249636 121518 249648
rect 129182 249636 129188 249648
rect 129240 249636 129246 249688
rect 119798 249092 119804 249144
rect 119856 249132 119862 249144
rect 130654 249132 130660 249144
rect 119856 249104 130660 249132
rect 119856 249092 119862 249104
rect 130654 249092 130660 249104
rect 130712 249092 130718 249144
rect 129734 249024 129740 249076
rect 129792 249064 129798 249076
rect 175918 249064 175924 249076
rect 129792 249036 175924 249064
rect 129792 249024 129798 249036
rect 175918 249024 175924 249036
rect 175976 249024 175982 249076
rect 65794 248616 65800 248668
rect 65852 248656 65858 248668
rect 68002 248656 68008 248668
rect 65852 248628 68008 248656
rect 65852 248616 65858 248628
rect 68002 248616 68008 248628
rect 68060 248616 68066 248668
rect 121454 248344 121460 248396
rect 121512 248384 121518 248396
rect 162118 248384 162124 248396
rect 121512 248356 162124 248384
rect 121512 248344 121518 248356
rect 162118 248344 162124 248356
rect 162176 248344 162182 248396
rect 295334 248344 295340 248396
rect 295392 248384 295398 248396
rect 316126 248384 316132 248396
rect 295392 248356 316132 248384
rect 295392 248344 295398 248356
rect 316126 248344 316132 248356
rect 316184 248384 316190 248396
rect 317230 248384 317236 248396
rect 316184 248356 317236 248384
rect 316184 248344 316190 248356
rect 317230 248344 317236 248356
rect 317288 248344 317294 248396
rect 317230 247664 317236 247716
rect 317288 247704 317294 247716
rect 373350 247704 373356 247716
rect 317288 247676 373356 247704
rect 317288 247664 317294 247676
rect 373350 247664 373356 247676
rect 373408 247664 373414 247716
rect 63218 247120 63224 247172
rect 63276 247160 63282 247172
rect 67634 247160 67640 247172
rect 63276 247132 67640 247160
rect 63276 247120 63282 247132
rect 67634 247120 67640 247132
rect 67692 247120 67698 247172
rect 59078 247052 59084 247104
rect 59136 247092 59142 247104
rect 67726 247092 67732 247104
rect 59136 247064 67732 247092
rect 59136 247052 59142 247064
rect 67726 247052 67732 247064
rect 67784 247052 67790 247104
rect 121546 247052 121552 247104
rect 121604 247092 121610 247104
rect 129182 247092 129188 247104
rect 121604 247064 129188 247092
rect 121604 247052 121610 247064
rect 129182 247052 129188 247064
rect 129240 247052 129246 247104
rect 362954 247052 362960 247104
rect 363012 247092 363018 247104
rect 376938 247092 376944 247104
rect 363012 247064 376944 247092
rect 363012 247052 363018 247064
rect 376938 247052 376944 247064
rect 376996 247052 377002 247104
rect 50798 246984 50804 247036
rect 50856 247024 50862 247036
rect 67634 247024 67640 247036
rect 50856 246996 67640 247024
rect 50856 246984 50862 246996
rect 67634 246984 67640 246996
rect 67692 246984 67698 247036
rect 65978 246916 65984 246968
rect 66036 246956 66042 246968
rect 68094 246956 68100 246968
rect 66036 246928 68100 246956
rect 66036 246916 66042 246928
rect 68094 246916 68100 246928
rect 68152 246916 68158 246968
rect 301038 246508 301044 246560
rect 301096 246548 301102 246560
rect 301590 246548 301596 246560
rect 301096 246520 301596 246548
rect 301096 246508 301102 246520
rect 301590 246508 301596 246520
rect 301648 246508 301654 246560
rect 294322 246304 294328 246356
rect 294380 246344 294386 246356
rect 301038 246344 301044 246356
rect 294380 246316 301044 246344
rect 294380 246304 294386 246316
rect 301038 246304 301044 246316
rect 301096 246304 301102 246356
rect 318702 246304 318708 246356
rect 318760 246344 318766 246356
rect 362954 246344 362960 246356
rect 318760 246316 362960 246344
rect 318760 246304 318766 246316
rect 362954 246304 362960 246316
rect 363012 246344 363018 246356
rect 363690 246344 363696 246356
rect 363012 246316 363696 246344
rect 363012 246304 363018 246316
rect 363690 246304 363696 246316
rect 363748 246304 363754 246356
rect 442902 246304 442908 246356
rect 442960 246344 442966 246356
rect 534074 246344 534080 246356
rect 442960 246316 534080 246344
rect 442960 246304 442966 246316
rect 534074 246304 534080 246316
rect 534132 246304 534138 246356
rect 121546 245760 121552 245812
rect 121604 245800 121610 245812
rect 124950 245800 124956 245812
rect 121604 245772 124956 245800
rect 121604 245760 121610 245772
rect 124950 245760 124956 245772
rect 125008 245760 125014 245812
rect 121454 245692 121460 245744
rect 121512 245732 121518 245744
rect 148410 245732 148416 245744
rect 121512 245704 148416 245732
rect 121512 245692 121518 245704
rect 148410 245692 148416 245704
rect 148468 245692 148474 245744
rect 131850 245624 131856 245676
rect 131908 245664 131914 245676
rect 164050 245664 164056 245676
rect 131908 245636 164056 245664
rect 131908 245624 131914 245636
rect 164050 245624 164056 245636
rect 164108 245664 164114 245676
rect 176654 245664 176660 245676
rect 164108 245636 176660 245664
rect 164108 245624 164114 245636
rect 176654 245624 176660 245636
rect 176712 245624 176718 245676
rect 318058 245624 318064 245676
rect 318116 245664 318122 245676
rect 318702 245664 318708 245676
rect 318116 245636 318708 245664
rect 318116 245624 318122 245636
rect 318702 245624 318708 245636
rect 318760 245624 318766 245676
rect 364702 245624 364708 245676
rect 364760 245664 364766 245676
rect 365622 245664 365628 245676
rect 364760 245636 365628 245664
rect 364760 245624 364766 245636
rect 365622 245624 365628 245636
rect 365680 245664 365686 245676
rect 376938 245664 376944 245676
rect 365680 245636 376944 245664
rect 365680 245624 365686 245636
rect 376938 245624 376944 245636
rect 376996 245624 377002 245676
rect 26142 245556 26148 245608
rect 26200 245596 26206 245608
rect 67634 245596 67640 245608
rect 26200 245568 67640 245596
rect 26200 245556 26206 245568
rect 67634 245556 67640 245568
rect 67692 245556 67698 245608
rect 121454 245556 121460 245608
rect 121512 245596 121518 245608
rect 166994 245596 167000 245608
rect 121512 245568 167000 245596
rect 121512 245556 121518 245568
rect 166994 245556 167000 245568
rect 167052 245556 167058 245608
rect 467098 245556 467104 245608
rect 467156 245596 467162 245608
rect 533982 245596 533988 245608
rect 467156 245568 533988 245596
rect 467156 245556 467162 245568
rect 533982 245556 533988 245568
rect 534040 245596 534046 245608
rect 580166 245596 580172 245608
rect 534040 245568 580172 245596
rect 534040 245556 534046 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 121546 244264 121552 244316
rect 121604 244304 121610 244316
rect 147490 244304 147496 244316
rect 121604 244276 147496 244304
rect 121604 244264 121610 244276
rect 147490 244264 147496 244276
rect 147548 244264 147554 244316
rect 35802 244196 35808 244248
rect 35860 244236 35866 244248
rect 67634 244236 67640 244248
rect 35860 244208 67640 244236
rect 35860 244196 35866 244208
rect 67634 244196 67640 244208
rect 67692 244196 67698 244248
rect 121638 244196 121644 244248
rect 121696 244236 121702 244248
rect 135990 244236 135996 244248
rect 121696 244208 135996 244236
rect 121696 244196 121702 244208
rect 135990 244196 135996 244208
rect 136048 244196 136054 244248
rect 17218 244128 17224 244180
rect 17276 244168 17282 244180
rect 43990 244168 43996 244180
rect 17276 244140 43996 244168
rect 17276 244128 17282 244140
rect 43990 244128 43996 244140
rect 44048 244168 44054 244180
rect 67726 244168 67732 244180
rect 44048 244140 67732 244168
rect 44048 244128 44054 244140
rect 67726 244128 67732 244140
rect 67784 244128 67790 244180
rect 121454 244128 121460 244180
rect 121512 244168 121518 244180
rect 126238 244168 126244 244180
rect 121512 244140 126244 244168
rect 121512 244128 121518 244140
rect 126238 244128 126244 244140
rect 126296 244128 126302 244180
rect 159450 243516 159456 243568
rect 159508 243556 159514 243568
rect 171778 243556 171784 243568
rect 159508 243528 171784 243556
rect 159508 243516 159514 243528
rect 171778 243516 171784 243528
rect 171836 243516 171842 243568
rect 128354 242904 128360 242956
rect 128412 242944 128418 242956
rect 129642 242944 129648 242956
rect 128412 242916 129648 242944
rect 128412 242904 128418 242916
rect 129642 242904 129648 242916
rect 129700 242944 129706 242956
rect 162118 242944 162124 242956
rect 129700 242916 162124 242944
rect 129700 242904 129706 242916
rect 162118 242904 162124 242916
rect 162176 242904 162182 242956
rect 296254 242904 296260 242956
rect 296312 242944 296318 242956
rect 300946 242944 300952 242956
rect 296312 242916 300952 242944
rect 296312 242904 296318 242916
rect 300946 242904 300952 242916
rect 301004 242904 301010 242956
rect 318150 242904 318156 242956
rect 318208 242944 318214 242956
rect 357526 242944 357532 242956
rect 318208 242916 357532 242944
rect 318208 242904 318214 242916
rect 357526 242904 357532 242916
rect 357584 242944 357590 242956
rect 358814 242944 358820 242956
rect 357584 242916 358820 242944
rect 357584 242904 357590 242916
rect 358814 242904 358820 242916
rect 358872 242904 358878 242956
rect 442166 242904 442172 242956
rect 442224 242944 442230 242956
rect 443270 242944 443276 242956
rect 442224 242916 443276 242944
rect 442224 242904 442230 242916
rect 443270 242904 443276 242916
rect 443328 242904 443334 242956
rect 121454 242836 121460 242888
rect 121512 242876 121518 242888
rect 138842 242876 138848 242888
rect 121512 242848 138848 242876
rect 121512 242836 121518 242848
rect 138842 242836 138848 242848
rect 138900 242836 138906 242888
rect 121546 242768 121552 242820
rect 121604 242808 121610 242820
rect 128354 242808 128360 242820
rect 121604 242780 128360 242808
rect 121604 242768 121610 242780
rect 128354 242768 128360 242780
rect 128412 242768 128418 242820
rect 142982 242292 142988 242344
rect 143040 242332 143046 242344
rect 174998 242332 175004 242344
rect 143040 242304 175004 242332
rect 143040 242292 143046 242304
rect 174998 242292 175004 242304
rect 175056 242292 175062 242344
rect 145650 242224 145656 242276
rect 145708 242264 145714 242276
rect 179874 242264 179880 242276
rect 145708 242236 179880 242264
rect 145708 242224 145714 242236
rect 179874 242224 179880 242236
rect 179932 242224 179938 242276
rect 63402 242156 63408 242208
rect 63460 242196 63466 242208
rect 69658 242196 69664 242208
rect 63460 242168 69664 242196
rect 63460 242156 63466 242168
rect 69658 242156 69664 242168
rect 69716 242156 69722 242208
rect 119982 242156 119988 242208
rect 120040 242196 120046 242208
rect 170490 242196 170496 242208
rect 120040 242168 170496 242196
rect 120040 242156 120046 242168
rect 170490 242156 170496 242168
rect 170548 242156 170554 242208
rect 442902 242156 442908 242208
rect 442960 242196 442966 242208
rect 444466 242196 444472 242208
rect 442960 242168 444472 242196
rect 442960 242156 442966 242168
rect 444466 242156 444472 242168
rect 444524 242156 444530 242208
rect 63310 241544 63316 241596
rect 63368 241584 63374 241596
rect 67634 241584 67640 241596
rect 63368 241556 67640 241584
rect 63368 241544 63374 241556
rect 67634 241544 67640 241556
rect 67692 241544 67698 241596
rect 61746 241476 61752 241528
rect 61804 241516 61810 241528
rect 67726 241516 67732 241528
rect 61804 241488 67732 241516
rect 61804 241476 61810 241488
rect 67726 241476 67732 241488
rect 67784 241476 67790 241528
rect 174998 241476 175004 241528
rect 175056 241516 175062 241528
rect 176654 241516 176660 241528
rect 175056 241488 176660 241516
rect 175056 241476 175062 241488
rect 176654 241476 176660 241488
rect 176712 241476 176718 241528
rect 53558 241408 53564 241460
rect 53616 241448 53622 241460
rect 67634 241448 67640 241460
rect 53616 241420 67640 241448
rect 53616 241408 53622 241420
rect 67634 241408 67640 241420
rect 67692 241408 67698 241460
rect 296438 241408 296444 241460
rect 296496 241448 296502 241460
rect 296622 241448 296628 241460
rect 296496 241420 296628 241448
rect 296496 241408 296502 241420
rect 296622 241408 296628 241420
rect 296680 241448 296686 241460
rect 300210 241448 300216 241460
rect 296680 241420 300216 241448
rect 296680 241408 296686 241420
rect 300210 241408 300216 241420
rect 300268 241408 300274 241460
rect 150066 240864 150072 240916
rect 150124 240904 150130 240916
rect 150124 240876 184244 240904
rect 150124 240864 150130 240876
rect 155770 240796 155776 240848
rect 155828 240836 155834 240848
rect 155828 240808 180794 240836
rect 155828 240796 155834 240808
rect 42702 240728 42708 240780
rect 42760 240768 42766 240780
rect 67634 240768 67640 240780
rect 42760 240740 67640 240768
rect 42760 240728 42766 240740
rect 67634 240728 67640 240740
rect 67692 240728 67698 240780
rect 127618 240728 127624 240780
rect 127676 240768 127682 240780
rect 179506 240768 179512 240780
rect 127676 240740 179512 240768
rect 127676 240728 127682 240740
rect 179506 240728 179512 240740
rect 179564 240728 179570 240780
rect 180766 240496 180794 240808
rect 184216 240644 184244 240876
rect 306374 240836 306380 240848
rect 287026 240808 306380 240836
rect 184198 240592 184204 240644
rect 184256 240592 184262 240644
rect 284202 240592 284208 240644
rect 284260 240632 284266 240644
rect 287026 240632 287054 240808
rect 306374 240796 306380 240808
rect 306432 240796 306438 240848
rect 372522 240796 372528 240848
rect 372580 240836 372586 240848
rect 372580 240808 377812 240836
rect 372580 240796 372586 240808
rect 301130 240728 301136 240780
rect 301188 240768 301194 240780
rect 301682 240768 301688 240780
rect 301188 240740 301688 240768
rect 301188 240728 301194 240740
rect 301682 240728 301688 240740
rect 301740 240768 301746 240780
rect 301740 240740 373994 240768
rect 301740 240728 301746 240740
rect 284260 240604 287054 240632
rect 373966 240632 373994 240740
rect 377784 240700 377812 240808
rect 476114 240768 476120 240780
rect 383626 240740 476120 240768
rect 381538 240700 381544 240712
rect 377784 240672 381544 240700
rect 381538 240660 381544 240672
rect 381596 240660 381602 240712
rect 383626 240632 383654 240740
rect 476114 240728 476120 240740
rect 476172 240728 476178 240780
rect 373966 240604 383654 240632
rect 284260 240592 284266 240604
rect 191926 240496 191932 240508
rect 180766 240468 191932 240496
rect 191926 240456 191932 240468
rect 191984 240456 191990 240508
rect 121454 240116 121460 240168
rect 121512 240156 121518 240168
rect 149882 240156 149888 240168
rect 121512 240128 149888 240156
rect 121512 240116 121518 240128
rect 149882 240116 149888 240128
rect 149940 240116 149946 240168
rect 3418 240048 3424 240100
rect 3476 240088 3482 240100
rect 48222 240088 48228 240100
rect 3476 240060 48228 240088
rect 3476 240048 3482 240060
rect 48222 240048 48228 240060
rect 48280 240048 48286 240100
rect 148502 240048 148508 240100
rect 148560 240088 148566 240100
rect 301130 240088 301136 240100
rect 148560 240060 301136 240088
rect 148560 240048 148566 240060
rect 301130 240048 301136 240060
rect 301188 240048 301194 240100
rect 310422 240048 310428 240100
rect 310480 240088 310486 240100
rect 310606 240088 310612 240100
rect 310480 240060 310612 240088
rect 310480 240048 310486 240060
rect 310606 240048 310612 240060
rect 310664 240048 310670 240100
rect 439498 239640 439504 239692
rect 439556 239680 439562 239692
rect 444558 239680 444564 239692
rect 439556 239652 444564 239680
rect 439556 239640 439562 239652
rect 444558 239640 444564 239652
rect 444616 239640 444622 239692
rect 395982 239504 395988 239556
rect 396040 239544 396046 239556
rect 440418 239544 440424 239556
rect 396040 239516 440424 239544
rect 396040 239504 396046 239516
rect 440418 239504 440424 239516
rect 440476 239504 440482 239556
rect 117130 239436 117136 239488
rect 117188 239476 117194 239488
rect 134610 239476 134616 239488
rect 117188 239448 134616 239476
rect 117188 239436 117194 239448
rect 134610 239436 134616 239448
rect 134668 239436 134674 239488
rect 158622 239436 158628 239488
rect 158680 239476 158686 239488
rect 220170 239476 220176 239488
rect 158680 239448 220176 239476
rect 158680 239436 158686 239448
rect 220170 239436 220176 239448
rect 220228 239436 220234 239488
rect 382182 239436 382188 239488
rect 382240 239476 382246 239488
rect 441706 239476 441712 239488
rect 382240 239448 441712 239476
rect 382240 239436 382246 239448
rect 441706 239436 441712 239448
rect 441764 239436 441770 239488
rect 48222 239368 48228 239420
rect 48280 239408 48286 239420
rect 71682 239408 71688 239420
rect 48280 239380 71688 239408
rect 48280 239368 48286 239380
rect 71682 239368 71688 239380
rect 71740 239368 71746 239420
rect 116762 239368 116768 239420
rect 116820 239408 116826 239420
rect 136726 239408 136732 239420
rect 116820 239380 136732 239408
rect 116820 239368 116826 239380
rect 136726 239368 136732 239380
rect 136784 239368 136790 239420
rect 161290 239368 161296 239420
rect 161348 239408 161354 239420
rect 323394 239408 323400 239420
rect 161348 239380 323400 239408
rect 161348 239368 161354 239380
rect 323394 239368 323400 239380
rect 323452 239368 323458 239420
rect 382090 239368 382096 239420
rect 382148 239408 382154 239420
rect 441614 239408 441620 239420
rect 382148 239380 441620 239408
rect 382148 239368 382154 239380
rect 441614 239368 441620 239380
rect 441672 239368 441678 239420
rect 443730 239368 443736 239420
rect 443788 239408 443794 239420
rect 580258 239408 580264 239420
rect 443788 239380 580264 239408
rect 443788 239368 443794 239380
rect 580258 239368 580264 239380
rect 580316 239368 580322 239420
rect 189074 239096 189080 239148
rect 189132 239136 189138 239148
rect 190178 239136 190184 239148
rect 189132 239108 190184 239136
rect 189132 239096 189138 239108
rect 190178 239096 190184 239108
rect 190236 239136 190242 239148
rect 382182 239136 382188 239148
rect 190236 239108 382188 239136
rect 190236 239096 190242 239108
rect 382182 239096 382188 239108
rect 382240 239096 382246 239148
rect 64690 239028 64696 239080
rect 64748 239068 64754 239080
rect 70026 239068 70032 239080
rect 64748 239040 70032 239068
rect 64748 239028 64754 239040
rect 70026 239028 70032 239040
rect 70084 239028 70090 239080
rect 316126 239028 316132 239080
rect 316184 239068 316190 239080
rect 317322 239068 317328 239080
rect 316184 239040 317328 239068
rect 316184 239028 316190 239040
rect 317322 239028 317328 239040
rect 317380 239068 317386 239080
rect 390462 239068 390468 239080
rect 317380 239040 390468 239068
rect 317380 239028 317386 239040
rect 390462 239028 390468 239040
rect 390520 239028 390526 239080
rect 60458 238960 60464 239012
rect 60516 239000 60522 239012
rect 80330 239000 80336 239012
rect 60516 238972 80336 239000
rect 60516 238960 60522 238972
rect 80330 238960 80336 238972
rect 80388 238960 80394 239012
rect 119982 238960 119988 239012
rect 120040 239000 120046 239012
rect 125042 239000 125048 239012
rect 120040 238972 125048 239000
rect 120040 238960 120046 238972
rect 125042 238960 125048 238972
rect 125100 238960 125106 239012
rect 263042 238960 263048 239012
rect 263100 239000 263106 239012
rect 297542 239000 297548 239012
rect 263100 238972 297548 239000
rect 263100 238960 263106 238972
rect 297542 238960 297548 238972
rect 297600 238960 297606 239012
rect 376018 238960 376024 239012
rect 376076 239000 376082 239012
rect 435358 239000 435364 239012
rect 376076 238972 435364 239000
rect 376076 238960 376082 238972
rect 435358 238960 435364 238972
rect 435416 239000 435422 239012
rect 438578 239000 438584 239012
rect 435416 238972 438584 239000
rect 435416 238960 435422 238972
rect 438578 238960 438584 238972
rect 438636 238960 438642 239012
rect 59262 238892 59268 238944
rect 59320 238932 59326 238944
rect 91278 238932 91284 238944
rect 59320 238904 91284 238932
rect 59320 238892 59326 238904
rect 91278 238892 91284 238904
rect 91336 238892 91342 238944
rect 117222 238892 117228 238944
rect 117280 238932 117286 238944
rect 210510 238932 210516 238944
rect 117280 238904 210516 238932
rect 117280 238892 117286 238904
rect 210510 238892 210516 238904
rect 210568 238892 210574 238944
rect 219434 238892 219440 238944
rect 219492 238932 219498 238944
rect 382090 238932 382096 238944
rect 219492 238904 382096 238932
rect 219492 238892 219498 238904
rect 382090 238892 382096 238904
rect 382148 238892 382154 238944
rect 390462 238892 390468 238944
rect 390520 238932 390526 238944
rect 438854 238932 438860 238944
rect 390520 238904 438860 238932
rect 390520 238892 390526 238904
rect 438854 238892 438860 238904
rect 438912 238892 438918 238944
rect 48958 238824 48964 238876
rect 49016 238864 49022 238876
rect 85574 238864 85580 238876
rect 49016 238836 85580 238864
rect 49016 238824 49022 238836
rect 85574 238824 85580 238836
rect 85632 238824 85638 238876
rect 99006 238824 99012 238876
rect 99064 238864 99070 238876
rect 120810 238864 120816 238876
rect 99064 238836 120816 238864
rect 99064 238824 99070 238836
rect 120810 238824 120816 238836
rect 120868 238824 120874 238876
rect 173342 238824 173348 238876
rect 173400 238864 173406 238876
rect 215294 238864 215300 238876
rect 173400 238836 215300 238864
rect 173400 238824 173406 238836
rect 215294 238824 215300 238836
rect 215352 238824 215358 238876
rect 269206 238824 269212 238876
rect 269264 238864 269270 238876
rect 395982 238864 395988 238876
rect 269264 238836 395988 238864
rect 269264 238824 269270 238836
rect 395982 238824 395988 238836
rect 396040 238824 396046 238876
rect 37090 238756 37096 238808
rect 37148 238796 37154 238808
rect 81618 238796 81624 238808
rect 37148 238768 81624 238796
rect 37148 238756 37154 238768
rect 81618 238756 81624 238768
rect 81676 238756 81682 238808
rect 91922 238756 91928 238808
rect 91980 238796 91986 238808
rect 144178 238796 144184 238808
rect 91980 238768 144184 238796
rect 91980 238756 91986 238768
rect 144178 238756 144184 238768
rect 144236 238756 144242 238808
rect 179506 238756 179512 238808
rect 179564 238796 179570 238808
rect 189074 238796 189080 238808
rect 179564 238768 189080 238796
rect 179564 238756 179570 238768
rect 189074 238756 189080 238768
rect 189132 238756 189138 238808
rect 223758 238756 223764 238808
rect 223816 238796 223822 238808
rect 269114 238796 269120 238808
rect 223816 238768 269120 238796
rect 223816 238756 223822 238768
rect 269114 238756 269120 238768
rect 269172 238756 269178 238808
rect 379606 238756 379612 238808
rect 379664 238796 379670 238808
rect 398926 238796 398932 238808
rect 379664 238768 398932 238796
rect 379664 238756 379670 238768
rect 398926 238756 398932 238768
rect 398984 238796 398990 238808
rect 399938 238796 399944 238808
rect 398984 238768 399944 238796
rect 398984 238756 398990 238768
rect 399938 238756 399944 238768
rect 399996 238756 400002 238808
rect 436738 238756 436744 238808
rect 436796 238796 436802 238808
rect 443086 238796 443092 238808
rect 436796 238768 443092 238796
rect 436796 238756 436802 238768
rect 443086 238756 443092 238768
rect 443144 238756 443150 238808
rect 3326 238688 3332 238740
rect 3384 238728 3390 238740
rect 55030 238728 55036 238740
rect 3384 238700 55036 238728
rect 3384 238688 3390 238700
rect 55030 238688 55036 238700
rect 55088 238728 55094 238740
rect 103514 238728 103520 238740
rect 55088 238700 103520 238728
rect 55088 238688 55094 238700
rect 103514 238688 103520 238700
rect 103572 238688 103578 238740
rect 114462 238688 114468 238740
rect 114520 238728 114526 238740
rect 117130 238728 117136 238740
rect 114520 238700 117136 238728
rect 114520 238688 114526 238700
rect 117130 238688 117136 238700
rect 117188 238688 117194 238740
rect 118970 238688 118976 238740
rect 119028 238728 119034 238740
rect 131850 238728 131856 238740
rect 119028 238700 131856 238728
rect 119028 238688 119034 238700
rect 131850 238688 131856 238700
rect 131908 238688 131914 238740
rect 178678 238688 178684 238740
rect 178736 238728 178742 238740
rect 196434 238728 196440 238740
rect 178736 238700 196440 238728
rect 178736 238688 178742 238700
rect 196434 238688 196440 238700
rect 196492 238688 196498 238740
rect 204806 238688 204812 238740
rect 204864 238728 204870 238740
rect 376570 238728 376576 238740
rect 204864 238700 376576 238728
rect 204864 238688 204870 238700
rect 376570 238688 376576 238700
rect 376628 238728 376634 238740
rect 424318 238728 424324 238740
rect 376628 238700 424324 238728
rect 376628 238688 376634 238700
rect 424318 238688 424324 238700
rect 424376 238688 424382 238740
rect 438578 238688 438584 238740
rect 438636 238728 438642 238740
rect 443730 238728 443736 238740
rect 438636 238700 443736 238728
rect 438636 238688 438642 238700
rect 443730 238688 443736 238700
rect 443788 238688 443794 238740
rect 71682 238620 71688 238672
rect 71740 238660 71746 238672
rect 112530 238660 112536 238672
rect 71740 238632 112536 238660
rect 71740 238620 71746 238632
rect 112530 238620 112536 238632
rect 112588 238660 112594 238672
rect 117222 238660 117228 238672
rect 112588 238632 117228 238660
rect 112588 238620 112594 238632
rect 117222 238620 117228 238632
rect 117280 238620 117286 238672
rect 117682 238620 117688 238672
rect 117740 238660 117746 238672
rect 250530 238660 250536 238672
rect 117740 238632 250536 238660
rect 117740 238620 117746 238632
rect 250530 238620 250536 238632
rect 250588 238620 250594 238672
rect 264974 238620 264980 238672
rect 265032 238660 265038 238672
rect 279418 238660 279424 238672
rect 265032 238632 279424 238660
rect 265032 238620 265038 238632
rect 279418 238620 279424 238632
rect 279476 238620 279482 238672
rect 296530 238620 296536 238672
rect 296588 238660 296594 238672
rect 387242 238660 387248 238672
rect 296588 238632 387248 238660
rect 296588 238620 296594 238632
rect 387242 238620 387248 238632
rect 387300 238620 387306 238672
rect 420178 238620 420184 238672
rect 420236 238660 420242 238672
rect 458266 238660 458272 238672
rect 420236 238632 458272 238660
rect 420236 238620 420242 238632
rect 458266 238620 458272 238632
rect 458324 238620 458330 238672
rect 57882 238552 57888 238604
rect 57940 238592 57946 238604
rect 74534 238592 74540 238604
rect 57940 238564 74540 238592
rect 57940 238552 57946 238564
rect 74534 238552 74540 238564
rect 74592 238552 74598 238604
rect 85574 238552 85580 238604
rect 85632 238592 85638 238604
rect 86770 238592 86776 238604
rect 85632 238564 86776 238592
rect 85632 238552 85638 238564
rect 86770 238552 86776 238564
rect 86828 238552 86834 238604
rect 117038 238552 117044 238604
rect 117096 238592 117102 238604
rect 123662 238592 123668 238604
rect 117096 238564 123668 238592
rect 117096 238552 117102 238564
rect 123662 238552 123668 238564
rect 123720 238552 123726 238604
rect 219342 238552 219348 238604
rect 219400 238592 219406 238604
rect 341518 238592 341524 238604
rect 219400 238564 341524 238592
rect 219400 238552 219406 238564
rect 341518 238552 341524 238564
rect 341576 238592 341582 238604
rect 407758 238592 407764 238604
rect 341576 238564 407764 238592
rect 341576 238552 341582 238564
rect 407758 238552 407764 238564
rect 407816 238552 407822 238604
rect 50890 238484 50896 238536
rect 50948 238524 50954 238536
rect 73246 238524 73252 238536
rect 50948 238496 73252 238524
rect 50948 238484 50954 238496
rect 73246 238484 73252 238496
rect 73304 238484 73310 238536
rect 118326 238484 118332 238536
rect 118384 238524 118390 238536
rect 240134 238524 240140 238536
rect 118384 238496 240140 238524
rect 118384 238484 118390 238496
rect 240134 238484 240140 238496
rect 240192 238484 240198 238536
rect 307202 238524 307208 238536
rect 302206 238496 307208 238524
rect 75822 238416 75828 238468
rect 75880 238456 75886 238468
rect 80882 238456 80888 238468
rect 75880 238428 80888 238456
rect 75880 238416 75886 238428
rect 80882 238416 80888 238428
rect 80940 238416 80946 238468
rect 115106 238416 115112 238468
rect 115164 238456 115170 238468
rect 236362 238456 236368 238468
rect 115164 238428 236368 238456
rect 115164 238416 115170 238428
rect 236362 238416 236368 238428
rect 236420 238456 236426 238468
rect 296530 238456 296536 238468
rect 236420 238428 296536 238456
rect 236420 238416 236426 238428
rect 296530 238416 296536 238428
rect 296588 238416 296594 238468
rect 108022 238348 108028 238400
rect 108080 238388 108086 238400
rect 119982 238388 119988 238400
rect 108080 238360 119988 238388
rect 108080 238348 108086 238360
rect 119982 238348 119988 238360
rect 120040 238348 120046 238400
rect 196434 238348 196440 238400
rect 196492 238388 196498 238400
rect 219434 238388 219440 238400
rect 196492 238360 219440 238388
rect 196492 238348 196498 238360
rect 219434 238348 219440 238360
rect 219492 238348 219498 238400
rect 253198 238348 253204 238400
rect 253256 238388 253262 238400
rect 302206 238388 302234 238496
rect 307202 238484 307208 238496
rect 307260 238524 307266 238536
rect 393590 238524 393596 238536
rect 307260 238496 393596 238524
rect 307260 238484 307266 238496
rect 393590 238484 393596 238496
rect 393648 238484 393654 238536
rect 312630 238416 312636 238468
rect 312688 238456 312694 238468
rect 384298 238456 384304 238468
rect 312688 238428 384304 238456
rect 312688 238416 312694 238428
rect 384298 238416 384304 238428
rect 384356 238416 384362 238468
rect 253256 238360 302234 238388
rect 253256 238348 253262 238360
rect 240134 238280 240140 238332
rect 240192 238320 240198 238332
rect 315298 238320 315304 238332
rect 240192 238292 315304 238320
rect 240192 238280 240198 238292
rect 315298 238280 315304 238292
rect 315356 238280 315362 238332
rect 46658 238008 46664 238060
rect 46716 238048 46722 238060
rect 77202 238048 77208 238060
rect 46716 238020 77208 238048
rect 46716 238008 46722 238020
rect 77202 238008 77208 238020
rect 77260 238008 77266 238060
rect 86770 238008 86776 238060
rect 86828 238048 86834 238060
rect 208486 238048 208492 238060
rect 86828 238020 208492 238048
rect 86828 238008 86834 238020
rect 208486 238008 208492 238020
rect 208544 238008 208550 238060
rect 257614 238008 257620 238060
rect 257672 238048 257678 238060
rect 262122 238048 262128 238060
rect 257672 238020 262128 238048
rect 257672 238008 257678 238020
rect 262122 238008 262128 238020
rect 262180 238008 262186 238060
rect 291194 238008 291200 238060
rect 291252 238048 291258 238060
rect 312630 238048 312636 238060
rect 291252 238020 312636 238048
rect 291252 238008 291258 238020
rect 312630 238008 312636 238020
rect 312688 238008 312694 238060
rect 315298 238008 315304 238060
rect 315356 238048 315362 238060
rect 405642 238048 405648 238060
rect 315356 238020 405648 238048
rect 315356 238008 315362 238020
rect 405642 238008 405648 238020
rect 405700 238008 405706 238060
rect 432230 238008 432236 238060
rect 432288 238048 432294 238060
rect 454034 238048 454040 238060
rect 432288 238020 454040 238048
rect 432288 238008 432294 238020
rect 454034 238008 454040 238020
rect 454092 238048 454098 238060
rect 456886 238048 456892 238060
rect 454092 238020 456892 238048
rect 454092 238008 454098 238020
rect 456886 238008 456892 238020
rect 456944 238008 456950 238060
rect 77202 237804 77208 237856
rect 77260 237844 77266 237856
rect 77754 237844 77760 237856
rect 77260 237816 77760 237844
rect 77260 237804 77266 237816
rect 77754 237804 77760 237816
rect 77812 237804 77818 237856
rect 422294 237668 422300 237720
rect 422352 237708 422358 237720
rect 426342 237708 426348 237720
rect 422352 237680 426348 237708
rect 422352 237668 422358 237680
rect 426342 237668 426348 237680
rect 426400 237668 426406 237720
rect 74534 237396 74540 237448
rect 74592 237436 74598 237448
rect 75178 237436 75184 237448
rect 74592 237408 75184 237436
rect 74592 237396 74598 237408
rect 75178 237396 75184 237408
rect 75236 237396 75242 237448
rect 79042 237396 79048 237448
rect 79100 237436 79106 237448
rect 80790 237436 80796 237448
rect 79100 237408 80796 237436
rect 79100 237396 79106 237408
rect 80790 237396 80796 237408
rect 80848 237396 80854 237448
rect 82078 237396 82084 237448
rect 82136 237436 82142 237448
rect 82906 237436 82912 237448
rect 82136 237408 82912 237436
rect 82136 237396 82142 237408
rect 82906 237396 82912 237408
rect 82964 237396 82970 237448
rect 208486 237396 208492 237448
rect 208544 237436 208550 237448
rect 209682 237436 209688 237448
rect 208544 237408 209688 237436
rect 208544 237396 208550 237408
rect 209682 237396 209688 237408
rect 209740 237436 209746 237448
rect 210602 237436 210608 237448
rect 209740 237408 210608 237436
rect 209740 237396 209746 237408
rect 210602 237396 210608 237408
rect 210660 237396 210666 237448
rect 432690 237396 432696 237448
rect 432748 237436 432754 237448
rect 434070 237436 434076 237448
rect 432748 237408 434076 237436
rect 432748 237396 432754 237408
rect 434070 237396 434076 237408
rect 434128 237396 434134 237448
rect 46750 237328 46756 237380
rect 46808 237368 46814 237380
rect 82096 237368 82124 237396
rect 46808 237340 82124 237368
rect 46808 237328 46814 237340
rect 107378 237328 107384 237380
rect 107436 237368 107442 237380
rect 116762 237368 116768 237380
rect 107436 237340 116768 237368
rect 107436 237328 107442 237340
rect 116762 237328 116768 237340
rect 116820 237328 116826 237380
rect 172330 237328 172336 237380
rect 172388 237368 172394 237380
rect 458358 237368 458364 237380
rect 172388 237340 458364 237368
rect 172388 237328 172394 237340
rect 458358 237328 458364 237340
rect 458416 237328 458422 237380
rect 54754 237260 54760 237312
rect 54812 237300 54818 237312
rect 325694 237300 325700 237312
rect 54812 237272 325700 237300
rect 54812 237260 54818 237272
rect 325694 237260 325700 237272
rect 325752 237300 325758 237312
rect 326338 237300 326344 237312
rect 325752 237272 326344 237300
rect 325752 237260 325758 237272
rect 326338 237260 326344 237272
rect 326396 237260 326402 237312
rect 357342 237260 357348 237312
rect 357400 237300 357406 237312
rect 411898 237300 411904 237312
rect 357400 237272 411904 237300
rect 357400 237260 357406 237272
rect 411898 237260 411904 237272
rect 411956 237260 411962 237312
rect 54938 237192 54944 237244
rect 54996 237232 55002 237244
rect 89346 237232 89352 237244
rect 54996 237204 89352 237232
rect 54996 237192 55002 237204
rect 89346 237192 89352 237204
rect 89404 237192 89410 237244
rect 106734 237192 106740 237244
rect 106792 237232 106798 237244
rect 140590 237232 140596 237244
rect 106792 237204 140596 237232
rect 106792 237192 106798 237204
rect 140590 237192 140596 237204
rect 140648 237192 140654 237244
rect 156690 237192 156696 237244
rect 156748 237232 156754 237244
rect 276014 237232 276020 237244
rect 156748 237204 276020 237232
rect 156748 237192 156754 237204
rect 276014 237192 276020 237204
rect 276072 237192 276078 237244
rect 288250 237192 288256 237244
rect 288308 237232 288314 237244
rect 313366 237232 313372 237244
rect 288308 237204 313372 237232
rect 288308 237192 288314 237204
rect 313366 237192 313372 237204
rect 313424 237192 313430 237244
rect 325142 237192 325148 237244
rect 325200 237232 325206 237244
rect 422294 237232 422300 237244
rect 325200 237204 422300 237232
rect 325200 237192 325206 237204
rect 422294 237192 422300 237204
rect 422352 237192 422358 237244
rect 45462 237124 45468 237176
rect 45520 237164 45526 237176
rect 77110 237164 77116 237176
rect 45520 237136 77116 237164
rect 45520 237124 45526 237136
rect 77110 237124 77116 237136
rect 77168 237124 77174 237176
rect 88702 237124 88708 237176
rect 88760 237164 88766 237176
rect 120718 237164 120724 237176
rect 88760 237136 120724 237164
rect 88760 237124 88766 237136
rect 120718 237124 120724 237136
rect 120776 237124 120782 237176
rect 179874 237124 179880 237176
rect 179932 237164 179938 237176
rect 204806 237164 204812 237176
rect 179932 237136 204812 237164
rect 179932 237124 179938 237136
rect 204806 237124 204812 237136
rect 204864 237124 204870 237176
rect 284662 237124 284668 237176
rect 284720 237164 284726 237176
rect 285582 237164 285588 237176
rect 284720 237136 285588 237164
rect 284720 237124 284726 237136
rect 285582 237124 285588 237136
rect 285640 237164 285646 237176
rect 308490 237164 308496 237176
rect 285640 237136 308496 237164
rect 285640 237124 285646 237136
rect 308490 237124 308496 237136
rect 308548 237124 308554 237176
rect 375098 237124 375104 237176
rect 375156 237164 375162 237176
rect 402974 237164 402980 237176
rect 375156 237136 402980 237164
rect 375156 237124 375162 237136
rect 402974 237124 402980 237136
rect 403032 237164 403038 237176
rect 403802 237164 403808 237176
rect 403032 237136 403808 237164
rect 403032 237124 403038 237136
rect 403802 237124 403808 237136
rect 403860 237124 403866 237176
rect 115842 237056 115848 237108
rect 115900 237096 115906 237108
rect 133322 237096 133328 237108
rect 115900 237068 133328 237096
rect 115900 237056 115906 237068
rect 133322 237056 133328 237068
rect 133380 237056 133386 237108
rect 86126 236988 86132 237040
rect 86184 237028 86190 237040
rect 130470 237028 130476 237040
rect 86184 237000 130476 237028
rect 86184 236988 86190 237000
rect 130470 236988 130476 237000
rect 130528 236988 130534 237040
rect 429102 236920 429108 236972
rect 429160 236960 429166 236972
rect 440234 236960 440240 236972
rect 429160 236932 440240 236960
rect 429160 236920 429166 236932
rect 440234 236920 440240 236932
rect 440292 236920 440298 236972
rect 443178 236920 443184 236972
rect 443236 236960 443242 236972
rect 459738 236960 459744 236972
rect 443236 236932 459744 236960
rect 443236 236920 443242 236932
rect 459738 236920 459744 236932
rect 459796 236920 459802 236972
rect 426434 236852 426440 236904
rect 426492 236892 426498 236904
rect 451274 236892 451280 236904
rect 426492 236864 451280 236892
rect 426492 236852 426498 236864
rect 451274 236852 451280 236864
rect 451332 236852 451338 236904
rect 414014 236784 414020 236836
rect 414072 236824 414078 236836
rect 449986 236824 449992 236836
rect 414072 236796 449992 236824
rect 414072 236784 414078 236796
rect 449986 236784 449992 236796
rect 450044 236784 450050 236836
rect 163682 236716 163688 236768
rect 163740 236756 163746 236768
rect 193950 236756 193956 236768
rect 163740 236728 193956 236756
rect 163740 236716 163746 236728
rect 193950 236716 193956 236728
rect 194008 236716 194014 236768
rect 261478 236716 261484 236768
rect 261536 236756 261542 236768
rect 291838 236756 291844 236768
rect 261536 236728 291844 236756
rect 261536 236716 261542 236728
rect 291838 236716 291844 236728
rect 291896 236716 291902 236768
rect 394602 236716 394608 236768
rect 394660 236756 394666 236768
rect 452838 236756 452844 236768
rect 394660 236728 452844 236756
rect 394660 236716 394666 236728
rect 452838 236716 452844 236728
rect 452896 236716 452902 236768
rect 140590 236648 140596 236700
rect 140648 236688 140654 236700
rect 288526 236688 288532 236700
rect 140648 236660 288532 236688
rect 140648 236648 140654 236660
rect 288526 236648 288532 236660
rect 288584 236648 288590 236700
rect 378042 236648 378048 236700
rect 378100 236688 378106 236700
rect 392578 236688 392584 236700
rect 378100 236660 392584 236688
rect 378100 236648 378106 236660
rect 392578 236648 392584 236660
rect 392636 236648 392642 236700
rect 432598 236648 432604 236700
rect 432656 236688 432662 236700
rect 561674 236688 561680 236700
rect 432656 236660 561680 236688
rect 432656 236648 432662 236660
rect 561674 236648 561680 236660
rect 561732 236648 561738 236700
rect 76558 235968 76564 236020
rect 76616 236008 76622 236020
rect 77110 236008 77116 236020
rect 76616 235980 77116 236008
rect 76616 235968 76622 235980
rect 77110 235968 77116 235980
rect 77168 235968 77174 236020
rect 393590 235968 393596 236020
rect 393648 236008 393654 236020
rect 395338 236008 395344 236020
rect 393648 235980 395344 236008
rect 393648 235968 393654 235980
rect 395338 235968 395344 235980
rect 395396 235968 395402 236020
rect 250530 235900 250536 235952
rect 250588 235940 250594 235952
rect 316126 235940 316132 235952
rect 250588 235912 316132 235940
rect 250588 235900 250594 235912
rect 316126 235900 316132 235912
rect 316184 235900 316190 235952
rect 373350 235900 373356 235952
rect 373408 235940 373414 235952
rect 467926 235940 467932 235952
rect 373408 235912 467932 235940
rect 373408 235900 373414 235912
rect 467926 235900 467932 235912
rect 467984 235900 467990 235952
rect 37182 235832 37188 235884
rect 37240 235872 37246 235884
rect 94406 235872 94412 235884
rect 37240 235844 94412 235872
rect 37240 235832 37246 235844
rect 94406 235832 94412 235844
rect 94464 235872 94470 235884
rect 95142 235872 95148 235884
rect 94464 235844 95148 235872
rect 94464 235832 94470 235844
rect 95142 235832 95148 235844
rect 95200 235832 95206 235884
rect 113818 235832 113824 235884
rect 113876 235872 113882 235884
rect 138014 235872 138020 235884
rect 113876 235844 138020 235872
rect 113876 235832 113882 235844
rect 138014 235832 138020 235844
rect 138072 235832 138078 235884
rect 166718 235832 166724 235884
rect 166776 235872 166782 235884
rect 358078 235872 358084 235884
rect 166776 235844 358084 235872
rect 166776 235832 166782 235844
rect 358078 235832 358084 235844
rect 358136 235832 358142 235884
rect 368382 235832 368388 235884
rect 368440 235872 368446 235884
rect 398098 235872 398104 235884
rect 368440 235844 398104 235872
rect 368440 235832 368446 235844
rect 398098 235832 398104 235844
rect 398156 235832 398162 235884
rect 48130 235764 48136 235816
rect 48188 235804 48194 235816
rect 79318 235804 79324 235816
rect 48188 235776 79324 235804
rect 48188 235764 48194 235776
rect 79318 235764 79324 235776
rect 79376 235764 79382 235816
rect 109678 235764 109684 235816
rect 109736 235804 109742 235816
rect 125134 235804 125140 235816
rect 109736 235776 125140 235804
rect 109736 235764 109742 235776
rect 125134 235764 125140 235776
rect 125192 235764 125198 235816
rect 155310 235764 155316 235816
rect 155368 235804 155374 235816
rect 269206 235804 269212 235816
rect 155368 235776 269212 235804
rect 155368 235764 155374 235776
rect 269206 235764 269212 235776
rect 269264 235764 269270 235816
rect 269298 235764 269304 235816
rect 269356 235804 269362 235816
rect 317414 235804 317420 235816
rect 269356 235776 317420 235804
rect 269356 235764 269362 235776
rect 317414 235764 317420 235776
rect 317472 235804 317478 235816
rect 377398 235804 377404 235816
rect 317472 235776 377404 235804
rect 317472 235764 317478 235776
rect 377398 235764 377404 235776
rect 377456 235764 377462 235816
rect 159542 235696 159548 235748
rect 159600 235736 159606 235748
rect 273990 235736 273996 235748
rect 159600 235708 273996 235736
rect 159600 235696 159606 235708
rect 273990 235696 273996 235708
rect 274048 235696 274054 235748
rect 286594 235696 286600 235748
rect 286652 235736 286658 235748
rect 286870 235736 286876 235748
rect 286652 235708 286876 235736
rect 286652 235696 286658 235708
rect 286870 235696 286876 235708
rect 286928 235736 286934 235748
rect 307110 235736 307116 235748
rect 286928 235708 307116 235736
rect 286928 235696 286934 235708
rect 307110 235696 307116 235708
rect 307168 235696 307174 235748
rect 347038 235696 347044 235748
rect 347096 235736 347102 235748
rect 402238 235736 402244 235748
rect 347096 235708 402244 235736
rect 347096 235696 347102 235708
rect 402238 235696 402244 235708
rect 402296 235696 402302 235748
rect 234062 235628 234068 235680
rect 234120 235668 234126 235680
rect 318058 235668 318064 235680
rect 234120 235640 318064 235668
rect 234120 235628 234126 235640
rect 318058 235628 318064 235640
rect 318116 235628 318122 235680
rect 352558 235628 352564 235680
rect 352616 235668 352622 235680
rect 391290 235668 391296 235680
rect 352616 235640 391296 235668
rect 352616 235628 352622 235640
rect 391290 235628 391296 235640
rect 391348 235628 391354 235680
rect 61930 235560 61936 235612
rect 61988 235600 61994 235612
rect 263042 235600 263048 235612
rect 61988 235572 263048 235600
rect 61988 235560 61994 235572
rect 263042 235560 263048 235572
rect 263100 235560 263106 235612
rect 67634 235220 67640 235272
rect 67692 235260 67698 235272
rect 242158 235260 242164 235272
rect 67692 235232 242164 235260
rect 67692 235220 67698 235232
rect 242158 235220 242164 235232
rect 242216 235220 242222 235272
rect 323394 235220 323400 235272
rect 323452 235260 323458 235272
rect 397362 235260 397368 235272
rect 323452 235232 397368 235260
rect 323452 235220 323458 235232
rect 397362 235220 397368 235232
rect 397420 235260 397426 235272
rect 448790 235260 448796 235272
rect 397420 235232 448796 235260
rect 397420 235220 397426 235232
rect 448790 235220 448796 235232
rect 448848 235220 448854 235272
rect 289814 234608 289820 234660
rect 289872 234648 289878 234660
rect 294138 234648 294144 234660
rect 289872 234620 294144 234648
rect 289872 234608 289878 234620
rect 294138 234608 294144 234620
rect 294196 234608 294202 234660
rect 349890 234608 349896 234660
rect 349948 234648 349954 234660
rect 353386 234648 353392 234660
rect 349948 234620 353392 234648
rect 349948 234608 349954 234620
rect 353386 234608 353392 234620
rect 353444 234608 353450 234660
rect 35158 234540 35164 234592
rect 35216 234580 35222 234592
rect 35710 234580 35716 234592
rect 35216 234552 35716 234580
rect 35216 234540 35222 234552
rect 35710 234540 35716 234552
rect 35768 234580 35774 234592
rect 303614 234580 303620 234592
rect 35768 234552 303620 234580
rect 35768 234540 35774 234552
rect 303614 234540 303620 234552
rect 303672 234540 303678 234592
rect 321370 234540 321376 234592
rect 321428 234580 321434 234592
rect 326522 234580 326528 234592
rect 321428 234552 326528 234580
rect 321428 234540 321434 234552
rect 326522 234540 326528 234552
rect 326580 234540 326586 234592
rect 331306 234540 331312 234592
rect 331364 234580 331370 234592
rect 332502 234580 332508 234592
rect 331364 234552 332508 234580
rect 331364 234540 331370 234552
rect 332502 234540 332508 234552
rect 332560 234580 332566 234592
rect 376110 234580 376116 234592
rect 332560 234552 376116 234580
rect 332560 234540 332566 234552
rect 376110 234540 376116 234552
rect 376168 234540 376174 234592
rect 95786 234472 95792 234524
rect 95844 234512 95850 234524
rect 146938 234512 146944 234524
rect 95844 234484 146944 234512
rect 95844 234472 95850 234484
rect 146938 234472 146944 234484
rect 146996 234472 147002 234524
rect 277946 234472 277952 234524
rect 278004 234512 278010 234524
rect 449894 234512 449900 234524
rect 278004 234484 449900 234512
rect 278004 234472 278010 234484
rect 449894 234472 449900 234484
rect 449952 234472 449958 234524
rect 162118 234404 162124 234456
rect 162176 234444 162182 234456
rect 331306 234444 331312 234456
rect 162176 234416 331312 234444
rect 162176 234404 162182 234416
rect 331306 234404 331312 234416
rect 331364 234404 331370 234456
rect 276014 234336 276020 234388
rect 276072 234376 276078 234388
rect 311894 234376 311900 234388
rect 276072 234348 311900 234376
rect 276072 234336 276078 234348
rect 311894 234336 311900 234348
rect 311952 234336 311958 234388
rect 100294 233996 100300 234048
rect 100352 234036 100358 234048
rect 117958 234036 117964 234048
rect 100352 234008 117964 234036
rect 100352 233996 100358 234008
rect 117958 233996 117964 234008
rect 118016 233996 118022 234048
rect 151354 233996 151360 234048
rect 151412 234036 151418 234048
rect 215938 234036 215944 234048
rect 151412 234008 215944 234036
rect 151412 233996 151418 234008
rect 215938 233996 215944 234008
rect 215996 233996 216002 234048
rect 84194 233928 84200 233980
rect 84252 233968 84258 233980
rect 84838 233968 84844 233980
rect 84252 233940 84844 233968
rect 84252 233928 84258 233940
rect 84838 233928 84844 233940
rect 84896 233928 84902 233980
rect 95234 233928 95240 233980
rect 95292 233968 95298 233980
rect 96430 233968 96436 233980
rect 95292 233940 96436 233968
rect 95292 233928 95298 233940
rect 96430 233928 96436 233940
rect 96488 233928 96494 233980
rect 104802 233928 104808 233980
rect 104860 233968 104866 233980
rect 210418 233968 210424 233980
rect 104860 233940 210424 233968
rect 104860 233928 104866 233940
rect 210418 233928 210424 233940
rect 210476 233928 210482 233980
rect 221550 233928 221556 233980
rect 221608 233968 221614 233980
rect 271230 233968 271236 233980
rect 221608 233940 271236 233968
rect 221608 233928 221614 233940
rect 271230 233928 271236 233940
rect 271288 233928 271294 233980
rect 311894 233928 311900 233980
rect 311952 233968 311958 233980
rect 312722 233968 312728 233980
rect 311952 233940 312728 233968
rect 311952 233928 311958 233940
rect 312722 233928 312728 233940
rect 312780 233968 312786 233980
rect 353938 233968 353944 233980
rect 312780 233940 353944 233968
rect 312780 233928 312786 233940
rect 353938 233928 353944 233940
rect 353996 233928 354002 233980
rect 377398 233928 377404 233980
rect 377456 233968 377462 233980
rect 387058 233968 387064 233980
rect 377456 233940 387064 233968
rect 377456 233928 377462 233940
rect 387058 233928 387064 233940
rect 387116 233928 387122 233980
rect 27522 233860 27528 233912
rect 27580 233900 27586 233912
rect 113082 233900 113088 233912
rect 27580 233872 113088 233900
rect 27580 233860 27586 233872
rect 113082 233860 113088 233872
rect 113140 233860 113146 233912
rect 169294 233860 169300 233912
rect 169352 233900 169358 233912
rect 321370 233900 321376 233912
rect 169352 233872 321376 233900
rect 169352 233860 169358 233872
rect 321370 233860 321376 233872
rect 321428 233860 321434 233912
rect 349798 233860 349804 233912
rect 349856 233900 349862 233912
rect 408494 233900 408500 233912
rect 349856 233872 408500 233900
rect 349856 233860 349862 233872
rect 408494 233860 408500 233872
rect 408552 233900 408558 233912
rect 444650 233900 444656 233912
rect 408552 233872 444656 233900
rect 408552 233860 408558 233872
rect 444650 233860 444656 233872
rect 444708 233860 444714 233912
rect 485774 233860 485780 233912
rect 485832 233900 485838 233912
rect 582374 233900 582380 233912
rect 485832 233872 582380 233900
rect 485832 233860 485838 233872
rect 582374 233860 582380 233872
rect 582432 233860 582438 233912
rect 385862 233248 385868 233300
rect 385920 233288 385926 233300
rect 385920 233260 397408 233288
rect 385920 233248 385926 233260
rect 71958 233220 71964 233232
rect 64846 233192 71964 233220
rect 39758 233112 39764 233164
rect 39816 233152 39822 233164
rect 64846 233152 64874 233192
rect 71958 233180 71964 233192
rect 72016 233220 72022 233232
rect 72418 233220 72424 233232
rect 72016 233192 72424 233220
rect 72016 233180 72022 233192
rect 72418 233180 72424 233192
rect 72476 233180 72482 233232
rect 102226 233180 102232 233232
rect 102284 233220 102290 233232
rect 103422 233220 103428 233232
rect 102284 233192 103428 233220
rect 102284 233180 102290 233192
rect 103422 233180 103428 233192
rect 103480 233220 103486 233232
rect 151078 233220 151084 233232
rect 103480 233192 151084 233220
rect 103480 233180 103486 233192
rect 151078 233180 151084 233192
rect 151136 233180 151142 233232
rect 158254 233180 158260 233232
rect 158312 233220 158318 233232
rect 321554 233220 321560 233232
rect 158312 233192 321560 233220
rect 158312 233180 158318 233192
rect 321554 233180 321560 233192
rect 321612 233180 321618 233232
rect 397380 233220 397408 233260
rect 579982 233220 579988 233232
rect 397380 233192 579988 233220
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 39816 233124 64874 233152
rect 39816 233112 39822 233124
rect 76466 233112 76472 233164
rect 76524 233152 76530 233164
rect 135898 233152 135904 233164
rect 76524 233124 135904 233152
rect 76524 233112 76530 233124
rect 135898 233112 135904 233124
rect 135956 233112 135962 233164
rect 152642 233112 152648 233164
rect 152700 233152 152706 233164
rect 299566 233152 299572 233164
rect 152700 233124 299572 233152
rect 152700 233112 152706 233124
rect 299566 233112 299572 233124
rect 299624 233112 299630 233164
rect 337378 233112 337384 233164
rect 337436 233152 337442 233164
rect 431954 233152 431960 233164
rect 337436 233124 431960 233152
rect 337436 233112 337442 233124
rect 431954 233112 431960 233124
rect 432012 233152 432018 233164
rect 432690 233152 432696 233164
rect 432012 233124 432696 233152
rect 432012 233112 432018 233124
rect 432690 233112 432696 233124
rect 432748 233112 432754 233164
rect 52362 233044 52368 233096
rect 52420 233084 52426 233096
rect 80698 233084 80704 233096
rect 52420 233056 80704 233084
rect 52420 233044 52426 233056
rect 80698 233044 80704 233056
rect 80756 233044 80762 233096
rect 98362 233044 98368 233096
rect 98420 233084 98426 233096
rect 234062 233084 234068 233096
rect 98420 233056 234068 233084
rect 98420 233044 98426 233056
rect 234062 233044 234068 233056
rect 234120 233044 234126 233096
rect 271230 233044 271236 233096
rect 271288 233084 271294 233096
rect 304258 233084 304264 233096
rect 271288 233056 304264 233084
rect 271288 233044 271294 233056
rect 304258 233044 304264 233056
rect 304316 233044 304322 233096
rect 382274 233044 382280 233096
rect 382332 233084 382338 233096
rect 450078 233084 450084 233096
rect 382332 233056 450084 233084
rect 382332 233044 382338 233056
rect 450078 233044 450084 233056
rect 450136 233044 450142 233096
rect 83550 232976 83556 233028
rect 83608 233016 83614 233028
rect 126330 233016 126336 233028
rect 83608 232988 126336 233016
rect 83608 232976 83614 232988
rect 126330 232976 126336 232988
rect 126388 232976 126394 233028
rect 129090 232976 129096 233028
rect 129148 233016 129154 233028
rect 223758 233016 223764 233028
rect 129148 232988 223764 233016
rect 129148 232976 129154 232988
rect 223758 232976 223764 232988
rect 223816 232976 223822 233028
rect 356790 232976 356796 233028
rect 356848 233016 356854 233028
rect 410518 233016 410524 233028
rect 356848 232988 410524 233016
rect 356848 232976 356854 232988
rect 410518 232976 410524 232988
rect 410576 232976 410582 233028
rect 32950 232908 32956 232960
rect 33008 232948 33014 232960
rect 104158 232948 104164 232960
rect 33008 232920 104164 232948
rect 33008 232908 33014 232920
rect 104158 232908 104164 232920
rect 104216 232908 104222 232960
rect 381998 232568 382004 232620
rect 382056 232608 382062 232620
rect 388438 232608 388444 232620
rect 382056 232580 388444 232608
rect 382056 232568 382062 232580
rect 388438 232568 388444 232580
rect 388496 232568 388502 232620
rect 369670 232500 369676 232552
rect 369728 232540 369734 232552
rect 387150 232540 387156 232552
rect 369728 232512 387156 232540
rect 369728 232500 369734 232512
rect 387150 232500 387156 232512
rect 387208 232500 387214 232552
rect 450078 232296 450084 232348
rect 450136 232336 450142 232348
rect 450538 232336 450544 232348
rect 450136 232308 450544 232336
rect 450136 232296 450142 232308
rect 450538 232296 450544 232308
rect 450596 232296 450602 232348
rect 110414 232160 110420 232212
rect 110472 232200 110478 232212
rect 111242 232200 111248 232212
rect 110472 232172 111248 232200
rect 110472 232160 110478 232172
rect 111242 232160 111248 232172
rect 111300 232160 111306 232212
rect 61746 231752 61752 231804
rect 61804 231792 61810 231804
rect 264054 231792 264060 231804
rect 61804 231764 264060 231792
rect 61804 231752 61810 231764
rect 264054 231752 264060 231764
rect 264112 231752 264118 231804
rect 314470 231752 314476 231804
rect 314528 231792 314534 231804
rect 314746 231792 314752 231804
rect 314528 231764 314752 231792
rect 314528 231752 314534 231764
rect 314746 231752 314752 231764
rect 314804 231752 314810 231804
rect 31662 231684 31668 231736
rect 31720 231724 31726 231736
rect 106182 231724 106188 231736
rect 31720 231696 106188 231724
rect 31720 231684 31726 231696
rect 106182 231684 106188 231696
rect 106240 231684 106246 231736
rect 166902 231684 166908 231736
rect 166960 231724 166966 231736
rect 198734 231724 198740 231736
rect 166960 231696 198740 231724
rect 166960 231684 166966 231696
rect 198734 231684 198740 231696
rect 198792 231724 198798 231736
rect 199378 231724 199384 231736
rect 198792 231696 199384 231724
rect 198792 231684 198798 231696
rect 199378 231684 199384 231696
rect 199436 231684 199442 231736
rect 214558 231684 214564 231736
rect 214616 231724 214622 231736
rect 362954 231724 362960 231736
rect 214616 231696 362960 231724
rect 214616 231684 214622 231696
rect 362954 231684 362960 231696
rect 363012 231684 363018 231736
rect 93946 231548 93952 231600
rect 94004 231588 94010 231600
rect 94498 231588 94504 231600
rect 94004 231560 94504 231588
rect 94004 231548 94010 231560
rect 94498 231548 94504 231560
rect 94556 231548 94562 231600
rect 278774 231344 278780 231396
rect 278832 231384 278838 231396
rect 294230 231384 294236 231396
rect 278832 231356 294236 231384
rect 278832 231344 278838 231356
rect 294230 231344 294236 231356
rect 294288 231344 294294 231396
rect 167730 231276 167736 231328
rect 167788 231316 167794 231328
rect 279418 231316 279424 231328
rect 167788 231288 279424 231316
rect 167788 231276 167794 231288
rect 279418 231276 279424 231288
rect 279476 231276 279482 231328
rect 106182 231208 106188 231260
rect 106240 231248 106246 231260
rect 243538 231248 243544 231260
rect 106240 231220 243544 231248
rect 106240 231208 106246 231220
rect 243538 231208 243544 231220
rect 243596 231208 243602 231260
rect 248414 231208 248420 231260
rect 248472 231248 248478 231260
rect 282178 231248 282184 231260
rect 248472 231220 282184 231248
rect 248472 231208 248478 231220
rect 282178 231208 282184 231220
rect 282236 231208 282242 231260
rect 296806 231208 296812 231260
rect 296864 231248 296870 231260
rect 301038 231248 301044 231260
rect 296864 231220 301044 231248
rect 296864 231208 296870 231220
rect 301038 231208 301044 231220
rect 301096 231248 301102 231260
rect 391198 231248 391204 231260
rect 301096 231220 391204 231248
rect 301096 231208 301102 231220
rect 391198 231208 391204 231220
rect 391256 231208 391262 231260
rect 141602 231140 141608 231192
rect 141660 231180 141666 231192
rect 314470 231180 314476 231192
rect 141660 231152 314476 231180
rect 141660 231140 141666 231152
rect 314470 231140 314476 231152
rect 314528 231140 314534 231192
rect 78398 231072 78404 231124
rect 78456 231112 78462 231124
rect 126238 231112 126244 231124
rect 78456 231084 126244 231112
rect 78456 231072 78462 231084
rect 126238 231072 126244 231084
rect 126296 231072 126302 231124
rect 158162 231072 158168 231124
rect 158220 231112 158226 231124
rect 220078 231112 220084 231124
rect 158220 231084 220084 231112
rect 158220 231072 158226 231084
rect 220078 231072 220084 231084
rect 220136 231072 220142 231124
rect 220170 231072 220176 231124
rect 220228 231112 220234 231124
rect 426618 231112 426624 231124
rect 220228 231084 426624 231112
rect 220228 231072 220234 231084
rect 426618 231072 426624 231084
rect 426676 231112 426682 231124
rect 451366 231112 451372 231124
rect 426676 231084 451372 231112
rect 426676 231072 426682 231084
rect 451366 231072 451372 231084
rect 451424 231072 451430 231124
rect 289078 231004 289084 231056
rect 289136 231044 289142 231056
rect 295610 231044 295616 231056
rect 289136 231016 295616 231044
rect 289136 231004 289142 231016
rect 295610 231004 295616 231016
rect 295668 231004 295674 231056
rect 59170 230392 59176 230444
rect 59228 230432 59234 230444
rect 288250 230432 288256 230444
rect 59228 230404 288256 230432
rect 59228 230392 59234 230404
rect 288250 230392 288256 230404
rect 288308 230392 288314 230444
rect 297358 230392 297364 230444
rect 297416 230432 297422 230444
rect 365070 230432 365076 230444
rect 297416 230404 365076 230432
rect 297416 230392 297422 230404
rect 365070 230392 365076 230404
rect 365128 230432 365134 230444
rect 396074 230432 396080 230444
rect 365128 230404 396080 230432
rect 365128 230392 365134 230404
rect 396074 230392 396080 230404
rect 396132 230392 396138 230444
rect 143074 230324 143080 230376
rect 143132 230364 143138 230376
rect 300854 230364 300860 230376
rect 143132 230336 300860 230364
rect 143132 230324 143138 230336
rect 300854 230324 300860 230336
rect 300912 230324 300918 230376
rect 184198 230256 184204 230308
rect 184256 230296 184262 230308
rect 310514 230296 310520 230308
rect 184256 230268 310520 230296
rect 184256 230256 184262 230268
rect 310514 230256 310520 230268
rect 310572 230256 310578 230308
rect 396074 229984 396080 230036
rect 396132 230024 396138 230036
rect 396718 230024 396724 230036
rect 396132 229996 396724 230024
rect 396132 229984 396138 229996
rect 396718 229984 396724 229996
rect 396776 229984 396782 230036
rect 171870 229848 171876 229900
rect 171928 229888 171934 229900
rect 189718 229888 189724 229900
rect 171928 229860 189724 229888
rect 171928 229848 171934 229860
rect 189718 229848 189724 229860
rect 189776 229848 189782 229900
rect 371142 229848 371148 229900
rect 371200 229888 371206 229900
rect 458266 229888 458272 229900
rect 371200 229860 458272 229888
rect 371200 229848 371206 229860
rect 458266 229848 458272 229860
rect 458324 229848 458330 229900
rect 64506 229780 64512 229832
rect 64564 229820 64570 229832
rect 98638 229820 98644 229832
rect 64564 229792 98644 229820
rect 64564 229780 64570 229792
rect 98638 229780 98644 229792
rect 98696 229780 98702 229832
rect 131942 229780 131948 229832
rect 132000 229820 132006 229832
rect 203518 229820 203524 229832
rect 132000 229792 203524 229820
rect 132000 229780 132006 229792
rect 203518 229780 203524 229792
rect 203576 229780 203582 229832
rect 244274 229780 244280 229832
rect 244332 229820 244338 229832
rect 266262 229820 266268 229832
rect 244332 229792 266268 229820
rect 244332 229780 244338 229792
rect 266262 229780 266268 229792
rect 266320 229820 266326 229832
rect 305730 229820 305736 229832
rect 266320 229792 305736 229820
rect 266320 229780 266326 229792
rect 305730 229780 305736 229792
rect 305788 229780 305794 229832
rect 386322 229820 386328 229832
rect 373966 229792 386328 229820
rect 3418 229712 3424 229764
rect 3476 229752 3482 229764
rect 120166 229752 120172 229764
rect 3476 229724 120172 229752
rect 3476 229712 3482 229724
rect 120166 229712 120172 229724
rect 120224 229712 120230 229764
rect 165062 229712 165068 229764
rect 165120 229752 165126 229764
rect 261478 229752 261484 229764
rect 165120 229724 261484 229752
rect 165120 229712 165126 229724
rect 261478 229712 261484 229724
rect 261536 229712 261542 229764
rect 281534 229712 281540 229764
rect 281592 229752 281598 229764
rect 373966 229752 373994 229792
rect 386322 229780 386328 229792
rect 386380 229820 386386 229832
rect 489178 229820 489184 229832
rect 386380 229792 489184 229820
rect 386380 229780 386386 229792
rect 489178 229780 489184 229792
rect 489236 229780 489242 229832
rect 281592 229724 373994 229752
rect 281592 229712 281598 229724
rect 418798 229712 418804 229764
rect 418856 229752 418862 229764
rect 533338 229752 533344 229764
rect 418856 229724 533344 229752
rect 418856 229712 418862 229724
rect 533338 229712 533344 229724
rect 533396 229712 533402 229764
rect 61654 229032 61660 229084
rect 61712 229072 61718 229084
rect 297358 229072 297364 229084
rect 61712 229044 297364 229072
rect 61712 229032 61718 229044
rect 297358 229032 297364 229044
rect 297416 229032 297422 229084
rect 56318 228488 56324 228540
rect 56376 228528 56382 228540
rect 158162 228528 158168 228540
rect 56376 228500 158168 228528
rect 56376 228488 56382 228500
rect 158162 228488 158168 228500
rect 158220 228488 158226 228540
rect 314562 228488 314568 228540
rect 314620 228528 314626 228540
rect 351178 228528 351184 228540
rect 314620 228500 351184 228528
rect 314620 228488 314626 228500
rect 351178 228488 351184 228500
rect 351236 228488 351242 228540
rect 122282 228420 122288 228472
rect 122340 228460 122346 228472
rect 320082 228460 320088 228472
rect 122340 228432 320088 228460
rect 122340 228420 122346 228432
rect 320082 228420 320088 228432
rect 320140 228420 320146 228472
rect 379238 228420 379244 228472
rect 379296 228460 379302 228472
rect 409874 228460 409880 228472
rect 379296 228432 409880 228460
rect 379296 228420 379302 228432
rect 409874 228420 409880 228432
rect 409932 228420 409938 228472
rect 157150 228352 157156 228404
rect 157208 228392 157214 228404
rect 377950 228392 377956 228404
rect 157208 228364 377956 228392
rect 157208 228352 157214 228364
rect 377950 228352 377956 228364
rect 378008 228392 378014 228404
rect 467098 228392 467104 228404
rect 378008 228364 467104 228392
rect 378008 228352 378014 228364
rect 467098 228352 467104 228364
rect 467156 228352 467162 228404
rect 231854 227740 231860 227792
rect 231912 227780 231918 227792
rect 233142 227780 233148 227792
rect 231912 227752 233148 227780
rect 231912 227740 231918 227752
rect 233142 227740 233148 227752
rect 233200 227740 233206 227792
rect 149974 227672 149980 227724
rect 150032 227712 150038 227724
rect 448698 227712 448704 227724
rect 150032 227684 448704 227712
rect 150032 227672 150038 227684
rect 448698 227672 448704 227684
rect 448756 227672 448762 227724
rect 56226 227604 56232 227656
rect 56284 227644 56290 227656
rect 242250 227644 242256 227656
rect 56284 227616 242256 227644
rect 56284 227604 56290 227616
rect 242250 227604 242256 227616
rect 242308 227604 242314 227656
rect 105446 227536 105452 227588
rect 105504 227576 105510 227588
rect 172422 227576 172428 227588
rect 105504 227548 172428 227576
rect 105504 227536 105510 227548
rect 172422 227536 172428 227548
rect 172480 227536 172486 227588
rect 185578 227536 185584 227588
rect 185636 227576 185642 227588
rect 323578 227576 323584 227588
rect 185636 227548 323584 227576
rect 185636 227536 185642 227548
rect 323578 227536 323584 227548
rect 323636 227536 323642 227588
rect 284110 227060 284116 227112
rect 284168 227100 284174 227112
rect 347774 227100 347780 227112
rect 284168 227072 347780 227100
rect 284168 227060 284174 227072
rect 347774 227060 347780 227072
rect 347832 227060 347838 227112
rect 172422 226992 172428 227044
rect 172480 227032 172486 227044
rect 345566 227032 345572 227044
rect 172480 227004 345572 227032
rect 172480 226992 172486 227004
rect 345566 226992 345572 227004
rect 345624 226992 345630 227044
rect 399110 226992 399116 227044
rect 399168 227032 399174 227044
rect 441614 227032 441620 227044
rect 399168 227004 441620 227032
rect 399168 226992 399174 227004
rect 441614 226992 441620 227004
rect 441672 226992 441678 227044
rect 448698 226380 448704 226432
rect 448756 226420 448762 226432
rect 449158 226420 449164 226432
rect 448756 226392 449164 226420
rect 448756 226380 448762 226392
rect 449158 226380 449164 226392
rect 449216 226380 449222 226432
rect 245654 226312 245660 226364
rect 245712 226352 245718 226364
rect 246942 226352 246948 226364
rect 245712 226324 246948 226352
rect 245712 226312 245718 226324
rect 246942 226312 246948 226324
rect 247000 226312 247006 226364
rect 323026 226312 323032 226364
rect 323084 226352 323090 226364
rect 323578 226352 323584 226364
rect 323084 226324 323584 226352
rect 323084 226312 323090 226324
rect 323578 226312 323584 226324
rect 323636 226312 323642 226364
rect 455506 226352 455512 226364
rect 416700 226324 455512 226352
rect 160002 226244 160008 226296
rect 160060 226284 160066 226296
rect 415394 226284 415400 226296
rect 160060 226256 415400 226284
rect 160060 226244 160066 226256
rect 415394 226244 415400 226256
rect 415452 226284 415458 226296
rect 416700 226284 416728 226324
rect 455506 226312 455512 226324
rect 455564 226312 455570 226364
rect 415452 226256 416728 226284
rect 415452 226244 415458 226256
rect 167822 226176 167828 226228
rect 167880 226216 167886 226228
rect 327258 226216 327264 226228
rect 167880 226188 327264 226216
rect 167880 226176 167886 226188
rect 327258 226176 327264 226188
rect 327316 226216 327322 226228
rect 327718 226216 327724 226228
rect 327316 226188 327724 226216
rect 327316 226176 327322 226188
rect 327718 226176 327724 226188
rect 327776 226176 327782 226228
rect 345566 226176 345572 226228
rect 345624 226216 345630 226228
rect 345750 226216 345756 226228
rect 345624 226188 345756 226216
rect 345624 226176 345630 226188
rect 345750 226176 345756 226188
rect 345808 226216 345814 226228
rect 474734 226216 474740 226228
rect 345808 226188 474740 226216
rect 345808 226176 345814 226188
rect 474734 226176 474740 226188
rect 474792 226176 474798 226228
rect 210510 226108 210516 226160
rect 210568 226148 210574 226160
rect 303706 226148 303712 226160
rect 210568 226120 303712 226148
rect 210568 226108 210574 226120
rect 303706 226108 303712 226120
rect 303764 226108 303770 226160
rect 123570 225632 123576 225684
rect 123628 225672 123634 225684
rect 270310 225672 270316 225684
rect 123628 225644 270316 225672
rect 123628 225632 123634 225644
rect 270310 225632 270316 225644
rect 270368 225632 270374 225684
rect 59078 225564 59084 225616
rect 59136 225604 59142 225616
rect 214558 225604 214564 225616
rect 59136 225576 214564 225604
rect 59136 225564 59142 225576
rect 214558 225564 214564 225576
rect 214616 225564 214622 225616
rect 319622 225564 319628 225616
rect 319680 225604 319686 225616
rect 341518 225604 341524 225616
rect 319680 225576 341524 225604
rect 319680 225564 319686 225576
rect 341518 225564 341524 225576
rect 341576 225564 341582 225616
rect 49602 224884 49608 224936
rect 49660 224924 49666 224936
rect 302326 224924 302332 224936
rect 49660 224896 302332 224924
rect 49660 224884 49666 224896
rect 302326 224884 302332 224896
rect 302384 224884 302390 224936
rect 54846 224816 54852 224868
rect 54904 224856 54910 224868
rect 253198 224856 253204 224868
rect 54904 224828 253204 224856
rect 54904 224816 54910 224828
rect 253198 224816 253204 224828
rect 253256 224816 253262 224868
rect 169202 224748 169208 224800
rect 169260 224788 169266 224800
rect 342990 224788 342996 224800
rect 169260 224760 342996 224788
rect 169260 224748 169266 224760
rect 342990 224748 342996 224760
rect 343048 224748 343054 224800
rect 88058 224272 88064 224324
rect 88116 224312 88122 224324
rect 249794 224312 249800 224324
rect 88116 224284 249800 224312
rect 88116 224272 88122 224284
rect 249794 224272 249800 224284
rect 249852 224272 249858 224324
rect 281442 224272 281448 224324
rect 281500 224312 281506 224324
rect 299474 224312 299480 224324
rect 281500 224284 299480 224312
rect 281500 224272 281506 224284
rect 299474 224272 299480 224284
rect 299532 224272 299538 224324
rect 175090 224204 175096 224256
rect 175148 224244 175154 224256
rect 579614 224244 579620 224256
rect 175148 224216 579620 224244
rect 175148 224204 175154 224216
rect 579614 224204 579620 224216
rect 579672 224204 579678 224256
rect 80882 223524 80888 223576
rect 80940 223564 80946 223576
rect 304994 223564 305000 223576
rect 80940 223536 305000 223564
rect 80940 223524 80946 223536
rect 304994 223524 305000 223536
rect 305052 223524 305058 223576
rect 93946 223456 93952 223508
rect 94004 223496 94010 223508
rect 136634 223496 136640 223508
rect 94004 223468 136640 223496
rect 94004 223456 94010 223468
rect 136634 223456 136640 223468
rect 136692 223496 136698 223508
rect 137094 223496 137100 223508
rect 136692 223468 137100 223496
rect 136692 223456 136698 223468
rect 137094 223456 137100 223468
rect 137152 223456 137158 223508
rect 193214 223456 193220 223508
rect 193272 223496 193278 223508
rect 194502 223496 194508 223508
rect 193272 223468 194508 223496
rect 193272 223456 193278 223468
rect 194502 223456 194508 223468
rect 194560 223456 194566 223508
rect 209682 223456 209688 223508
rect 209740 223496 209746 223508
rect 371970 223496 371976 223508
rect 209740 223468 371976 223496
rect 209740 223456 209746 223468
rect 371970 223456 371976 223468
rect 372028 223456 372034 223508
rect 144454 223388 144460 223440
rect 144512 223428 144518 223440
rect 296806 223428 296812 223440
rect 144512 223400 296812 223428
rect 144512 223388 144518 223400
rect 296806 223388 296812 223400
rect 296864 223388 296870 223440
rect 194502 223320 194508 223372
rect 194560 223360 194566 223372
rect 345842 223360 345848 223372
rect 194560 223332 345848 223360
rect 194560 223320 194566 223332
rect 345842 223320 345848 223332
rect 345900 223320 345906 223372
rect 170582 222980 170588 223032
rect 170640 223020 170646 223032
rect 196618 223020 196624 223032
rect 170640 222992 196624 223020
rect 170640 222980 170646 222992
rect 196618 222980 196624 222992
rect 196676 222980 196682 223032
rect 137094 222912 137100 222964
rect 137152 222952 137158 222964
rect 170674 222952 170680 222964
rect 137152 222924 170680 222952
rect 137152 222912 137158 222924
rect 170674 222912 170680 222924
rect 170732 222912 170738 222964
rect 300118 222912 300124 222964
rect 300176 222952 300182 222964
rect 334710 222952 334716 222964
rect 300176 222924 334716 222952
rect 300176 222912 300182 222924
rect 334710 222912 334716 222924
rect 334768 222912 334774 222964
rect 104158 222844 104164 222896
rect 104216 222884 104222 222896
rect 264238 222884 264244 222896
rect 104216 222856 264244 222884
rect 104216 222844 104222 222856
rect 264238 222844 264244 222856
rect 264296 222844 264302 222896
rect 270310 222844 270316 222896
rect 270368 222884 270374 222896
rect 315942 222884 315948 222896
rect 270368 222856 315948 222884
rect 270368 222844 270374 222856
rect 315942 222844 315948 222856
rect 316000 222884 316006 222896
rect 318794 222884 318800 222896
rect 316000 222856 318800 222884
rect 316000 222844 316006 222856
rect 318794 222844 318800 222856
rect 318852 222844 318858 222896
rect 153930 222096 153936 222148
rect 153988 222136 153994 222148
rect 434714 222136 434720 222148
rect 153988 222108 434720 222136
rect 153988 222096 153994 222108
rect 434714 222096 434720 222108
rect 434772 222136 434778 222148
rect 436002 222136 436008 222148
rect 434772 222108 436008 222136
rect 434772 222096 434778 222108
rect 436002 222096 436008 222108
rect 436060 222096 436066 222148
rect 57698 222028 57704 222080
rect 57756 222068 57762 222080
rect 328546 222068 328552 222080
rect 57756 222040 328552 222068
rect 57756 222028 57762 222040
rect 328546 222028 328552 222040
rect 328604 222068 328610 222080
rect 329190 222068 329196 222080
rect 328604 222040 329196 222068
rect 328604 222028 328610 222040
rect 329190 222028 329196 222040
rect 329248 222028 329254 222080
rect 82078 221960 82084 222012
rect 82136 222000 82142 222012
rect 298278 222000 298284 222012
rect 82136 221972 298284 222000
rect 82136 221960 82142 221972
rect 298278 221960 298284 221972
rect 298336 221960 298342 222012
rect 101582 221484 101588 221536
rect 101640 221524 101646 221536
rect 253934 221524 253940 221536
rect 101640 221496 253940 221524
rect 101640 221484 101646 221496
rect 253934 221484 253940 221496
rect 253992 221484 253998 221536
rect 63310 221416 63316 221468
rect 63368 221456 63374 221468
rect 240778 221456 240784 221468
rect 63368 221428 240784 221456
rect 63368 221416 63374 221428
rect 240778 221416 240784 221428
rect 240836 221416 240842 221468
rect 436002 221416 436008 221468
rect 436060 221456 436066 221468
rect 461026 221456 461032 221468
rect 436060 221428 461032 221456
rect 436060 221416 436066 221428
rect 461026 221416 461032 221428
rect 461084 221416 461090 221468
rect 99650 220736 99656 220788
rect 99708 220776 99714 220788
rect 168926 220776 168932 220788
rect 99708 220748 168932 220776
rect 99708 220736 99714 220748
rect 168926 220736 168932 220748
rect 168984 220736 168990 220788
rect 173250 220260 173256 220312
rect 173308 220300 173314 220312
rect 236638 220300 236644 220312
rect 173308 220272 236644 220300
rect 173308 220260 173314 220272
rect 236638 220260 236644 220272
rect 236696 220260 236702 220312
rect 67358 220192 67364 220244
rect 67416 220232 67422 220244
rect 156690 220232 156696 220244
rect 67416 220204 156696 220232
rect 67416 220192 67422 220204
rect 156690 220192 156696 220204
rect 156748 220192 156754 220244
rect 168926 220192 168932 220244
rect 168984 220232 168990 220244
rect 169570 220232 169576 220244
rect 168984 220204 169576 220232
rect 168984 220192 168990 220204
rect 169570 220192 169576 220204
rect 169628 220232 169634 220244
rect 318058 220232 318064 220244
rect 169628 220204 318064 220232
rect 169628 220192 169634 220204
rect 318058 220192 318064 220204
rect 318116 220192 318122 220244
rect 64598 220124 64604 220176
rect 64656 220164 64662 220176
rect 251174 220164 251180 220176
rect 64656 220136 251180 220164
rect 64656 220124 64662 220136
rect 251174 220124 251180 220136
rect 251232 220124 251238 220176
rect 154390 220056 154396 220108
rect 154448 220096 154454 220108
rect 393222 220096 393228 220108
rect 154448 220068 393228 220096
rect 154448 220056 154454 220068
rect 393222 220056 393228 220068
rect 393280 220096 393286 220108
rect 414198 220096 414204 220108
rect 393280 220068 414204 220096
rect 393280 220056 393286 220068
rect 414198 220056 414204 220068
rect 414256 220056 414262 220108
rect 69658 219376 69664 219428
rect 69716 219416 69722 219428
rect 331858 219416 331864 219428
rect 69716 219388 331864 219416
rect 69716 219376 69722 219388
rect 331858 219376 331864 219388
rect 331916 219376 331922 219428
rect 162762 219308 162768 219360
rect 162820 219348 162826 219360
rect 420914 219348 420920 219360
rect 162820 219320 420920 219348
rect 162820 219308 162826 219320
rect 420914 219308 420920 219320
rect 420972 219308 420978 219360
rect 148318 218832 148324 218884
rect 148376 218872 148382 218884
rect 210510 218872 210516 218884
rect 148376 218844 210516 218872
rect 148376 218832 148382 218844
rect 210510 218832 210516 218844
rect 210568 218832 210574 218884
rect 130562 218764 130568 218816
rect 130620 218804 130626 218816
rect 221458 218804 221464 218816
rect 130620 218776 221464 218804
rect 130620 218764 130626 218776
rect 221458 218764 221464 218776
rect 221516 218764 221522 218816
rect 229094 218764 229100 218816
rect 229152 218804 229158 218816
rect 275922 218804 275928 218816
rect 229152 218776 275928 218804
rect 229152 218764 229158 218776
rect 275922 218764 275928 218776
rect 275980 218804 275986 218816
rect 324958 218804 324964 218816
rect 275980 218776 324964 218804
rect 275980 218764 275986 218776
rect 324958 218764 324964 218776
rect 325016 218764 325022 218816
rect 331306 218764 331312 218816
rect 331364 218804 331370 218816
rect 331858 218804 331864 218816
rect 331364 218776 331864 218804
rect 331364 218764 331370 218776
rect 331858 218764 331864 218776
rect 331916 218764 331922 218816
rect 361482 218764 361488 218816
rect 361540 218804 361546 218816
rect 388622 218804 388628 218816
rect 361540 218776 388628 218804
rect 361540 218764 361546 218776
rect 388622 218764 388628 218776
rect 388680 218764 388686 218816
rect 153838 218696 153844 218748
rect 153896 218736 153902 218748
rect 300118 218736 300124 218748
rect 153896 218708 300124 218736
rect 153896 218696 153902 218708
rect 300118 218696 300124 218708
rect 300176 218696 300182 218748
rect 364242 218696 364248 218748
rect 364300 218736 364306 218748
rect 380158 218736 380164 218748
rect 364300 218708 380164 218736
rect 364300 218696 364306 218708
rect 380158 218696 380164 218708
rect 380216 218696 380222 218748
rect 380802 218696 380808 218748
rect 380860 218736 380866 218748
rect 433978 218736 433984 218748
rect 380860 218708 433984 218736
rect 380860 218696 380866 218708
rect 433978 218696 433984 218708
rect 434036 218696 434042 218748
rect 420914 218084 420920 218136
rect 420972 218124 420978 218136
rect 421650 218124 421656 218136
rect 420972 218096 421656 218124
rect 420972 218084 420978 218096
rect 421650 218084 421656 218096
rect 421708 218084 421714 218136
rect 388622 218016 388628 218068
rect 388680 218056 388686 218068
rect 389082 218056 389088 218068
rect 388680 218028 389088 218056
rect 388680 218016 388686 218028
rect 389082 218016 389088 218028
rect 389140 218056 389146 218068
rect 580166 218056 580172 218068
rect 389140 218028 580172 218056
rect 389140 218016 389146 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 142890 217948 142896 218000
rect 142948 217988 142954 218000
rect 300946 217988 300952 218000
rect 142948 217960 300952 217988
rect 142948 217948 142954 217960
rect 300946 217948 300952 217960
rect 301004 217988 301010 218000
rect 385678 217988 385684 218000
rect 301004 217960 385684 217988
rect 301004 217948 301010 217960
rect 385678 217948 385684 217960
rect 385736 217948 385742 218000
rect 111886 217268 111892 217320
rect 111944 217308 111950 217320
rect 270494 217308 270500 217320
rect 111944 217280 270500 217308
rect 111944 217268 111950 217280
rect 270494 217268 270500 217280
rect 270552 217268 270558 217320
rect 419442 217268 419448 217320
rect 419500 217308 419506 217320
rect 526438 217308 526444 217320
rect 419500 217280 526444 217308
rect 419500 217268 419506 217280
rect 526438 217268 526444 217280
rect 526496 217268 526502 217320
rect 164050 216588 164056 216640
rect 164108 216628 164114 216640
rect 378962 216628 378968 216640
rect 164108 216600 378968 216628
rect 164108 216588 164114 216600
rect 378962 216588 378968 216600
rect 379020 216588 379026 216640
rect 160922 216520 160928 216572
rect 160980 216560 160986 216572
rect 334802 216560 334808 216572
rect 160980 216532 334808 216560
rect 160980 216520 160986 216532
rect 334802 216520 334808 216532
rect 334860 216520 334866 216572
rect 3510 216112 3516 216164
rect 3568 216152 3574 216164
rect 8938 216152 8944 216164
rect 3568 216124 8944 216152
rect 3568 216112 3574 216124
rect 8938 216112 8944 216124
rect 8996 216112 9002 216164
rect 151170 215976 151176 216028
rect 151228 216016 151234 216028
rect 276014 216016 276020 216028
rect 151228 215988 276020 216016
rect 151228 215976 151234 215988
rect 276014 215976 276020 215988
rect 276072 215976 276078 216028
rect 337378 215976 337384 216028
rect 337436 216016 337442 216028
rect 439498 216016 439504 216028
rect 337436 215988 439504 216016
rect 337436 215976 337442 215988
rect 439498 215976 439504 215988
rect 439556 215976 439562 216028
rect 74718 215908 74724 215960
rect 74776 215948 74782 215960
rect 252554 215948 252560 215960
rect 74776 215920 252560 215948
rect 74776 215908 74782 215920
rect 252554 215908 252560 215920
rect 252612 215908 252618 215960
rect 423582 215908 423588 215960
rect 423640 215948 423646 215960
rect 530578 215948 530584 215960
rect 423640 215920 530584 215948
rect 423640 215908 423646 215920
rect 530578 215908 530584 215920
rect 530636 215908 530642 215960
rect 333974 215500 333980 215552
rect 334032 215540 334038 215552
rect 334802 215540 334808 215552
rect 334032 215512 334808 215540
rect 334032 215500 334038 215512
rect 334802 215500 334808 215512
rect 334860 215500 334866 215552
rect 42794 215228 42800 215280
rect 42852 215268 42858 215280
rect 44082 215268 44088 215280
rect 42852 215240 44088 215268
rect 42852 215228 42858 215240
rect 44082 215228 44088 215240
rect 44140 215268 44146 215280
rect 120074 215268 120080 215280
rect 44140 215240 120080 215268
rect 44140 215228 44146 215240
rect 120074 215228 120080 215240
rect 120132 215228 120138 215280
rect 147674 215228 147680 215280
rect 147732 215268 147738 215280
rect 358814 215268 358820 215280
rect 147732 215240 358820 215268
rect 147732 215228 147738 215240
rect 358814 215228 358820 215240
rect 358872 215268 358878 215280
rect 359458 215268 359464 215280
rect 358872 215240 359464 215268
rect 358872 215228 358878 215240
rect 359458 215228 359464 215240
rect 359516 215228 359522 215280
rect 60366 215160 60372 215212
rect 60424 215200 60430 215212
rect 291194 215200 291200 215212
rect 60424 215172 291200 215200
rect 60424 215160 60430 215172
rect 291194 215160 291200 215172
rect 291252 215160 291258 215212
rect 96706 215092 96712 215144
rect 96764 215132 96770 215144
rect 147674 215132 147680 215144
rect 96764 215104 147680 215132
rect 96764 215092 96770 215104
rect 147674 215092 147680 215104
rect 147732 215092 147738 215144
rect 1302 214548 1308 214600
rect 1360 214588 1366 214600
rect 42794 214588 42800 214600
rect 1360 214560 42800 214588
rect 1360 214548 1366 214560
rect 42794 214548 42800 214560
rect 42852 214548 42858 214600
rect 86954 213868 86960 213920
rect 87012 213908 87018 213920
rect 144914 213908 144920 213920
rect 87012 213880 144920 213908
rect 87012 213868 87018 213880
rect 144914 213868 144920 213880
rect 144972 213908 144978 213920
rect 146202 213908 146208 213920
rect 144972 213880 146208 213908
rect 144972 213868 144978 213880
rect 146202 213868 146208 213880
rect 146260 213868 146266 213920
rect 146202 213460 146208 213512
rect 146260 213500 146266 213512
rect 202138 213500 202144 213512
rect 146260 213472 202144 213500
rect 146260 213460 146266 213472
rect 202138 213460 202144 213472
rect 202196 213460 202202 213512
rect 141510 213392 141516 213444
rect 141568 213432 141574 213444
rect 229738 213432 229744 213444
rect 141568 213404 229744 213432
rect 141568 213392 141574 213404
rect 229738 213392 229744 213404
rect 229796 213392 229802 213444
rect 133230 213324 133236 213376
rect 133288 213364 133294 213376
rect 247678 213364 247684 213376
rect 133288 213336 247684 213364
rect 133288 213324 133294 213336
rect 247678 213324 247684 213336
rect 247736 213324 247742 213376
rect 271874 213324 271880 213376
rect 271932 213364 271938 213376
rect 293126 213364 293132 213376
rect 271932 213336 293132 213364
rect 271932 213324 271938 213336
rect 293126 213324 293132 213336
rect 293184 213324 293190 213376
rect 126882 213256 126888 213308
rect 126940 213296 126946 213308
rect 273898 213296 273904 213308
rect 126940 213268 273904 213296
rect 126940 213256 126946 213268
rect 273898 213256 273904 213268
rect 273956 213256 273962 213308
rect 311250 213256 311256 213308
rect 311308 213296 311314 213308
rect 404354 213296 404360 213308
rect 311308 213268 404360 213296
rect 311308 213256 311314 213268
rect 404354 213256 404360 213268
rect 404412 213256 404418 213308
rect 14458 213188 14464 213240
rect 14516 213228 14522 213240
rect 83458 213228 83464 213240
rect 14516 213200 83464 213228
rect 14516 213188 14522 213200
rect 83458 213188 83464 213200
rect 83516 213188 83522 213240
rect 147582 213188 147588 213240
rect 147640 213228 147646 213240
rect 391842 213228 391848 213240
rect 147640 213200 391848 213228
rect 147640 213188 147646 213200
rect 391842 213188 391848 213200
rect 391900 213228 391906 213240
rect 429194 213228 429200 213240
rect 391900 213200 429200 213228
rect 391900 213188 391906 213200
rect 429194 213188 429200 213200
rect 429252 213188 429258 213240
rect 77202 212440 77208 212492
rect 77260 212480 77266 212492
rect 367094 212480 367100 212492
rect 77260 212452 367100 212480
rect 77260 212440 77266 212452
rect 367094 212440 367100 212452
rect 367152 212440 367158 212492
rect 164142 212372 164148 212424
rect 164200 212412 164206 212424
rect 376662 212412 376668 212424
rect 164200 212384 376668 212412
rect 164200 212372 164206 212384
rect 376662 212372 376668 212384
rect 376720 212412 376726 212424
rect 382918 212412 382924 212424
rect 376720 212384 382924 212412
rect 376720 212372 376726 212384
rect 382918 212372 382924 212384
rect 382976 212372 382982 212424
rect 162210 211896 162216 211948
rect 162268 211936 162274 211948
rect 274634 211936 274640 211948
rect 162268 211908 274640 211936
rect 162268 211896 162274 211908
rect 274634 211896 274640 211908
rect 274692 211896 274698 211948
rect 48038 211828 48044 211880
rect 48096 211868 48102 211880
rect 211890 211868 211896 211880
rect 48096 211840 211896 211868
rect 48096 211828 48102 211840
rect 211890 211828 211896 211840
rect 211948 211828 211954 211880
rect 170674 211760 170680 211812
rect 170732 211800 170738 211812
rect 346578 211800 346584 211812
rect 170732 211772 346584 211800
rect 170732 211760 170738 211772
rect 346578 211760 346584 211772
rect 346636 211760 346642 211812
rect 210418 211080 210424 211132
rect 210476 211120 210482 211132
rect 335446 211120 335452 211132
rect 210476 211092 335452 211120
rect 210476 211080 210482 211092
rect 335446 211080 335452 211092
rect 335504 211080 335510 211132
rect 84378 210468 84384 210520
rect 84436 210508 84442 210520
rect 264974 210508 264980 210520
rect 84436 210480 264980 210508
rect 84436 210468 84442 210480
rect 264974 210468 264980 210480
rect 265032 210468 265038 210520
rect 128998 210400 129004 210452
rect 129056 210440 129062 210452
rect 345014 210440 345020 210452
rect 129056 210412 345020 210440
rect 129056 210400 129062 210412
rect 345014 210400 345020 210412
rect 345072 210440 345078 210452
rect 351914 210440 351920 210452
rect 345072 210412 351920 210440
rect 345072 210400 345078 210412
rect 351914 210400 351920 210412
rect 351972 210400 351978 210452
rect 377858 210400 377864 210452
rect 377916 210440 377922 210452
rect 451642 210440 451648 210452
rect 377916 210412 451648 210440
rect 377916 210400 377922 210412
rect 451642 210400 451648 210412
rect 451700 210400 451706 210452
rect 41230 209720 41236 209772
rect 41288 209760 41294 209772
rect 322842 209760 322848 209772
rect 41288 209732 322848 209760
rect 41288 209720 41294 209732
rect 322842 209720 322848 209732
rect 322900 209720 322906 209772
rect 95234 209652 95240 209704
rect 95292 209692 95298 209704
rect 140682 209692 140688 209704
rect 95292 209664 140688 209692
rect 95292 209652 95298 209664
rect 140682 209652 140688 209664
rect 140740 209652 140746 209704
rect 147030 209244 147036 209296
rect 147088 209284 147094 209296
rect 239490 209284 239496 209296
rect 147088 209256 239496 209284
rect 147088 209244 147094 209256
rect 239490 209244 239496 209256
rect 239548 209244 239554 209296
rect 171778 209176 171784 209228
rect 171836 209216 171842 209228
rect 304258 209216 304264 209228
rect 171836 209188 304264 209216
rect 171836 209176 171842 209188
rect 304258 209176 304264 209188
rect 304316 209176 304322 209228
rect 140682 209108 140688 209160
rect 140740 209148 140746 209160
rect 319438 209148 319444 209160
rect 140740 209120 319444 209148
rect 140740 209108 140746 209120
rect 319438 209108 319444 209120
rect 319496 209108 319502 209160
rect 398926 209108 398932 209160
rect 398984 209148 398990 209160
rect 449986 209148 449992 209160
rect 398984 209120 449992 209148
rect 398984 209108 398990 209120
rect 449986 209108 449992 209120
rect 450044 209108 450050 209160
rect 43806 209040 43812 209092
rect 43864 209080 43870 209092
rect 233878 209080 233884 209092
rect 43864 209052 233884 209080
rect 43864 209040 43870 209052
rect 233878 209040 233884 209052
rect 233936 209040 233942 209092
rect 371050 209040 371056 209092
rect 371108 209080 371114 209092
rect 431218 209080 431224 209092
rect 371108 209052 431224 209080
rect 371108 209040 371114 209052
rect 431218 209040 431224 209052
rect 431276 209040 431282 209092
rect 311158 208360 311164 208412
rect 311216 208400 311222 208412
rect 316034 208400 316040 208412
rect 311216 208372 316040 208400
rect 311216 208360 311222 208372
rect 316034 208360 316040 208372
rect 316092 208360 316098 208412
rect 49510 208292 49516 208344
rect 49568 208332 49574 208344
rect 322934 208332 322940 208344
rect 49568 208304 322940 208332
rect 49568 208292 49574 208304
rect 322934 208292 322940 208304
rect 322992 208292 322998 208344
rect 124858 207816 124864 207868
rect 124916 207856 124922 207868
rect 265066 207856 265072 207868
rect 124916 207828 265072 207856
rect 124916 207816 124922 207828
rect 265066 207816 265072 207828
rect 265124 207816 265130 207868
rect 131758 207748 131764 207800
rect 131816 207788 131822 207800
rect 281534 207788 281540 207800
rect 131816 207760 281540 207788
rect 131816 207748 131822 207760
rect 281534 207748 281540 207760
rect 281592 207748 281598 207800
rect 102134 207680 102140 207732
rect 102192 207720 102198 207732
rect 252738 207720 252744 207732
rect 102192 207692 252744 207720
rect 102192 207680 102198 207692
rect 252738 207680 252744 207692
rect 252796 207680 252802 207732
rect 61838 207612 61844 207664
rect 61896 207652 61902 207664
rect 277486 207652 277492 207664
rect 61896 207624 277492 207652
rect 61896 207612 61902 207624
rect 277486 207612 277492 207624
rect 277544 207612 277550 207664
rect 110506 206932 110512 206984
rect 110564 206972 110570 206984
rect 111058 206972 111064 206984
rect 110564 206944 111064 206972
rect 110564 206932 110570 206944
rect 111058 206932 111064 206944
rect 111116 206972 111122 206984
rect 153102 206972 153108 206984
rect 111116 206944 153108 206972
rect 111116 206932 111122 206944
rect 153102 206932 153108 206944
rect 153160 206972 153166 206984
rect 443086 206972 443092 206984
rect 153160 206944 443092 206972
rect 153160 206932 153166 206944
rect 443086 206932 443092 206944
rect 443144 206932 443150 206984
rect 476206 206932 476212 206984
rect 476264 206972 476270 206984
rect 579982 206972 579988 206984
rect 476264 206944 579988 206972
rect 476264 206932 476270 206944
rect 579982 206932 579988 206944
rect 580040 206932 580046 206984
rect 107654 206864 107660 206916
rect 107712 206904 107718 206916
rect 155862 206904 155868 206916
rect 107712 206876 155868 206904
rect 107712 206864 107718 206876
rect 155862 206864 155868 206876
rect 155920 206864 155926 206916
rect 227714 206864 227720 206916
rect 227772 206904 227778 206916
rect 346486 206904 346492 206916
rect 227772 206876 346492 206904
rect 227772 206864 227778 206876
rect 346486 206864 346492 206876
rect 346544 206904 346550 206916
rect 347682 206904 347688 206916
rect 346544 206876 347688 206904
rect 346544 206864 346550 206876
rect 347682 206864 347688 206876
rect 347740 206864 347746 206916
rect 155862 206388 155868 206440
rect 155920 206428 155926 206440
rect 257338 206428 257344 206440
rect 155920 206400 257344 206428
rect 155920 206388 155926 206400
rect 257338 206388 257344 206400
rect 257396 206388 257402 206440
rect 89806 206320 89812 206372
rect 89864 206360 89870 206372
rect 252646 206360 252652 206372
rect 89864 206332 252652 206360
rect 89864 206320 89870 206332
rect 252646 206320 252652 206332
rect 252704 206320 252710 206372
rect 67542 206252 67548 206304
rect 67600 206292 67606 206304
rect 280154 206292 280160 206304
rect 67600 206264 280160 206292
rect 67600 206252 67606 206264
rect 280154 206252 280160 206264
rect 280212 206252 280218 206304
rect 347682 206252 347688 206304
rect 347740 206292 347746 206304
rect 452838 206292 452844 206304
rect 347740 206264 452844 206292
rect 347740 206252 347746 206264
rect 452838 206252 452844 206264
rect 452896 206252 452902 206304
rect 467098 206252 467104 206304
rect 467156 206292 467162 206304
rect 476206 206292 476212 206304
rect 467156 206264 476212 206292
rect 467156 206252 467162 206264
rect 476206 206252 476212 206264
rect 476264 206252 476270 206304
rect 84286 205572 84292 205624
rect 84344 205612 84350 205624
rect 125778 205612 125784 205624
rect 84344 205584 125784 205612
rect 84344 205572 84350 205584
rect 125778 205572 125784 205584
rect 125836 205612 125842 205624
rect 126882 205612 126888 205624
rect 125836 205584 126888 205612
rect 125836 205572 125842 205584
rect 126882 205572 126888 205584
rect 126940 205572 126946 205624
rect 158070 205164 158076 205216
rect 158128 205204 158134 205216
rect 247770 205204 247776 205216
rect 158128 205176 247776 205204
rect 158128 205164 158134 205176
rect 247770 205164 247776 205176
rect 247828 205164 247834 205216
rect 151262 205096 151268 205148
rect 151320 205136 151326 205148
rect 263594 205136 263600 205148
rect 151320 205108 263600 205136
rect 151320 205096 151326 205108
rect 263594 205096 263600 205108
rect 263652 205096 263658 205148
rect 126238 205028 126244 205080
rect 126296 205068 126302 205080
rect 259546 205068 259552 205080
rect 126296 205040 259552 205068
rect 126296 205028 126302 205040
rect 259546 205028 259552 205040
rect 259604 205028 259610 205080
rect 66070 204960 66076 205012
rect 66128 205000 66134 205012
rect 251266 205000 251272 205012
rect 66128 204972 251272 205000
rect 66128 204960 66134 204972
rect 251266 204960 251272 204972
rect 251324 204960 251330 205012
rect 373810 204960 373816 205012
rect 373868 205000 373874 205012
rect 435450 205000 435456 205012
rect 373868 204972 435456 205000
rect 373868 204960 373874 204972
rect 435450 204960 435456 204972
rect 435508 204960 435514 205012
rect 179138 204892 179144 204944
rect 179196 204932 179202 204944
rect 405734 204932 405740 204944
rect 179196 204904 405740 204932
rect 179196 204892 179202 204904
rect 405734 204892 405740 204904
rect 405792 204892 405798 204944
rect 421558 204892 421564 204944
rect 421616 204932 421622 204944
rect 464338 204932 464344 204944
rect 421616 204904 464344 204932
rect 421616 204892 421622 204904
rect 464338 204892 464344 204904
rect 464396 204892 464402 204944
rect 126882 204280 126888 204332
rect 126940 204320 126946 204332
rect 193858 204320 193864 204332
rect 126940 204292 193864 204320
rect 126940 204280 126946 204292
rect 193858 204280 193864 204292
rect 193916 204280 193922 204332
rect 84194 204212 84200 204264
rect 84252 204252 84258 204264
rect 126974 204252 126980 204264
rect 84252 204224 126980 204252
rect 84252 204212 84258 204224
rect 126974 204212 126980 204224
rect 127032 204252 127038 204264
rect 127434 204252 127440 204264
rect 127032 204224 127440 204252
rect 127032 204212 127038 204224
rect 127434 204212 127440 204224
rect 127492 204212 127498 204264
rect 144362 203872 144368 203924
rect 144420 203912 144426 203924
rect 242250 203912 242256 203924
rect 144420 203884 242256 203912
rect 144420 203872 144426 203884
rect 242250 203872 242256 203884
rect 242308 203872 242314 203924
rect 242158 203804 242164 203856
rect 242216 203844 242222 203856
rect 351914 203844 351920 203856
rect 242216 203816 351920 203844
rect 242216 203804 242222 203816
rect 351914 203804 351920 203816
rect 351972 203804 351978 203856
rect 142798 203736 142804 203788
rect 142856 203776 142862 203788
rect 277394 203776 277400 203788
rect 142856 203748 277400 203776
rect 142856 203736 142862 203748
rect 277394 203736 277400 203748
rect 277452 203736 277458 203788
rect 115934 203668 115940 203720
rect 115992 203708 115998 203720
rect 254118 203708 254124 203720
rect 115992 203680 254124 203708
rect 115992 203668 115998 203680
rect 254118 203668 254124 203680
rect 254176 203668 254182 203720
rect 53650 203600 53656 203652
rect 53708 203640 53714 203652
rect 267826 203640 267832 203652
rect 53708 203612 267832 203640
rect 53708 203600 53714 203612
rect 267826 203600 267832 203612
rect 267884 203600 267890 203652
rect 127434 203532 127440 203584
rect 127492 203572 127498 203584
rect 352006 203572 352012 203584
rect 127492 203544 352012 203572
rect 127492 203532 127498 203544
rect 352006 203532 352012 203544
rect 352064 203532 352070 203584
rect 381538 203532 381544 203584
rect 381596 203572 381602 203584
rect 458818 203572 458824 203584
rect 381596 203544 458824 203572
rect 381596 203532 381602 203544
rect 458818 203532 458824 203544
rect 458876 203532 458882 203584
rect 130654 202376 130660 202428
rect 130712 202416 130718 202428
rect 246298 202416 246304 202428
rect 130712 202388 246304 202416
rect 130712 202376 130718 202388
rect 246298 202376 246304 202388
rect 246356 202376 246362 202428
rect 144270 202308 144276 202360
rect 144328 202348 144334 202360
rect 192478 202348 192484 202360
rect 144328 202320 192484 202348
rect 144328 202308 144334 202320
rect 192478 202308 192484 202320
rect 192536 202308 192542 202360
rect 193950 202308 193956 202360
rect 194008 202348 194014 202360
rect 335446 202348 335452 202360
rect 194008 202320 335452 202348
rect 194008 202308 194014 202320
rect 335446 202308 335452 202320
rect 335504 202308 335510 202360
rect 170398 202240 170404 202292
rect 170456 202280 170462 202292
rect 316678 202280 316684 202292
rect 170456 202252 316684 202280
rect 170456 202240 170462 202252
rect 316678 202240 316684 202252
rect 316736 202240 316742 202292
rect 89714 202172 89720 202224
rect 89772 202212 89778 202224
rect 252830 202212 252836 202224
rect 89772 202184 252836 202212
rect 89772 202172 89778 202184
rect 252830 202172 252836 202184
rect 252888 202172 252894 202224
rect 39942 202104 39948 202156
rect 40000 202144 40006 202156
rect 287698 202144 287704 202156
rect 40000 202116 287704 202144
rect 40000 202104 40006 202116
rect 287698 202104 287704 202116
rect 287756 202104 287762 202156
rect 395890 202104 395896 202156
rect 395948 202144 395954 202156
rect 444466 202144 444472 202156
rect 395948 202116 444472 202144
rect 395948 202104 395954 202116
rect 444466 202104 444472 202116
rect 444524 202104 444530 202156
rect 421650 201492 421656 201544
rect 421708 201532 421714 201544
rect 422202 201532 422208 201544
rect 421708 201504 422208 201532
rect 421708 201492 421714 201504
rect 422202 201492 422208 201504
rect 422260 201532 422266 201544
rect 427078 201532 427084 201544
rect 422260 201504 427084 201532
rect 422260 201492 422266 201504
rect 427078 201492 427084 201504
rect 427136 201492 427142 201544
rect 246942 201424 246948 201476
rect 247000 201464 247006 201476
rect 298002 201464 298008 201476
rect 247000 201436 298008 201464
rect 247000 201424 247006 201436
rect 298002 201424 298008 201436
rect 298060 201424 298066 201476
rect 196618 200948 196624 201000
rect 196676 200988 196682 201000
rect 271966 200988 271972 201000
rect 196676 200960 271972 200988
rect 196676 200948 196682 200960
rect 271966 200948 271972 200960
rect 272024 200948 272030 201000
rect 110414 200880 110420 200932
rect 110472 200920 110478 200932
rect 255590 200920 255596 200932
rect 110472 200892 255596 200920
rect 110472 200880 110478 200892
rect 255590 200880 255596 200892
rect 255648 200880 255654 200932
rect 57790 200812 57796 200864
rect 57848 200852 57854 200864
rect 222838 200852 222844 200864
rect 57848 200824 222844 200852
rect 57848 200812 57854 200824
rect 222838 200812 222844 200824
rect 222896 200812 222902 200864
rect 79318 200744 79324 200796
rect 79376 200784 79382 200796
rect 322934 200784 322940 200796
rect 79376 200756 322940 200784
rect 79376 200744 79382 200756
rect 322934 200744 322940 200756
rect 322992 200744 322998 200796
rect 298002 200132 298008 200184
rect 298060 200172 298066 200184
rect 451366 200172 451372 200184
rect 298060 200144 451372 200172
rect 298060 200132 298066 200144
rect 451366 200132 451372 200144
rect 451424 200132 451430 200184
rect 233142 200064 233148 200116
rect 233200 200104 233206 200116
rect 284110 200104 284116 200116
rect 233200 200076 284116 200104
rect 233200 200064 233206 200076
rect 284110 200064 284116 200076
rect 284168 200064 284174 200116
rect 117958 199452 117964 199504
rect 118016 199492 118022 199504
rect 273254 199492 273260 199504
rect 118016 199464 273260 199492
rect 118016 199452 118022 199464
rect 273254 199452 273260 199464
rect 273312 199452 273318 199504
rect 94038 199384 94044 199436
rect 94096 199424 94102 199436
rect 255406 199424 255412 199436
rect 94096 199396 255412 199424
rect 94096 199384 94102 199396
rect 255406 199384 255412 199396
rect 255464 199384 255470 199436
rect 282914 198704 282920 198756
rect 282972 198744 282978 198756
rect 284110 198744 284116 198756
rect 282972 198716 284116 198744
rect 282972 198704 282978 198716
rect 284110 198704 284116 198716
rect 284168 198744 284174 198756
rect 451458 198744 451464 198756
rect 284168 198716 451464 198744
rect 284168 198704 284174 198716
rect 451458 198704 451464 198716
rect 451516 198704 451522 198756
rect 76558 198636 76564 198688
rect 76616 198676 76622 198688
rect 330570 198676 330576 198688
rect 76616 198648 330576 198676
rect 76616 198636 76622 198648
rect 330570 198636 330576 198648
rect 330628 198636 330634 198688
rect 145558 198160 145564 198212
rect 145616 198200 145622 198212
rect 232498 198200 232504 198212
rect 145616 198172 232504 198200
rect 145616 198160 145622 198172
rect 232498 198160 232504 198172
rect 232556 198160 232562 198212
rect 149698 198092 149704 198144
rect 149756 198132 149762 198144
rect 269206 198132 269212 198144
rect 149756 198104 269212 198132
rect 149756 198092 149762 198104
rect 269206 198092 269212 198104
rect 269264 198092 269270 198144
rect 92474 198024 92480 198076
rect 92532 198064 92538 198076
rect 261018 198064 261024 198076
rect 92532 198036 261024 198064
rect 92532 198024 92538 198036
rect 261018 198024 261024 198036
rect 261076 198024 261082 198076
rect 292666 198024 292672 198076
rect 292724 198064 292730 198076
rect 441614 198064 441620 198076
rect 292724 198036 441620 198064
rect 292724 198024 292730 198036
rect 441614 198024 441620 198036
rect 441672 198024 441678 198076
rect 93762 197956 93768 198008
rect 93820 197996 93826 198008
rect 356238 197996 356244 198008
rect 93820 197968 356244 197996
rect 93820 197956 93826 197968
rect 356238 197956 356244 197968
rect 356296 197956 356302 198008
rect 439498 197956 439504 198008
rect 439556 197996 439562 198008
rect 538214 197996 538220 198008
rect 439556 197968 538220 197996
rect 439556 197956 439562 197968
rect 538214 197956 538220 197968
rect 538272 197956 538278 198008
rect 329834 197684 329840 197736
rect 329892 197724 329898 197736
rect 330570 197724 330576 197736
rect 329892 197696 330576 197724
rect 329892 197684 329898 197696
rect 330570 197684 330576 197696
rect 330628 197684 330634 197736
rect 94498 197276 94504 197328
rect 94556 197316 94562 197328
rect 354766 197316 354772 197328
rect 94556 197288 354772 197316
rect 94556 197276 94562 197288
rect 354766 197276 354772 197288
rect 354824 197316 354830 197328
rect 355318 197316 355324 197328
rect 354824 197288 355324 197316
rect 354824 197276 354830 197288
rect 355318 197276 355324 197288
rect 355376 197276 355382 197328
rect 335446 197208 335452 197260
rect 335504 197248 335510 197260
rect 535454 197248 535460 197260
rect 335504 197220 535460 197248
rect 335504 197208 335510 197220
rect 535454 197208 535460 197220
rect 535512 197208 535518 197260
rect 141418 196732 141424 196784
rect 141476 196772 141482 196784
rect 269114 196772 269120 196784
rect 141476 196744 269120 196772
rect 141476 196732 141482 196744
rect 269114 196732 269120 196744
rect 269172 196732 269178 196784
rect 133138 196664 133144 196716
rect 133196 196704 133202 196716
rect 263686 196704 263692 196716
rect 133196 196676 263692 196704
rect 133196 196664 133202 196676
rect 263686 196664 263692 196676
rect 263744 196664 263750 196716
rect 70394 196596 70400 196648
rect 70452 196636 70458 196648
rect 254026 196636 254032 196648
rect 70452 196608 254032 196636
rect 70452 196596 70458 196608
rect 254026 196596 254032 196608
rect 254084 196596 254090 196648
rect 98638 195916 98644 195968
rect 98696 195956 98702 195968
rect 354858 195956 354864 195968
rect 98696 195928 354864 195956
rect 98696 195916 98702 195928
rect 354858 195916 354864 195928
rect 354916 195956 354922 195968
rect 355410 195956 355416 195968
rect 354916 195928 355416 195956
rect 354916 195916 354922 195928
rect 355410 195916 355416 195928
rect 355468 195916 355474 195968
rect 162302 195372 162308 195424
rect 162360 195412 162366 195424
rect 267734 195412 267740 195424
rect 162360 195384 267740 195412
rect 162360 195372 162366 195384
rect 267734 195372 267740 195384
rect 267792 195372 267798 195424
rect 138658 195304 138664 195356
rect 138716 195344 138722 195356
rect 281626 195344 281632 195356
rect 138716 195316 281632 195344
rect 138716 195304 138722 195316
rect 281626 195304 281632 195316
rect 281684 195304 281690 195356
rect 52178 195236 52184 195288
rect 52236 195276 52242 195288
rect 236730 195276 236736 195288
rect 52236 195248 236736 195276
rect 52236 195236 52242 195248
rect 236730 195236 236736 195248
rect 236788 195236 236794 195288
rect 264238 195236 264244 195288
rect 264296 195276 264302 195288
rect 356146 195276 356152 195288
rect 264296 195248 356152 195276
rect 264296 195236 264302 195248
rect 356146 195236 356152 195248
rect 356204 195236 356210 195288
rect 134702 194080 134708 194132
rect 134760 194120 134766 194132
rect 262306 194120 262312 194132
rect 134760 194092 262312 194120
rect 134760 194080 134766 194092
rect 262306 194080 262312 194092
rect 262364 194080 262370 194132
rect 100754 194012 100760 194064
rect 100812 194052 100818 194064
rect 278866 194052 278872 194064
rect 100812 194024 278872 194052
rect 100812 194012 100818 194024
rect 278866 194012 278872 194024
rect 278924 194012 278930 194064
rect 55122 193944 55128 193996
rect 55180 193984 55186 193996
rect 239582 193984 239588 193996
rect 55180 193956 239588 193984
rect 55180 193944 55186 193956
rect 239582 193944 239588 193956
rect 239640 193944 239646 193996
rect 177666 193876 177672 193928
rect 177724 193916 177730 193928
rect 376018 193916 376024 193928
rect 177724 193888 376024 193916
rect 177724 193876 177730 193888
rect 376018 193876 376024 193888
rect 376076 193876 376082 193928
rect 391290 193876 391296 193928
rect 391348 193916 391354 193928
rect 454126 193916 454132 193928
rect 391348 193888 454132 193916
rect 391348 193876 391354 193888
rect 454126 193876 454132 193888
rect 454184 193876 454190 193928
rect 136082 193808 136088 193860
rect 136140 193848 136146 193860
rect 338114 193848 338120 193860
rect 136140 193820 338120 193848
rect 136140 193808 136146 193820
rect 338114 193808 338120 193820
rect 338172 193808 338178 193860
rect 390370 193808 390376 193860
rect 390428 193848 390434 193860
rect 520918 193848 520924 193860
rect 390428 193820 520924 193848
rect 390428 193808 390434 193820
rect 520918 193808 520924 193820
rect 520976 193808 520982 193860
rect 427078 193128 427084 193180
rect 427136 193168 427142 193180
rect 580166 193168 580172 193180
rect 427136 193140 580172 193168
rect 427136 193128 427142 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 243538 192720 243544 192772
rect 243596 192760 243602 192772
rect 327074 192760 327080 192772
rect 243596 192732 327080 192760
rect 243596 192720 243602 192732
rect 327074 192720 327080 192732
rect 327132 192720 327138 192772
rect 137278 192652 137284 192704
rect 137336 192692 137342 192704
rect 247862 192692 247868 192704
rect 137336 192664 247868 192692
rect 137336 192652 137342 192664
rect 247862 192652 247868 192664
rect 247920 192652 247926 192704
rect 96614 192584 96620 192636
rect 96672 192624 96678 192636
rect 258166 192624 258172 192636
rect 96672 192596 258172 192624
rect 96672 192584 96678 192596
rect 258166 192584 258172 192596
rect 258224 192584 258230 192636
rect 67450 192516 67456 192568
rect 67508 192556 67514 192568
rect 251358 192556 251364 192568
rect 67508 192528 251364 192556
rect 67508 192516 67514 192528
rect 251358 192516 251364 192528
rect 251416 192516 251422 192568
rect 402238 192516 402244 192568
rect 402296 192556 402302 192568
rect 435542 192556 435548 192568
rect 402296 192528 435548 192556
rect 402296 192516 402302 192528
rect 435542 192516 435548 192528
rect 435600 192516 435606 192568
rect 80790 192448 80796 192500
rect 80848 192488 80854 192500
rect 270586 192488 270592 192500
rect 80848 192460 270592 192488
rect 80848 192448 80854 192460
rect 270586 192448 270592 192460
rect 270644 192448 270650 192500
rect 275830 192448 275836 192500
rect 275888 192488 275894 192500
rect 293034 192488 293040 192500
rect 275888 192460 293040 192488
rect 275888 192448 275894 192460
rect 293034 192448 293040 192460
rect 293092 192448 293098 192500
rect 350626 192448 350632 192500
rect 350684 192488 350690 192500
rect 416958 192488 416964 192500
rect 350684 192460 416964 192488
rect 350684 192448 350690 192460
rect 416958 192448 416964 192460
rect 417016 192448 417022 192500
rect 212534 191768 212540 191820
rect 212592 191808 212598 191820
rect 368474 191808 368480 191820
rect 212592 191780 368480 191808
rect 212592 191768 212598 191780
rect 368474 191768 368480 191780
rect 368532 191808 368538 191820
rect 368934 191808 368940 191820
rect 368532 191780 368940 191808
rect 368532 191768 368538 191780
rect 368934 191768 368940 191780
rect 368992 191768 368998 191820
rect 398098 191768 398104 191820
rect 398156 191808 398162 191820
rect 399478 191808 399484 191820
rect 398156 191780 399484 191808
rect 398156 191768 398162 191780
rect 399478 191768 399484 191780
rect 399536 191768 399542 191820
rect 161382 191224 161388 191276
rect 161440 191264 161446 191276
rect 197998 191264 198004 191276
rect 161440 191236 198004 191264
rect 161440 191224 161446 191236
rect 197998 191224 198004 191236
rect 198056 191224 198062 191276
rect 149882 191156 149888 191208
rect 149940 191196 149946 191208
rect 242158 191196 242164 191208
rect 149940 191168 242164 191196
rect 149940 191156 149946 191168
rect 242158 191156 242164 191168
rect 242216 191156 242222 191208
rect 63218 191088 63224 191140
rect 63276 191128 63282 191140
rect 260834 191128 260840 191140
rect 63276 191100 260840 191128
rect 63276 191088 63282 191100
rect 260834 191088 260840 191100
rect 260892 191088 260898 191140
rect 368934 191088 368940 191140
rect 368992 191128 368998 191140
rect 396074 191128 396080 191140
rect 368992 191100 396080 191128
rect 368992 191088 368998 191100
rect 396074 191088 396080 191100
rect 396132 191088 396138 191140
rect 407758 191088 407764 191140
rect 407816 191128 407822 191140
rect 452930 191128 452936 191140
rect 407816 191100 452936 191128
rect 407816 191088 407822 191100
rect 452930 191088 452936 191100
rect 452988 191088 452994 191140
rect 148410 190000 148416 190052
rect 148468 190040 148474 190052
rect 260926 190040 260932 190052
rect 148468 190012 260932 190040
rect 148468 190000 148474 190012
rect 260926 190000 260932 190012
rect 260984 190000 260990 190052
rect 46842 189932 46848 189984
rect 46900 189972 46906 189984
rect 162118 189972 162124 189984
rect 46900 189944 162124 189972
rect 46900 189932 46906 189944
rect 162118 189932 162124 189944
rect 162176 189932 162182 189984
rect 203518 189932 203524 189984
rect 203576 189972 203582 189984
rect 267918 189972 267924 189984
rect 203576 189944 267924 189972
rect 203576 189932 203582 189944
rect 267918 189932 267924 189944
rect 267976 189932 267982 189984
rect 129182 189864 129188 189916
rect 129240 189904 129246 189916
rect 246390 189904 246396 189916
rect 129240 189876 246396 189904
rect 129240 189864 129246 189876
rect 246390 189864 246396 189876
rect 246448 189864 246454 189916
rect 134794 189796 134800 189848
rect 134852 189836 134858 189848
rect 259454 189836 259460 189848
rect 134852 189808 259460 189836
rect 134852 189796 134858 189808
rect 259454 189796 259460 189808
rect 259512 189796 259518 189848
rect 261478 189796 261484 189848
rect 261536 189836 261542 189848
rect 318150 189836 318156 189848
rect 261536 189808 318156 189836
rect 261536 189796 261542 189808
rect 318150 189796 318156 189808
rect 318208 189796 318214 189848
rect 420270 189796 420276 189848
rect 420328 189836 420334 189848
rect 536926 189836 536932 189848
rect 420328 189808 536932 189836
rect 420328 189796 420334 189808
rect 536926 189796 536932 189808
rect 536984 189796 536990 189848
rect 136174 189728 136180 189780
rect 136232 189768 136238 189780
rect 263778 189768 263784 189780
rect 136232 189740 263784 189768
rect 136232 189728 136238 189740
rect 263778 189728 263784 189740
rect 263836 189728 263842 189780
rect 307018 189728 307024 189780
rect 307076 189768 307082 189780
rect 460198 189768 460204 189780
rect 307076 189740 460204 189768
rect 307076 189728 307082 189740
rect 460198 189728 460204 189740
rect 460256 189728 460262 189780
rect 107562 189048 107568 189100
rect 107620 189088 107626 189100
rect 189902 189088 189908 189100
rect 107620 189060 189908 189088
rect 107620 189048 107626 189060
rect 189902 189048 189908 189060
rect 189960 189048 189966 189100
rect 307018 189048 307024 189100
rect 307076 189088 307082 189100
rect 307662 189088 307668 189100
rect 307076 189060 307668 189088
rect 307076 189048 307082 189060
rect 307662 189048 307668 189060
rect 307720 189048 307726 189100
rect 459554 189048 459560 189100
rect 459612 189088 459618 189100
rect 460198 189088 460204 189100
rect 459612 189060 460204 189088
rect 459612 189048 459618 189060
rect 460198 189048 460204 189060
rect 460256 189048 460262 189100
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 58710 189020 58716 189032
rect 3476 188992 58716 189020
rect 3476 188980 3482 188992
rect 58710 188980 58716 188992
rect 58768 188980 58774 189032
rect 214558 188640 214564 188692
rect 214616 188680 214622 188692
rect 256970 188680 256976 188692
rect 214616 188652 256976 188680
rect 214616 188640 214622 188652
rect 256970 188640 256976 188652
rect 257028 188640 257034 188692
rect 239398 188572 239404 188624
rect 239456 188612 239462 188624
rect 343818 188612 343824 188624
rect 239456 188584 343824 188612
rect 239456 188572 239462 188584
rect 343818 188572 343824 188584
rect 343876 188572 343882 188624
rect 123478 188504 123484 188556
rect 123536 188544 123542 188556
rect 247954 188544 247960 188556
rect 123536 188516 247960 188544
rect 123536 188504 123542 188516
rect 247954 188504 247960 188516
rect 248012 188504 248018 188556
rect 124950 188436 124956 188488
rect 125008 188476 125014 188488
rect 258074 188476 258080 188488
rect 125008 188448 258080 188476
rect 125008 188436 125014 188448
rect 258074 188436 258080 188448
rect 258132 188436 258138 188488
rect 160830 188368 160836 188420
rect 160888 188408 160894 188420
rect 324590 188408 324596 188420
rect 160888 188380 324596 188408
rect 160888 188368 160894 188380
rect 324590 188368 324596 188380
rect 324648 188368 324654 188420
rect 72418 188300 72424 188352
rect 72476 188340 72482 188352
rect 323118 188340 323124 188352
rect 72476 188312 323124 188340
rect 72476 188300 72482 188312
rect 323118 188300 323124 188312
rect 323176 188300 323182 188352
rect 363782 188300 363788 188352
rect 363840 188340 363846 188352
rect 470594 188340 470600 188352
rect 363840 188312 470600 188340
rect 363840 188300 363846 188312
rect 470594 188300 470600 188312
rect 470652 188300 470658 188352
rect 106182 187688 106188 187740
rect 106240 187728 106246 187740
rect 189810 187728 189816 187740
rect 106240 187700 189816 187728
rect 106240 187688 106246 187700
rect 189810 187688 189816 187700
rect 189868 187688 189874 187740
rect 236638 187144 236644 187196
rect 236696 187184 236702 187196
rect 332686 187184 332692 187196
rect 236696 187156 332692 187184
rect 236696 187144 236702 187156
rect 332686 187144 332692 187156
rect 332744 187144 332750 187196
rect 41322 187076 41328 187128
rect 41380 187116 41386 187128
rect 171502 187116 171508 187128
rect 41380 187088 171508 187116
rect 41380 187076 41386 187088
rect 171502 187076 171508 187088
rect 171560 187076 171566 187128
rect 203518 187076 203524 187128
rect 203576 187116 203582 187128
rect 310606 187116 310612 187128
rect 203576 187088 310612 187116
rect 203576 187076 203582 187088
rect 310606 187076 310612 187088
rect 310664 187076 310670 187128
rect 164878 187008 164884 187060
rect 164936 187048 164942 187060
rect 324682 187048 324688 187060
rect 164936 187020 324688 187048
rect 164936 187008 164942 187020
rect 324682 187008 324688 187020
rect 324740 187008 324746 187060
rect 339402 187008 339408 187060
rect 339460 187048 339466 187060
rect 416866 187048 416872 187060
rect 339460 187020 416872 187048
rect 339460 187008 339466 187020
rect 416866 187008 416872 187020
rect 416924 187008 416930 187060
rect 147490 186940 147496 186992
rect 147548 186980 147554 186992
rect 346486 186980 346492 186992
rect 147548 186952 346492 186980
rect 147548 186940 147554 186952
rect 346486 186940 346492 186952
rect 346544 186940 346550 186992
rect 417418 186940 417424 186992
rect 417476 186980 417482 186992
rect 440234 186980 440240 186992
rect 417476 186952 440240 186980
rect 417476 186940 417482 186952
rect 440234 186940 440240 186952
rect 440292 186940 440298 186992
rect 134610 186396 134616 186448
rect 134668 186436 134674 186448
rect 214558 186436 214564 186448
rect 134668 186408 214564 186436
rect 134668 186396 134674 186408
rect 214558 186396 214564 186408
rect 214616 186396 214622 186448
rect 114462 186328 114468 186380
rect 114520 186368 114526 186380
rect 196618 186368 196624 186380
rect 114520 186340 196624 186368
rect 114520 186328 114526 186340
rect 196618 186328 196624 186340
rect 196676 186328 196682 186380
rect 321462 186260 321468 186312
rect 321520 186300 321526 186312
rect 325878 186300 325884 186312
rect 321520 186272 325884 186300
rect 321520 186260 321526 186272
rect 325878 186260 325884 186272
rect 325936 186260 325942 186312
rect 189718 185784 189724 185836
rect 189776 185824 189782 185836
rect 266538 185824 266544 185836
rect 189776 185796 266544 185824
rect 189776 185784 189782 185796
rect 266538 185784 266544 185796
rect 266596 185784 266602 185836
rect 152734 185716 152740 185768
rect 152792 185756 152798 185768
rect 242342 185756 242348 185768
rect 152792 185728 242348 185756
rect 152792 185716 152798 185728
rect 242342 185716 242348 185728
rect 242400 185716 242406 185768
rect 120718 185648 120724 185700
rect 120776 185688 120782 185700
rect 338298 185688 338304 185700
rect 120776 185660 338304 185688
rect 120776 185648 120782 185660
rect 338298 185648 338304 185660
rect 338356 185648 338362 185700
rect 80698 185580 80704 185632
rect 80756 185620 80762 185632
rect 323210 185620 323216 185632
rect 80756 185592 323216 185620
rect 80756 185580 80762 185592
rect 323210 185580 323216 185592
rect 323268 185580 323274 185632
rect 365070 185580 365076 185632
rect 365128 185620 365134 185632
rect 506474 185620 506480 185632
rect 365128 185592 506480 185620
rect 365128 185580 365134 185592
rect 506474 185580 506480 185592
rect 506532 185580 506538 185632
rect 100662 184900 100668 184952
rect 100720 184940 100726 184952
rect 170398 184940 170404 184952
rect 100720 184912 170404 184940
rect 100720 184900 100726 184912
rect 170398 184900 170404 184912
rect 170456 184900 170462 184952
rect 221458 184356 221464 184408
rect 221516 184396 221522 184408
rect 261110 184396 261116 184408
rect 221516 184368 261116 184396
rect 221516 184356 221522 184368
rect 261110 184356 261116 184368
rect 261168 184356 261174 184408
rect 140130 184288 140136 184340
rect 140188 184328 140194 184340
rect 259638 184328 259644 184340
rect 140188 184300 259644 184328
rect 140188 184288 140194 184300
rect 259638 184288 259644 184300
rect 259696 184288 259702 184340
rect 48958 184220 48964 184272
rect 49016 184260 49022 184272
rect 109678 184260 109684 184272
rect 49016 184232 109684 184260
rect 49016 184220 49022 184232
rect 109678 184220 109684 184232
rect 109736 184220 109742 184272
rect 125042 184220 125048 184272
rect 125100 184260 125106 184272
rect 341058 184260 341064 184272
rect 125100 184232 341064 184260
rect 125100 184220 125106 184232
rect 341058 184220 341064 184232
rect 341116 184220 341122 184272
rect 103422 184152 103428 184204
rect 103480 184192 103486 184204
rect 321278 184192 321284 184204
rect 103480 184164 321284 184192
rect 103480 184152 103486 184164
rect 321278 184152 321284 184164
rect 321336 184152 321342 184204
rect 327074 184152 327080 184204
rect 327132 184192 327138 184204
rect 334158 184192 334164 184204
rect 327132 184164 334164 184192
rect 327132 184152 327138 184164
rect 334158 184152 334164 184164
rect 334216 184192 334222 184204
rect 480254 184192 480260 184204
rect 334216 184164 480260 184192
rect 334216 184152 334222 184164
rect 480254 184152 480260 184164
rect 480312 184152 480318 184204
rect 124122 183540 124128 183592
rect 124180 183580 124186 183592
rect 169202 183580 169208 183592
rect 124180 183552 169208 183580
rect 124180 183540 124186 183552
rect 169202 183540 169208 183552
rect 169260 183540 169266 183592
rect 211890 183132 211896 183184
rect 211948 183172 211954 183184
rect 265158 183172 265164 183184
rect 211948 183144 265164 183172
rect 211948 183132 211954 183144
rect 265158 183132 265164 183144
rect 265216 183132 265222 183184
rect 173158 183064 173164 183116
rect 173216 183104 173222 183116
rect 249886 183104 249892 183116
rect 173216 183076 249892 183104
rect 173216 183064 173222 183076
rect 249886 183064 249892 183076
rect 249944 183064 249950 183116
rect 319530 183064 319536 183116
rect 319588 183104 319594 183116
rect 330018 183104 330024 183116
rect 319588 183076 330024 183104
rect 319588 183064 319594 183076
rect 330018 183064 330024 183076
rect 330076 183064 330082 183116
rect 154482 182996 154488 183048
rect 154540 183036 154546 183048
rect 338206 183036 338212 183048
rect 154540 183008 338212 183036
rect 154540 182996 154546 183008
rect 338206 182996 338212 183008
rect 338264 182996 338270 183048
rect 157978 182928 157984 182980
rect 158036 182968 158042 182980
rect 345106 182968 345112 182980
rect 158036 182940 345112 182968
rect 158036 182928 158042 182940
rect 345106 182928 345112 182940
rect 345164 182928 345170 182980
rect 60550 182860 60556 182912
rect 60608 182900 60614 182912
rect 272058 182900 272064 182912
rect 60608 182872 272064 182900
rect 60608 182860 60614 182872
rect 272058 182860 272064 182872
rect 272116 182860 272122 182912
rect 315390 182860 315396 182912
rect 315448 182900 315454 182912
rect 339678 182900 339684 182912
rect 315448 182872 339684 182900
rect 315448 182860 315454 182872
rect 339678 182860 339684 182872
rect 339736 182860 339742 182912
rect 75178 182792 75184 182844
rect 75236 182832 75242 182844
rect 321646 182832 321652 182844
rect 75236 182804 321652 182832
rect 75236 182792 75242 182804
rect 321646 182792 321652 182804
rect 321704 182792 321710 182844
rect 389818 182792 389824 182844
rect 389876 182832 389882 182844
rect 436278 182832 436284 182844
rect 389876 182804 436284 182832
rect 389876 182792 389882 182804
rect 436278 182792 436284 182804
rect 436336 182792 436342 182844
rect 127802 182180 127808 182232
rect 127860 182220 127866 182232
rect 167914 182220 167920 182232
rect 127860 182192 167920 182220
rect 127860 182180 127866 182192
rect 167914 182180 167920 182192
rect 167972 182180 167978 182232
rect 309042 182220 309048 182232
rect 308955 182192 309048 182220
rect 309042 182180 309048 182192
rect 309100 182220 309106 182232
rect 339586 182220 339592 182232
rect 309100 182192 339592 182220
rect 309100 182180 309106 182192
rect 339586 182180 339592 182192
rect 339644 182180 339650 182232
rect 122098 182112 122104 182164
rect 122156 182152 122162 182164
rect 309060 182152 309088 182180
rect 122156 182124 309088 182152
rect 122156 182112 122162 182124
rect 269758 181840 269764 181892
rect 269816 181880 269822 181892
rect 270402 181880 270408 181892
rect 269816 181852 270408 181880
rect 269816 181840 269822 181852
rect 270402 181840 270408 181852
rect 270460 181840 270466 181892
rect 222838 181500 222844 181552
rect 222896 181540 222902 181552
rect 266446 181540 266452 181552
rect 222896 181512 266452 181540
rect 222896 181500 222902 181512
rect 266446 181500 266452 181512
rect 266504 181500 266510 181552
rect 156690 181432 156696 181484
rect 156748 181472 156754 181484
rect 276106 181472 276112 181484
rect 156748 181444 276112 181472
rect 156748 181432 156754 181444
rect 276106 181432 276112 181444
rect 276164 181432 276170 181484
rect 392670 181432 392676 181484
rect 392728 181472 392734 181484
rect 487154 181472 487160 181484
rect 392728 181444 487160 181472
rect 392728 181432 392734 181444
rect 487154 181432 487160 181444
rect 487212 181432 487218 181484
rect 121178 180888 121184 180940
rect 121236 180928 121242 180940
rect 169294 180928 169300 180940
rect 121236 180900 169300 180928
rect 121236 180888 121242 180900
rect 169294 180888 169300 180900
rect 169352 180888 169358 180940
rect 112622 180820 112628 180872
rect 112680 180860 112686 180872
rect 167730 180860 167736 180872
rect 112680 180832 167736 180860
rect 112680 180820 112686 180832
rect 167730 180820 167736 180832
rect 167788 180820 167794 180872
rect 269758 180820 269764 180872
rect 269816 180860 269822 180872
rect 431310 180860 431316 180872
rect 269816 180832 431316 180860
rect 269816 180820 269822 180832
rect 431310 180820 431316 180832
rect 431368 180820 431374 180872
rect 242158 180412 242164 180464
rect 242216 180452 242222 180464
rect 259730 180452 259736 180464
rect 242216 180424 259736 180452
rect 242216 180412 242222 180424
rect 259730 180412 259736 180424
rect 259788 180412 259794 180464
rect 236730 180344 236736 180396
rect 236788 180384 236794 180396
rect 262398 180384 262404 180396
rect 236788 180356 262404 180384
rect 236788 180344 236794 180356
rect 262398 180344 262404 180356
rect 262456 180344 262462 180396
rect 313182 180344 313188 180396
rect 313240 180384 313246 180396
rect 346670 180384 346676 180396
rect 313240 180356 346676 180384
rect 313240 180344 313246 180356
rect 346670 180344 346676 180356
rect 346728 180344 346734 180396
rect 237374 180276 237380 180328
rect 237432 180316 237438 180328
rect 276658 180316 276664 180328
rect 237432 180288 276664 180316
rect 237432 180276 237438 180288
rect 276658 180276 276664 180288
rect 276716 180276 276722 180328
rect 300118 180276 300124 180328
rect 300176 180316 300182 180328
rect 335446 180316 335452 180328
rect 300176 180288 335452 180316
rect 300176 180276 300182 180288
rect 335446 180276 335452 180288
rect 335504 180276 335510 180328
rect 215938 180208 215944 180260
rect 215996 180248 216002 180260
rect 258350 180248 258356 180260
rect 215996 180220 258356 180248
rect 215996 180208 216002 180220
rect 258350 180208 258356 180220
rect 258408 180208 258414 180260
rect 304258 180208 304264 180260
rect 304316 180248 304322 180260
rect 351362 180248 351368 180260
rect 304316 180220 351368 180248
rect 304316 180208 304322 180220
rect 351362 180208 351368 180220
rect 351420 180208 351426 180260
rect 210510 180140 210516 180192
rect 210568 180180 210574 180192
rect 245654 180180 245660 180192
rect 210568 180152 245660 180180
rect 210568 180140 210574 180152
rect 245654 180140 245660 180152
rect 245712 180140 245718 180192
rect 257338 180140 257344 180192
rect 257396 180180 257402 180192
rect 349338 180180 349344 180192
rect 257396 180152 349344 180180
rect 257396 180140 257402 180152
rect 349338 180140 349344 180152
rect 349396 180140 349402 180192
rect 169110 180072 169116 180124
rect 169168 180112 169174 180124
rect 324498 180112 324504 180124
rect 169168 180084 324504 180112
rect 169168 180072 169174 180084
rect 324498 180072 324504 180084
rect 324556 180072 324562 180124
rect 403618 180072 403624 180124
rect 403676 180112 403682 180124
rect 427814 180112 427820 180124
rect 403676 180084 427820 180112
rect 403676 180072 403682 180084
rect 427814 180072 427820 180084
rect 427872 180072 427878 180124
rect 124950 179664 124956 179716
rect 125008 179704 125014 179716
rect 166442 179704 166448 179716
rect 125008 179676 166448 179704
rect 125008 179664 125014 179676
rect 166442 179664 166448 179676
rect 166500 179664 166506 179716
rect 115842 179596 115848 179648
rect 115900 179636 115906 179648
rect 167822 179636 167828 179648
rect 115900 179608 167828 179636
rect 115900 179596 115906 179608
rect 167822 179596 167828 179608
rect 167880 179596 167886 179648
rect 116946 179528 116952 179580
rect 117004 179568 117010 179580
rect 173158 179568 173164 179580
rect 117004 179540 173164 179568
rect 117004 179528 117010 179540
rect 173158 179528 173164 179540
rect 173216 179528 173222 179580
rect 148226 179460 148232 179512
rect 148284 179500 148290 179512
rect 214650 179500 214656 179512
rect 148284 179472 214656 179500
rect 148284 179460 148290 179472
rect 214650 179460 214656 179472
rect 214708 179460 214714 179512
rect 110046 179392 110052 179444
rect 110104 179432 110110 179444
rect 211890 179432 211896 179444
rect 110104 179404 211896 179432
rect 110104 179392 110110 179404
rect 211890 179392 211896 179404
rect 211948 179392 211954 179444
rect 285582 179392 285588 179444
rect 285640 179432 285646 179444
rect 393958 179432 393964 179444
rect 285640 179404 393964 179432
rect 285640 179392 285646 179404
rect 393958 179392 393964 179404
rect 394016 179392 394022 179444
rect 185578 179324 185584 179376
rect 185636 179364 185642 179376
rect 336826 179364 336832 179376
rect 185636 179336 336832 179364
rect 185636 179324 185642 179336
rect 336826 179324 336832 179336
rect 336884 179324 336890 179376
rect 246390 178848 246396 178900
rect 246448 178888 246454 178900
rect 249334 178888 249340 178900
rect 246448 178860 249340 178888
rect 246448 178848 246454 178860
rect 249334 178848 249340 178860
rect 249392 178848 249398 178900
rect 229738 178780 229744 178832
rect 229796 178820 229802 178832
rect 246942 178820 246948 178832
rect 229796 178792 246948 178820
rect 229796 178780 229802 178792
rect 246942 178780 246948 178792
rect 247000 178780 247006 178832
rect 247954 178780 247960 178832
rect 248012 178820 248018 178832
rect 249058 178820 249064 178832
rect 248012 178792 249064 178820
rect 248012 178780 248018 178792
rect 249058 178780 249064 178792
rect 249116 178780 249122 178832
rect 216582 178712 216588 178764
rect 216640 178752 216646 178764
rect 224954 178752 224960 178764
rect 216640 178724 224960 178752
rect 216640 178712 216646 178724
rect 224954 178712 224960 178724
rect 225012 178712 225018 178764
rect 240778 178712 240784 178764
rect 240836 178752 240842 178764
rect 262214 178752 262220 178764
rect 240836 178724 262220 178752
rect 240836 178712 240842 178724
rect 262214 178712 262220 178724
rect 262272 178712 262278 178764
rect 220078 178644 220084 178696
rect 220136 178684 220142 178696
rect 256878 178684 256884 178696
rect 220136 178656 256884 178684
rect 220136 178644 220142 178656
rect 256878 178644 256884 178656
rect 256936 178644 256942 178696
rect 279418 178644 279424 178696
rect 279476 178684 279482 178696
rect 334066 178684 334072 178696
rect 279476 178656 334072 178684
rect 279476 178644 279482 178656
rect 334066 178644 334072 178656
rect 334124 178644 334130 178696
rect 348418 178644 348424 178696
rect 348476 178684 348482 178696
rect 445846 178684 445852 178696
rect 348476 178656 445852 178684
rect 348476 178644 348482 178656
rect 445846 178644 445852 178656
rect 445904 178644 445910 178696
rect 132034 178372 132040 178424
rect 132092 178412 132098 178424
rect 165246 178412 165252 178424
rect 132092 178384 165252 178412
rect 132092 178372 132098 178384
rect 165246 178372 165252 178384
rect 165304 178372 165310 178424
rect 159266 178304 159272 178356
rect 159324 178344 159330 178356
rect 206370 178344 206376 178356
rect 159324 178316 206376 178344
rect 159324 178304 159330 178316
rect 206370 178304 206376 178316
rect 206428 178304 206434 178356
rect 118418 178236 118424 178288
rect 118476 178276 118482 178288
rect 166350 178276 166356 178288
rect 118476 178248 166356 178276
rect 118476 178236 118482 178248
rect 166350 178236 166356 178248
rect 166408 178236 166414 178288
rect 99190 178168 99196 178220
rect 99248 178208 99254 178220
rect 171778 178208 171784 178220
rect 99248 178180 171784 178208
rect 99248 178168 99254 178180
rect 171778 178168 171784 178180
rect 171836 178168 171842 178220
rect 130746 178100 130752 178152
rect 130804 178140 130810 178152
rect 214098 178140 214104 178152
rect 130804 178112 214104 178140
rect 130804 178100 130810 178112
rect 214098 178100 214104 178112
rect 214156 178100 214162 178152
rect 308398 178100 308404 178152
rect 308456 178140 308462 178152
rect 316034 178140 316040 178152
rect 308456 178112 316040 178140
rect 308456 178100 308462 178112
rect 316034 178100 316040 178112
rect 316092 178100 316098 178152
rect 125778 178032 125784 178084
rect 125836 178072 125842 178084
rect 214926 178072 214932 178084
rect 125836 178044 214932 178072
rect 125836 178032 125842 178044
rect 214926 178032 214932 178044
rect 214984 178032 214990 178084
rect 309686 178032 309692 178084
rect 309744 178072 309750 178084
rect 331490 178072 331496 178084
rect 309744 178044 331496 178072
rect 309744 178032 309750 178044
rect 331490 178032 331496 178044
rect 331548 178032 331554 178084
rect 464338 178032 464344 178084
rect 464396 178072 464402 178084
rect 580166 178072 580172 178084
rect 464396 178044 580172 178072
rect 464396 178032 464402 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 97810 177964 97816 178016
rect 97868 178004 97874 178016
rect 134610 178004 134616 178016
rect 97868 177976 134616 178004
rect 97868 177964 97874 177976
rect 134610 177964 134616 177976
rect 134668 177964 134674 178016
rect 166258 177964 166264 178016
rect 166316 178004 166322 178016
rect 309704 178004 309732 178032
rect 166316 177976 309732 178004
rect 166316 177964 166322 177976
rect 247678 177896 247684 177948
rect 247736 177936 247742 177948
rect 249242 177936 249248 177948
rect 247736 177908 249248 177936
rect 247736 177896 247742 177908
rect 249242 177896 249248 177908
rect 249300 177896 249306 177948
rect 316678 177556 316684 177608
rect 316736 177596 316742 177608
rect 325786 177596 325792 177608
rect 316736 177568 325792 177596
rect 316736 177556 316742 177568
rect 325786 177556 325792 177568
rect 325844 177556 325850 177608
rect 239490 177488 239496 177540
rect 239548 177528 239554 177540
rect 250070 177528 250076 177540
rect 239548 177500 250076 177528
rect 239548 177488 239554 177500
rect 250070 177488 250076 177500
rect 250128 177488 250134 177540
rect 320082 177488 320088 177540
rect 320140 177528 320146 177540
rect 329926 177528 329932 177540
rect 320140 177500 329932 177528
rect 320140 177488 320146 177500
rect 329926 177488 329932 177500
rect 329984 177488 329990 177540
rect 242250 177420 242256 177472
rect 242308 177460 242314 177472
rect 258258 177460 258264 177472
rect 242308 177432 258264 177460
rect 242308 177420 242314 177432
rect 258258 177420 258264 177432
rect 258316 177420 258322 177472
rect 318058 177420 318064 177472
rect 318116 177460 318122 177472
rect 332870 177460 332876 177472
rect 318116 177432 332876 177460
rect 318116 177420 318122 177432
rect 332870 177420 332876 177432
rect 332928 177420 332934 177472
rect 239582 177352 239588 177404
rect 239640 177392 239646 177404
rect 256786 177392 256792 177404
rect 239640 177364 256792 177392
rect 239640 177352 239646 177364
rect 256786 177352 256792 177364
rect 256844 177352 256850 177404
rect 309962 177352 309968 177404
rect 310020 177392 310026 177404
rect 329190 177392 329196 177404
rect 310020 177364 329196 177392
rect 310020 177352 310026 177364
rect 329190 177352 329196 177364
rect 329248 177352 329254 177404
rect 167638 177284 167644 177336
rect 167696 177324 167702 177336
rect 251450 177324 251456 177336
rect 167696 177296 251456 177324
rect 167696 177284 167702 177296
rect 251450 177284 251456 177296
rect 251508 177284 251514 177336
rect 299290 177284 299296 177336
rect 299348 177324 299354 177336
rect 311158 177324 311164 177336
rect 299348 177296 311164 177324
rect 299348 177284 299354 177296
rect 311158 177284 311164 177296
rect 311216 177284 311222 177336
rect 318702 177284 318708 177336
rect 318760 177324 318766 177336
rect 342346 177324 342352 177336
rect 318760 177296 342352 177324
rect 318760 177284 318766 177296
rect 342346 177284 342352 177296
rect 342404 177284 342410 177336
rect 134426 176876 134432 176928
rect 134484 176916 134490 176928
rect 164510 176916 164516 176928
rect 134484 176888 164516 176916
rect 134484 176876 134490 176888
rect 164510 176876 164516 176888
rect 164568 176876 164574 176928
rect 128170 176808 128176 176860
rect 128228 176848 128234 176860
rect 166994 176848 167000 176860
rect 128228 176820 167000 176848
rect 128228 176808 128234 176820
rect 166994 176808 167000 176820
rect 167052 176808 167058 176860
rect 108114 176740 108120 176792
rect 108172 176780 108178 176792
rect 169018 176780 169024 176792
rect 108172 176752 169024 176780
rect 108172 176740 108178 176752
rect 169018 176740 169024 176752
rect 169076 176740 169082 176792
rect 309778 176740 309784 176792
rect 309836 176780 309842 176792
rect 313274 176780 313280 176792
rect 309836 176752 313280 176780
rect 309836 176740 309842 176752
rect 313274 176740 313280 176752
rect 313332 176740 313338 176792
rect 344278 176740 344284 176792
rect 344336 176780 344342 176792
rect 429194 176780 429200 176792
rect 344336 176752 429200 176780
rect 344336 176740 344342 176752
rect 429194 176740 429200 176752
rect 429252 176740 429258 176792
rect 100754 176672 100760 176724
rect 100812 176712 100818 176724
rect 171870 176712 171876 176724
rect 100812 176684 171876 176712
rect 100812 176672 100818 176684
rect 171870 176672 171876 176684
rect 171928 176672 171934 176724
rect 295334 176672 295340 176724
rect 295392 176712 295398 176724
rect 296622 176712 296628 176724
rect 295392 176684 296628 176712
rect 295392 176672 295398 176684
rect 296622 176672 296628 176684
rect 296680 176712 296686 176724
rect 444558 176712 444564 176724
rect 296680 176684 444564 176712
rect 296680 176672 296686 176684
rect 444558 176672 444564 176684
rect 444616 176672 444622 176724
rect 135714 176604 135720 176656
rect 135772 176644 135778 176656
rect 213914 176644 213920 176656
rect 135772 176616 213920 176644
rect 135772 176604 135778 176616
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 233878 176604 233884 176656
rect 233936 176644 233942 176656
rect 261202 176644 261208 176656
rect 233936 176616 261208 176644
rect 233936 176604 233942 176616
rect 261202 176604 261208 176616
rect 261260 176604 261266 176656
rect 287698 176604 287704 176656
rect 287756 176644 287762 176656
rect 321462 176644 321468 176656
rect 287756 176616 321468 176644
rect 287756 176604 287762 176616
rect 321462 176604 321468 176616
rect 321520 176604 321526 176656
rect 242342 176536 242348 176588
rect 242400 176576 242406 176588
rect 249150 176576 249156 176588
rect 242400 176548 249156 176576
rect 242400 176536 242406 176548
rect 249150 176536 249156 176548
rect 249208 176536 249214 176588
rect 319438 176468 319444 176520
rect 319496 176508 319502 176520
rect 327074 176508 327080 176520
rect 319496 176480 327080 176508
rect 319496 176468 319502 176480
rect 327074 176468 327080 176480
rect 327132 176468 327138 176520
rect 133138 176196 133144 176248
rect 133196 176236 133202 176248
rect 165522 176236 165528 176248
rect 133196 176208 165528 176236
rect 133196 176196 133202 176208
rect 165522 176196 165528 176208
rect 165580 176196 165586 176248
rect 129458 176128 129464 176180
rect 129516 176168 129522 176180
rect 166166 176168 166172 176180
rect 129516 176140 166172 176168
rect 129516 176128 129522 176140
rect 166166 176128 166172 176140
rect 166224 176128 166230 176180
rect 121914 176060 121920 176112
rect 121972 176100 121978 176112
rect 166258 176100 166264 176112
rect 121972 176072 166264 176100
rect 121972 176060 121978 176072
rect 166258 176060 166264 176072
rect 166316 176060 166322 176112
rect 321370 176060 321376 176112
rect 321428 176100 321434 176112
rect 321738 176100 321744 176112
rect 321428 176072 321744 176100
rect 321428 176060 321434 176072
rect 321738 176060 321744 176072
rect 321796 176060 321802 176112
rect 396718 176060 396724 176112
rect 396776 176100 396782 176112
rect 409966 176100 409972 176112
rect 396776 176072 409972 176100
rect 396776 176060 396782 176072
rect 409966 176060 409972 176072
rect 410024 176060 410030 176112
rect 104618 175992 104624 176044
rect 104676 176032 104682 176044
rect 170490 176032 170496 176044
rect 104676 176004 170496 176032
rect 104676 175992 104682 176004
rect 170490 175992 170496 176004
rect 170548 175992 170554 176044
rect 266262 175992 266268 176044
rect 266320 176032 266326 176044
rect 428458 176032 428464 176044
rect 266320 176004 428464 176032
rect 266320 175992 266326 176004
rect 428458 175992 428464 176004
rect 428516 175992 428522 176044
rect 8938 175924 8944 175976
rect 8996 175964 9002 175976
rect 111058 175964 111064 175976
rect 8996 175936 111064 175964
rect 8996 175924 9002 175936
rect 111058 175924 111064 175936
rect 111116 175924 111122 175976
rect 119430 175924 119436 175976
rect 119488 175964 119494 175976
rect 170582 175964 170588 175976
rect 119488 175936 170588 175964
rect 119488 175924 119494 175936
rect 170582 175924 170588 175936
rect 170640 175924 170646 175976
rect 247770 175924 247776 175976
rect 247828 175964 247834 175976
rect 255498 175964 255504 175976
rect 247828 175936 255504 175964
rect 247828 175924 247834 175936
rect 255498 175924 255504 175936
rect 255556 175924 255562 175976
rect 278038 175924 278044 175976
rect 278096 175964 278102 175976
rect 295334 175964 295340 175976
rect 278096 175936 295340 175964
rect 278096 175924 278102 175936
rect 295334 175924 295340 175936
rect 295392 175924 295398 175976
rect 297358 175924 297364 175976
rect 297416 175964 297422 175976
rect 307662 175964 307668 175976
rect 297416 175936 307668 175964
rect 297416 175924 297422 175936
rect 307662 175924 307668 175936
rect 307720 175924 307726 175976
rect 313918 175924 313924 175976
rect 313976 175964 313982 175976
rect 347958 175964 347964 175976
rect 313976 175936 347964 175964
rect 313976 175924 313982 175936
rect 347958 175924 347964 175936
rect 348016 175964 348022 175976
rect 553394 175964 553400 175976
rect 348016 175936 553400 175964
rect 348016 175924 348022 175936
rect 553394 175924 553400 175936
rect 553452 175924 553458 175976
rect 165522 175176 165528 175228
rect 165580 175216 165586 175228
rect 214006 175216 214012 175228
rect 165580 175188 214012 175216
rect 165580 175176 165586 175188
rect 214006 175176 214012 175188
rect 214064 175176 214070 175228
rect 164510 175108 164516 175160
rect 164568 175148 164574 175160
rect 213914 175148 213920 175160
rect 164568 175120 213920 175148
rect 164568 175108 164574 175120
rect 213914 175108 213920 175120
rect 213972 175108 213978 175160
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 57238 164200 57244 164212
rect 3292 164172 57244 164200
rect 3292 164160 3298 164172
rect 57238 164160 57244 164172
rect 57296 164160 57302 164212
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 13078 150396 13084 150408
rect 3476 150368 13084 150396
rect 3476 150356 3482 150368
rect 13078 150356 13084 150368
rect 13136 150356 13142 150408
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 18598 137952 18604 137964
rect 3292 137924 18604 137952
rect 3292 137912 3298 137924
rect 18598 137912 18604 137924
rect 18656 137912 18662 137964
rect 63402 126964 63408 127016
rect 63460 127004 63466 127016
rect 65518 127004 65524 127016
rect 63460 126976 65524 127004
rect 63460 126964 63466 126976
rect 65518 126964 65524 126976
rect 65576 126964 65582 127016
rect 62022 121456 62028 121508
rect 62080 121496 62086 121508
rect 66070 121496 66076 121508
rect 62080 121468 66076 121496
rect 62080 121456 62086 121468
rect 66070 121456 66076 121468
rect 66128 121456 66134 121508
rect 3418 111528 3424 111580
rect 3476 111568 3482 111580
rect 8938 111568 8944 111580
rect 3476 111540 8944 111568
rect 3476 111528 3482 111540
rect 8938 111528 8944 111540
rect 8996 111528 9002 111580
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 14458 97968 14464 97980
rect 3476 97940 14464 97968
rect 3476 97928 3482 97940
rect 14458 97928 14464 97940
rect 14516 97928 14522 97980
rect 287698 174020 287704 174072
rect 287756 174060 287762 174072
rect 307478 174060 307484 174072
rect 287756 174032 307484 174060
rect 287756 174020 287762 174032
rect 307478 174020 307484 174032
rect 307536 174020 307542 174072
rect 279418 173952 279424 174004
rect 279476 173992 279482 174004
rect 307570 173992 307576 174004
rect 279476 173964 307576 173992
rect 279476 173952 279482 173964
rect 307570 173952 307576 173964
rect 307628 173952 307634 174004
rect 264238 173884 264244 173936
rect 264296 173924 264302 173936
rect 307662 173924 307668 173936
rect 264296 173896 307668 173924
rect 264296 173884 264302 173896
rect 307662 173884 307668 173896
rect 307720 173884 307726 173936
rect 165246 173816 165252 173868
rect 165304 173856 165310 173868
rect 213914 173856 213920 173868
rect 165304 173828 213920 173856
rect 165304 173816 165310 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 340138 173136 340144 173188
rect 340196 173176 340202 173188
rect 516134 173176 516140 173188
rect 340196 173148 516140 173176
rect 340196 173136 340202 173148
rect 516134 173136 516140 173148
rect 516192 173136 516198 173188
rect 290642 172660 290648 172712
rect 290700 172700 290706 172712
rect 307294 172700 307300 172712
rect 290700 172672 307300 172700
rect 290700 172660 290706 172672
rect 307294 172660 307300 172672
rect 307352 172660 307358 172712
rect 287790 172592 287796 172644
rect 287848 172632 287854 172644
rect 307662 172632 307668 172644
rect 287848 172604 307668 172632
rect 287848 172592 287854 172604
rect 307662 172592 307668 172604
rect 307720 172592 307726 172644
rect 271230 172524 271236 172576
rect 271288 172564 271294 172576
rect 306926 172564 306932 172576
rect 271288 172536 306932 172564
rect 271288 172524 271294 172536
rect 306926 172524 306932 172536
rect 306984 172524 306990 172576
rect 166166 172456 166172 172508
rect 166224 172496 166230 172508
rect 213914 172496 213920 172508
rect 166224 172468 213920 172496
rect 166224 172456 166230 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 166994 172388 167000 172440
rect 167052 172428 167058 172440
rect 214006 172428 214012 172440
rect 167052 172400 214012 172428
rect 167052 172388 167058 172400
rect 214006 172388 214012 172400
rect 214064 172388 214070 172440
rect 324314 172388 324320 172440
rect 324372 172428 324378 172440
rect 327074 172428 327080 172440
rect 324372 172400 327080 172428
rect 324372 172388 324378 172400
rect 327074 172388 327080 172400
rect 327132 172388 327138 172440
rect 384298 171776 384304 171828
rect 384356 171816 384362 171828
rect 450078 171816 450084 171828
rect 384356 171788 450084 171816
rect 384356 171776 384362 171788
rect 450078 171776 450084 171788
rect 450136 171776 450142 171828
rect 321738 171368 321744 171420
rect 321796 171408 321802 171420
rect 325786 171408 325792 171420
rect 321796 171380 325792 171408
rect 321796 171368 321802 171380
rect 325786 171368 325792 171380
rect 325844 171368 325850 171420
rect 300118 171232 300124 171284
rect 300176 171272 300182 171284
rect 307478 171272 307484 171284
rect 300176 171244 307484 171272
rect 300176 171232 300182 171244
rect 307478 171232 307484 171244
rect 307536 171232 307542 171284
rect 282362 171164 282368 171216
rect 282420 171204 282426 171216
rect 307570 171204 307576 171216
rect 282420 171176 307576 171204
rect 282420 171164 282426 171176
rect 307570 171164 307576 171176
rect 307628 171164 307634 171216
rect 168006 171096 168012 171148
rect 168064 171136 168070 171148
rect 211798 171136 211804 171148
rect 168064 171108 211804 171136
rect 168064 171096 168070 171108
rect 211798 171096 211804 171108
rect 211856 171096 211862 171148
rect 269942 171096 269948 171148
rect 270000 171136 270006 171148
rect 307662 171136 307668 171148
rect 270000 171108 307668 171136
rect 270000 171096 270006 171108
rect 307662 171096 307668 171108
rect 307720 171096 307726 171148
rect 167914 171028 167920 171080
rect 167972 171068 167978 171080
rect 213914 171068 213920 171080
rect 167972 171040 213920 171068
rect 167972 171028 167978 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 324314 171028 324320 171080
rect 324372 171068 324378 171080
rect 349890 171068 349896 171080
rect 324372 171040 349896 171068
rect 324372 171028 324378 171040
rect 349890 171028 349896 171040
rect 349948 171028 349954 171080
rect 351362 171028 351368 171080
rect 351420 171068 351426 171080
rect 498838 171068 498844 171080
rect 351420 171040 498844 171068
rect 351420 171028 351426 171040
rect 498838 171028 498844 171040
rect 498896 171028 498902 171080
rect 252462 170620 252468 170672
rect 252520 170660 252526 170672
rect 256970 170660 256976 170672
rect 252520 170632 256976 170660
rect 252520 170620 252526 170632
rect 256970 170620 256976 170632
rect 257028 170620 257034 170672
rect 389082 170348 389088 170400
rect 389140 170388 389146 170400
rect 422754 170388 422760 170400
rect 389140 170360 422760 170388
rect 389140 170348 389146 170360
rect 422754 170348 422760 170360
rect 422812 170348 422818 170400
rect 274082 169872 274088 169924
rect 274140 169912 274146 169924
rect 307662 169912 307668 169924
rect 274140 169884 307668 169912
rect 274140 169872 274146 169884
rect 307662 169872 307668 169884
rect 307720 169872 307726 169924
rect 268470 169804 268476 169856
rect 268528 169844 268534 169856
rect 306558 169844 306564 169856
rect 268528 169816 306564 169844
rect 268528 169804 268534 169816
rect 306558 169804 306564 169816
rect 306616 169804 306622 169856
rect 257522 169736 257528 169788
rect 257580 169776 257586 169788
rect 307662 169776 307668 169788
rect 257580 169748 307668 169776
rect 257580 169736 257586 169748
rect 307662 169736 307668 169748
rect 307720 169736 307726 169788
rect 166442 169668 166448 169720
rect 166500 169708 166506 169720
rect 213914 169708 213920 169720
rect 166500 169680 213920 169708
rect 166500 169668 166506 169680
rect 213914 169668 213920 169680
rect 213972 169668 213978 169720
rect 324314 169668 324320 169720
rect 324372 169708 324378 169720
rect 369118 169708 369124 169720
rect 324372 169680 369124 169708
rect 324372 169668 324378 169680
rect 369118 169668 369124 169680
rect 369176 169668 369182 169720
rect 169202 169600 169208 169652
rect 169260 169640 169266 169652
rect 214006 169640 214012 169652
rect 169260 169612 214012 169640
rect 169260 169600 169266 169612
rect 214006 169600 214012 169612
rect 214064 169600 214070 169652
rect 324406 169600 324412 169652
rect 324464 169640 324470 169652
rect 328454 169640 328460 169652
rect 324464 169612 328460 169640
rect 324464 169600 324470 169612
rect 328454 169600 328460 169612
rect 328512 169600 328518 169652
rect 252370 169532 252376 169584
rect 252428 169572 252434 169584
rect 263778 169572 263784 169584
rect 252428 169544 263784 169572
rect 252428 169532 252434 169544
rect 263778 169532 263784 169544
rect 263836 169532 263842 169584
rect 252462 169464 252468 169516
rect 252520 169504 252526 169516
rect 258166 169504 258172 169516
rect 252520 169476 258172 169504
rect 252520 169464 252526 169476
rect 258166 169464 258172 169476
rect 258224 169464 258230 169516
rect 401594 169056 401600 169108
rect 401652 169096 401658 169108
rect 422294 169096 422300 169108
rect 401652 169068 422300 169096
rect 401652 169056 401658 169068
rect 422294 169056 422300 169068
rect 422352 169056 422358 169108
rect 265618 168988 265624 169040
rect 265676 169028 265682 169040
rect 307294 169028 307300 169040
rect 265676 169000 307300 169028
rect 265676 168988 265682 169000
rect 307294 168988 307300 169000
rect 307352 168988 307358 169040
rect 407758 168988 407764 169040
rect 407816 169028 407822 169040
rect 539594 169028 539600 169040
rect 407816 169000 539600 169028
rect 407816 168988 407822 169000
rect 539594 168988 539600 169000
rect 539652 168988 539658 169040
rect 304258 168444 304264 168496
rect 304316 168484 304322 168496
rect 306558 168484 306564 168496
rect 304316 168456 306564 168484
rect 304316 168444 304322 168456
rect 306558 168444 306564 168456
rect 306616 168444 306622 168496
rect 284938 168376 284944 168428
rect 284996 168416 285002 168428
rect 307662 168416 307668 168428
rect 284996 168388 307668 168416
rect 284996 168376 285002 168388
rect 307662 168376 307668 168388
rect 307720 168376 307726 168428
rect 327810 168376 327816 168428
rect 327868 168416 327874 168428
rect 334158 168416 334164 168428
rect 327868 168388 334164 168416
rect 327868 168376 327874 168388
rect 334158 168376 334164 168388
rect 334216 168376 334222 168428
rect 166258 168308 166264 168360
rect 166316 168348 166322 168360
rect 213914 168348 213920 168360
rect 166316 168320 213920 168348
rect 166316 168308 166322 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 252370 168308 252376 168360
rect 252428 168348 252434 168360
rect 263686 168348 263692 168360
rect 252428 168320 263692 168348
rect 252428 168308 252434 168320
rect 263686 168308 263692 168320
rect 263744 168308 263750 168360
rect 169294 168240 169300 168292
rect 169352 168280 169358 168292
rect 214006 168280 214012 168292
rect 169352 168252 214012 168280
rect 169352 168240 169358 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 252462 168240 252468 168292
rect 252520 168280 252526 168292
rect 262306 168280 262312 168292
rect 252520 168252 262312 168280
rect 252520 168240 252526 168252
rect 262306 168240 262312 168252
rect 262364 168240 262370 168292
rect 337286 168172 337292 168224
rect 337344 168212 337350 168224
rect 339494 168212 339500 168224
rect 337344 168184 339500 168212
rect 337344 168172 337350 168184
rect 339494 168172 339500 168184
rect 339552 168172 339558 168224
rect 252002 167696 252008 167748
rect 252060 167736 252066 167748
rect 256878 167736 256884 167748
rect 252060 167708 256884 167736
rect 252060 167696 252066 167708
rect 256878 167696 256884 167708
rect 256936 167696 256942 167748
rect 415394 167628 415400 167680
rect 415452 167668 415458 167680
rect 440326 167668 440332 167680
rect 415452 167640 440332 167668
rect 415452 167628 415458 167640
rect 440326 167628 440332 167640
rect 440384 167628 440390 167680
rect 295978 167152 295984 167204
rect 296036 167192 296042 167204
rect 307662 167192 307668 167204
rect 296036 167164 307668 167192
rect 296036 167152 296042 167164
rect 307662 167152 307668 167164
rect 307720 167152 307726 167204
rect 267090 167084 267096 167136
rect 267148 167124 267154 167136
rect 307478 167124 307484 167136
rect 267148 167096 307484 167124
rect 267148 167084 267154 167096
rect 307478 167084 307484 167096
rect 307536 167084 307542 167136
rect 264330 167016 264336 167068
rect 264388 167056 264394 167068
rect 307570 167056 307576 167068
rect 264388 167028 307576 167056
rect 264388 167016 264394 167028
rect 307570 167016 307576 167028
rect 307628 167016 307634 167068
rect 166350 166948 166356 167000
rect 166408 166988 166414 167000
rect 214098 166988 214104 167000
rect 166408 166960 214104 166988
rect 166408 166948 166414 166960
rect 214098 166948 214104 166960
rect 214156 166948 214162 167000
rect 252370 166948 252376 167000
rect 252428 166988 252434 167000
rect 261018 166988 261024 167000
rect 252428 166960 261024 166988
rect 252428 166948 252434 166960
rect 261018 166948 261024 166960
rect 261076 166948 261082 167000
rect 170582 166880 170588 166932
rect 170640 166920 170646 166932
rect 213914 166920 213920 166932
rect 170640 166892 213920 166920
rect 170640 166880 170646 166892
rect 213914 166880 213920 166892
rect 213972 166880 213978 166932
rect 173158 166812 173164 166864
rect 173216 166852 173222 166864
rect 214006 166852 214012 166864
rect 173216 166824 214012 166852
rect 173216 166812 173222 166824
rect 214006 166812 214012 166824
rect 214064 166812 214070 166864
rect 251910 166268 251916 166320
rect 251968 166308 251974 166320
rect 256786 166308 256792 166320
rect 251968 166280 256792 166308
rect 251968 166268 251974 166280
rect 256786 166268 256792 166280
rect 256844 166268 256850 166320
rect 412634 166268 412640 166320
rect 412692 166308 412698 166320
rect 435358 166308 435364 166320
rect 412692 166280 435364 166308
rect 412692 166268 412698 166280
rect 435358 166268 435364 166280
rect 435416 166268 435422 166320
rect 449158 166268 449164 166320
rect 449216 166308 449222 166320
rect 476206 166308 476212 166320
rect 449216 166280 476212 166308
rect 449216 166268 449222 166280
rect 476206 166268 476212 166280
rect 476264 166268 476270 166320
rect 252462 165860 252468 165912
rect 252520 165900 252526 165912
rect 259730 165900 259736 165912
rect 252520 165872 259736 165900
rect 252520 165860 252526 165872
rect 259730 165860 259736 165872
rect 259788 165860 259794 165912
rect 293218 165724 293224 165776
rect 293276 165764 293282 165776
rect 306374 165764 306380 165776
rect 293276 165736 306380 165764
rect 293276 165724 293282 165736
rect 306374 165724 306380 165736
rect 306432 165724 306438 165776
rect 273990 165656 273996 165708
rect 274048 165696 274054 165708
rect 306558 165696 306564 165708
rect 274048 165668 306564 165696
rect 274048 165656 274054 165668
rect 306558 165656 306564 165668
rect 306616 165656 306622 165708
rect 257614 165588 257620 165640
rect 257672 165628 257678 165640
rect 306466 165628 306472 165640
rect 257672 165600 306472 165628
rect 257672 165588 257678 165600
rect 306466 165588 306472 165600
rect 306524 165588 306530 165640
rect 476206 165588 476212 165640
rect 476264 165628 476270 165640
rect 580166 165628 580172 165640
rect 476264 165600 580172 165628
rect 476264 165588 476270 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 167822 165520 167828 165572
rect 167880 165560 167886 165572
rect 213914 165560 213920 165572
rect 167880 165532 213920 165560
rect 167880 165520 167886 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 251910 165520 251916 165572
rect 251968 165560 251974 165572
rect 267826 165560 267832 165572
rect 251968 165532 267832 165560
rect 251968 165520 251974 165532
rect 267826 165520 267832 165532
rect 267884 165520 267890 165572
rect 324314 165520 324320 165572
rect 324372 165560 324378 165572
rect 337286 165560 337292 165572
rect 324372 165532 337292 165560
rect 324372 165520 324378 165532
rect 337286 165520 337292 165532
rect 337344 165520 337350 165572
rect 251450 165180 251456 165232
rect 251508 165220 251514 165232
rect 252830 165220 252836 165232
rect 251508 165192 252836 165220
rect 251508 165180 251514 165192
rect 252830 165180 252836 165192
rect 252888 165180 252894 165232
rect 252462 164908 252468 164960
rect 252520 164948 252526 164960
rect 258350 164948 258356 164960
rect 252520 164920 258356 164948
rect 252520 164908 252526 164920
rect 258350 164908 258356 164920
rect 258408 164908 258414 164960
rect 268378 164840 268384 164892
rect 268436 164880 268442 164892
rect 307294 164880 307300 164892
rect 268436 164852 307300 164880
rect 268436 164840 268442 164852
rect 307294 164840 307300 164852
rect 307352 164840 307358 164892
rect 337930 164840 337936 164892
rect 337988 164880 337994 164892
rect 426526 164880 426532 164892
rect 337988 164852 426532 164880
rect 337988 164840 337994 164852
rect 426526 164840 426532 164852
rect 426584 164840 426590 164892
rect 306466 164472 306472 164484
rect 296686 164444 306472 164472
rect 275370 164296 275376 164348
rect 275428 164336 275434 164348
rect 296686 164336 296714 164444
rect 306466 164432 306472 164444
rect 306524 164432 306530 164484
rect 306374 164404 306380 164416
rect 275428 164308 296714 164336
rect 300136 164376 306380 164404
rect 275428 164296 275434 164308
rect 258902 164228 258908 164280
rect 258960 164268 258966 164280
rect 300136 164268 300164 164376
rect 306374 164364 306380 164376
rect 306432 164364 306438 164416
rect 258960 164240 300164 164268
rect 258960 164228 258966 164240
rect 300302 164228 300308 164280
rect 300360 164268 300366 164280
rect 306374 164268 306380 164280
rect 300360 164240 306380 164268
rect 300360 164228 300366 164240
rect 306374 164228 306380 164240
rect 306432 164228 306438 164280
rect 167730 164160 167736 164212
rect 167788 164200 167794 164212
rect 214006 164200 214012 164212
rect 167788 164172 214012 164200
rect 167788 164160 167794 164172
rect 214006 164160 214012 164172
rect 214064 164160 214070 164212
rect 252186 164160 252192 164212
rect 252244 164200 252250 164212
rect 266538 164200 266544 164212
rect 252244 164172 266544 164200
rect 252244 164160 252250 164172
rect 266538 164160 266544 164172
rect 266596 164160 266602 164212
rect 324406 164160 324412 164212
rect 324464 164200 324470 164212
rect 331214 164200 331220 164212
rect 324464 164172 331220 164200
rect 324464 164160 324470 164172
rect 331214 164160 331220 164172
rect 331272 164160 331278 164212
rect 196618 164092 196624 164144
rect 196676 164132 196682 164144
rect 213914 164132 213920 164144
rect 196676 164104 213920 164132
rect 196676 164092 196682 164104
rect 213914 164092 213920 164104
rect 213972 164092 213978 164144
rect 251910 164092 251916 164144
rect 251968 164132 251974 164144
rect 265158 164132 265164 164144
rect 251968 164104 265164 164132
rect 251968 164092 251974 164104
rect 265158 164092 265164 164104
rect 265216 164092 265222 164144
rect 324314 164024 324320 164076
rect 324372 164064 324378 164076
rect 327166 164064 327172 164076
rect 324372 164036 327172 164064
rect 324372 164024 324378 164036
rect 327166 164024 327172 164036
rect 327224 164024 327230 164076
rect 332410 163480 332416 163532
rect 332468 163520 332474 163532
rect 340966 163520 340972 163532
rect 332468 163492 340972 163520
rect 332468 163480 332474 163492
rect 340966 163480 340972 163492
rect 341024 163480 341030 163532
rect 410518 163480 410524 163532
rect 410576 163520 410582 163532
rect 443638 163520 443644 163532
rect 410576 163492 443644 163520
rect 410576 163480 410582 163492
rect 443638 163480 443644 163492
rect 443696 163480 443702 163532
rect 283558 163004 283564 163056
rect 283616 163044 283622 163056
rect 306374 163044 306380 163056
rect 283616 163016 306380 163044
rect 283616 163004 283622 163016
rect 306374 163004 306380 163016
rect 306432 163004 306438 163056
rect 263042 162936 263048 162988
rect 263100 162976 263106 162988
rect 306558 162976 306564 162988
rect 263100 162948 306564 162976
rect 263100 162936 263106 162948
rect 306558 162936 306564 162948
rect 306616 162936 306622 162988
rect 253290 162868 253296 162920
rect 253348 162908 253354 162920
rect 306466 162908 306472 162920
rect 253348 162880 306472 162908
rect 253348 162868 253354 162880
rect 306466 162868 306472 162880
rect 306524 162868 306530 162920
rect 211890 162800 211896 162852
rect 211948 162840 211954 162852
rect 213914 162840 213920 162852
rect 211948 162812 213920 162840
rect 211948 162800 211954 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 252462 162800 252468 162852
rect 252520 162840 252526 162852
rect 262398 162840 262404 162852
rect 252520 162812 262404 162840
rect 252520 162800 252526 162812
rect 262398 162800 262404 162812
rect 262456 162800 262462 162852
rect 252094 162732 252100 162784
rect 252152 162772 252158 162784
rect 261110 162772 261116 162784
rect 252152 162744 261116 162772
rect 252152 162732 252158 162744
rect 261110 162732 261116 162744
rect 261168 162732 261174 162784
rect 439590 162120 439596 162172
rect 439648 162160 439654 162172
rect 447134 162160 447140 162172
rect 439648 162132 447140 162160
rect 439648 162120 439654 162132
rect 447134 162120 447140 162132
rect 447192 162120 447198 162172
rect 287882 161576 287888 161628
rect 287940 161616 287946 161628
rect 306466 161616 306472 161628
rect 287940 161588 306472 161616
rect 287940 161576 287946 161588
rect 306466 161576 306472 161588
rect 306524 161576 306530 161628
rect 252462 161508 252468 161560
rect 252520 161548 252526 161560
rect 259546 161548 259552 161560
rect 252520 161520 259552 161548
rect 252520 161508 252526 161520
rect 259546 161508 259552 161520
rect 259604 161508 259610 161560
rect 264606 161508 264612 161560
rect 264664 161548 264670 161560
rect 306374 161548 306380 161560
rect 264664 161520 306380 161548
rect 264664 161508 264670 161520
rect 306374 161508 306380 161520
rect 306432 161508 306438 161560
rect 254578 161440 254584 161492
rect 254636 161480 254642 161492
rect 306558 161480 306564 161492
rect 254636 161452 306564 161480
rect 254636 161440 254642 161452
rect 306558 161440 306564 161452
rect 306616 161440 306622 161492
rect 169018 161372 169024 161424
rect 169076 161412 169082 161424
rect 213914 161412 213920 161424
rect 169076 161384 213920 161412
rect 169076 161372 169082 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 324314 161372 324320 161424
rect 324372 161412 324378 161424
rect 335630 161412 335636 161424
rect 324372 161384 335636 161412
rect 324372 161372 324378 161384
rect 335630 161372 335636 161384
rect 335688 161372 335694 161424
rect 189902 161304 189908 161356
rect 189960 161344 189966 161356
rect 214006 161344 214012 161356
rect 189960 161316 214012 161344
rect 189960 161304 189966 161316
rect 214006 161304 214012 161316
rect 214064 161304 214070 161356
rect 251358 160828 251364 160880
rect 251416 160868 251422 160880
rect 254118 160868 254124 160880
rect 251416 160840 254124 160868
rect 251416 160828 251422 160840
rect 254118 160828 254124 160840
rect 254176 160828 254182 160880
rect 252462 160692 252468 160744
rect 252520 160732 252526 160744
rect 258258 160732 258264 160744
rect 252520 160704 258264 160732
rect 252520 160692 252526 160704
rect 258258 160692 258264 160704
rect 258316 160692 258322 160744
rect 326430 160692 326436 160744
rect 326488 160732 326494 160744
rect 338298 160732 338304 160744
rect 326488 160704 338304 160732
rect 326488 160692 326494 160704
rect 338298 160692 338304 160704
rect 338356 160692 338362 160744
rect 398650 160692 398656 160744
rect 398708 160732 398714 160744
rect 536834 160732 536840 160744
rect 398708 160704 536840 160732
rect 398708 160692 398714 160704
rect 536834 160692 536840 160704
rect 536892 160692 536898 160744
rect 251910 160352 251916 160404
rect 251968 160392 251974 160404
rect 255498 160392 255504 160404
rect 251968 160364 255504 160392
rect 251968 160352 251974 160364
rect 255498 160352 255504 160364
rect 255556 160352 255562 160404
rect 302970 160216 302976 160268
rect 303028 160256 303034 160268
rect 306558 160256 306564 160268
rect 303028 160228 306564 160256
rect 303028 160216 303034 160228
rect 306558 160216 306564 160228
rect 306616 160216 306622 160268
rect 280890 160148 280896 160200
rect 280948 160188 280954 160200
rect 306466 160188 306472 160200
rect 280948 160160 306472 160188
rect 280948 160148 280954 160160
rect 306466 160148 306472 160160
rect 306524 160148 306530 160200
rect 261570 160080 261576 160132
rect 261628 160120 261634 160132
rect 306374 160120 306380 160132
rect 261628 160092 306380 160120
rect 261628 160080 261634 160092
rect 306374 160080 306380 160092
rect 306432 160080 306438 160132
rect 170490 160012 170496 160064
rect 170548 160052 170554 160064
rect 214006 160052 214012 160064
rect 170548 160024 214012 160052
rect 170548 160012 170554 160024
rect 214006 160012 214012 160024
rect 214064 160012 214070 160064
rect 324314 160012 324320 160064
rect 324372 160052 324378 160064
rect 332410 160052 332416 160064
rect 324372 160024 332416 160052
rect 324372 160012 324378 160024
rect 332410 160012 332416 160024
rect 332468 160012 332474 160064
rect 189810 159944 189816 159996
rect 189868 159984 189874 159996
rect 213914 159984 213920 159996
rect 189868 159956 213920 159984
rect 189868 159944 189874 159956
rect 213914 159944 213920 159956
rect 213972 159944 213978 159996
rect 424318 159400 424324 159452
rect 424376 159440 424382 159452
rect 449066 159440 449072 159452
rect 424376 159412 449072 159440
rect 424376 159400 424382 159412
rect 449066 159400 449072 159412
rect 449124 159400 449130 159452
rect 171870 159332 171876 159384
rect 171928 159372 171934 159384
rect 214098 159372 214104 159384
rect 171928 159344 214104 159372
rect 171928 159332 171934 159344
rect 214098 159332 214104 159344
rect 214156 159332 214162 159384
rect 376110 159332 376116 159384
rect 376168 159372 376174 159384
rect 455598 159372 455604 159384
rect 376168 159344 455604 159372
rect 376168 159332 376174 159344
rect 455598 159332 455604 159344
rect 455656 159332 455662 159384
rect 292206 158856 292212 158908
rect 292264 158896 292270 158908
rect 306374 158896 306380 158908
rect 292264 158868 306380 158896
rect 292264 158856 292270 158868
rect 306374 158856 306380 158868
rect 306432 158856 306438 158908
rect 272518 158788 272524 158840
rect 272576 158828 272582 158840
rect 306558 158828 306564 158840
rect 272576 158800 306564 158828
rect 272576 158788 272582 158800
rect 306558 158788 306564 158800
rect 306616 158788 306622 158840
rect 260282 158720 260288 158772
rect 260340 158760 260346 158772
rect 306466 158760 306472 158772
rect 260340 158732 306472 158760
rect 260340 158720 260346 158732
rect 306466 158720 306472 158732
rect 306524 158720 306530 158772
rect 252370 158652 252376 158704
rect 252428 158692 252434 158704
rect 272058 158692 272064 158704
rect 252428 158664 272064 158692
rect 252428 158652 252434 158664
rect 272058 158652 272064 158664
rect 272116 158652 272122 158704
rect 324406 158652 324412 158704
rect 324464 158692 324470 158704
rect 334066 158692 334072 158704
rect 324464 158664 334072 158692
rect 324464 158652 324470 158664
rect 334066 158652 334072 158664
rect 334124 158652 334130 158704
rect 252462 158584 252468 158636
rect 252520 158624 252526 158636
rect 265066 158624 265072 158636
rect 252520 158596 265072 158624
rect 252520 158584 252526 158596
rect 265066 158584 265072 158596
rect 265124 158584 265130 158636
rect 324314 158584 324320 158636
rect 324372 158624 324378 158636
rect 330018 158624 330024 158636
rect 324372 158596 330024 158624
rect 324372 158584 324378 158596
rect 330018 158584 330024 158596
rect 330076 158584 330082 158636
rect 293402 157496 293408 157548
rect 293460 157536 293466 157548
rect 306374 157536 306380 157548
rect 293460 157508 306380 157536
rect 293460 157496 293466 157508
rect 306374 157496 306380 157508
rect 306432 157496 306438 157548
rect 262858 157428 262864 157480
rect 262916 157468 262922 157480
rect 306558 157468 306564 157480
rect 262916 157440 306564 157468
rect 262916 157428 262922 157440
rect 306558 157428 306564 157440
rect 306616 157428 306622 157480
rect 257338 157360 257344 157412
rect 257396 157400 257402 157412
rect 306466 157400 306472 157412
rect 257396 157372 306472 157400
rect 257396 157360 257402 157372
rect 306466 157360 306472 157372
rect 306524 157360 306530 157412
rect 170398 157292 170404 157344
rect 170456 157332 170462 157344
rect 213914 157332 213920 157344
rect 170456 157304 213920 157332
rect 170456 157292 170462 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 252462 157292 252468 157344
rect 252520 157332 252526 157344
rect 267918 157332 267924 157344
rect 252520 157304 267924 157332
rect 252520 157292 252526 157304
rect 267918 157292 267924 157304
rect 267976 157292 267982 157344
rect 324406 157292 324412 157344
rect 324464 157332 324470 157344
rect 332870 157332 332876 157344
rect 324464 157304 332876 157332
rect 324464 157292 324470 157304
rect 332870 157292 332876 157304
rect 332928 157292 332934 157344
rect 324314 157020 324320 157072
rect 324372 157060 324378 157072
rect 325970 157060 325976 157072
rect 324372 157032 325976 157060
rect 324372 157020 324378 157032
rect 325970 157020 325976 157032
rect 326028 157020 326034 157072
rect 411898 156612 411904 156664
rect 411956 156652 411962 156664
rect 449250 156652 449256 156664
rect 411956 156624 449256 156652
rect 411956 156612 411962 156624
rect 449250 156612 449256 156624
rect 449308 156612 449314 156664
rect 285122 156068 285128 156120
rect 285180 156108 285186 156120
rect 307662 156108 307668 156120
rect 285180 156080 307668 156108
rect 285180 156068 285186 156080
rect 307662 156068 307668 156080
rect 307720 156068 307726 156120
rect 258994 156000 259000 156052
rect 259052 156040 259058 156052
rect 307478 156040 307484 156052
rect 259052 156012 307484 156040
rect 259052 156000 259058 156012
rect 307478 156000 307484 156012
rect 307536 156000 307542 156052
rect 258810 155932 258816 155984
rect 258868 155972 258874 155984
rect 307570 155972 307576 155984
rect 258868 155944 307576 155972
rect 258868 155932 258874 155944
rect 307570 155932 307576 155944
rect 307628 155932 307634 155984
rect 171778 155864 171784 155916
rect 171836 155904 171842 155916
rect 213914 155904 213920 155916
rect 171836 155876 213920 155904
rect 171836 155864 171842 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 252462 155864 252468 155916
rect 252520 155904 252526 155916
rect 278866 155904 278872 155916
rect 252520 155876 278872 155904
rect 252520 155864 252526 155876
rect 278866 155864 278872 155876
rect 278924 155864 278930 155916
rect 324314 155864 324320 155916
rect 324372 155904 324378 155916
rect 356054 155904 356060 155916
rect 324372 155876 356060 155904
rect 324372 155864 324378 155876
rect 356054 155864 356060 155876
rect 356112 155864 356118 155916
rect 252370 155796 252376 155848
rect 252428 155836 252434 155848
rect 274634 155836 274640 155848
rect 252428 155808 274640 155836
rect 252428 155796 252434 155808
rect 274634 155796 274640 155808
rect 274692 155796 274698 155848
rect 252462 155728 252468 155780
rect 252520 155768 252526 155780
rect 264974 155768 264980 155780
rect 252520 155740 264980 155768
rect 252520 155728 252526 155740
rect 264974 155728 264980 155740
rect 265032 155728 265038 155780
rect 261662 155184 261668 155236
rect 261720 155224 261726 155236
rect 306926 155224 306932 155236
rect 261720 155196 306932 155224
rect 261720 155184 261726 155196
rect 306926 155184 306932 155196
rect 306984 155184 306990 155236
rect 351270 155184 351276 155236
rect 351328 155224 351334 155236
rect 451550 155224 451556 155236
rect 351328 155196 451556 155224
rect 351328 155184 351334 155196
rect 451550 155184 451556 155196
rect 451608 155184 451614 155236
rect 279510 154640 279516 154692
rect 279568 154680 279574 154692
rect 307478 154680 307484 154692
rect 279568 154652 307484 154680
rect 279568 154640 279574 154652
rect 307478 154640 307484 154652
rect 307536 154640 307542 154692
rect 262950 154572 262956 154624
rect 263008 154612 263014 154624
rect 306742 154612 306748 154624
rect 263008 154584 306748 154612
rect 263008 154572 263014 154584
rect 306742 154572 306748 154584
rect 306800 154572 306806 154624
rect 251726 154504 251732 154556
rect 251784 154544 251790 154556
rect 277486 154544 277492 154556
rect 251784 154516 277492 154544
rect 251784 154504 251790 154516
rect 277486 154504 277492 154516
rect 277544 154504 277550 154556
rect 324314 154300 324320 154352
rect 324372 154340 324378 154352
rect 326430 154340 326436 154352
rect 324372 154312 326436 154340
rect 324372 154300 324378 154312
rect 326430 154300 326436 154312
rect 326488 154300 326494 154352
rect 251174 154232 251180 154284
rect 251232 154272 251238 154284
rect 254026 154272 254032 154284
rect 251232 154244 254032 154272
rect 251232 154232 251238 154244
rect 254026 154232 254032 154244
rect 254084 154232 254090 154284
rect 254762 153824 254768 153876
rect 254820 153864 254826 153876
rect 307386 153864 307392 153876
rect 254820 153836 307392 153864
rect 254820 153824 254826 153836
rect 307386 153824 307392 153836
rect 307444 153824 307450 153876
rect 408402 153824 408408 153876
rect 408460 153864 408466 153876
rect 426618 153864 426624 153876
rect 408460 153836 426624 153864
rect 408460 153824 408466 153836
rect 426618 153824 426624 153836
rect 426676 153824 426682 153876
rect 195238 153280 195244 153332
rect 195296 153320 195302 153332
rect 214006 153320 214012 153332
rect 195296 153292 214012 153320
rect 195296 153280 195302 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 301498 153280 301504 153332
rect 301556 153320 301562 153332
rect 307570 153320 307576 153332
rect 301556 153292 307576 153320
rect 301556 153280 301562 153292
rect 307570 153280 307576 153292
rect 307628 153280 307634 153332
rect 431586 153320 431592 153332
rect 412606 153292 431592 153320
rect 185578 153212 185584 153264
rect 185636 153252 185642 153264
rect 213914 153252 213920 153264
rect 185636 153224 213920 153252
rect 185636 153212 185642 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 271138 153212 271144 153264
rect 271196 153252 271202 153264
rect 307662 153252 307668 153264
rect 271196 153224 307668 153252
rect 271196 153212 271202 153224
rect 307662 153212 307668 153224
rect 307720 153212 307726 153264
rect 329190 153212 329196 153264
rect 329248 153252 329254 153264
rect 412606 153252 412634 153292
rect 431586 153280 431592 153292
rect 431644 153280 431650 153332
rect 329248 153224 412634 153252
rect 329248 153212 329254 153224
rect 429654 153212 429660 153264
rect 429712 153252 429718 153264
rect 431954 153252 431960 153264
rect 429712 153224 431960 153252
rect 429712 153212 429718 153224
rect 431954 153212 431960 153224
rect 432012 153212 432018 153264
rect 252002 153144 252008 153196
rect 252060 153184 252066 153196
rect 271966 153184 271972 153196
rect 252060 153156 271972 153184
rect 252060 153144 252066 153156
rect 271966 153144 271972 153156
rect 272024 153144 272030 153196
rect 324314 153144 324320 153196
rect 324372 153184 324378 153196
rect 339678 153184 339684 153196
rect 324372 153156 339684 153184
rect 324372 153144 324378 153156
rect 339678 153144 339684 153156
rect 339736 153144 339742 153196
rect 252462 153076 252468 153128
rect 252520 153116 252526 153128
rect 269206 153116 269212 153128
rect 252520 153088 269212 153116
rect 252520 153076 252526 153088
rect 269206 153076 269212 153088
rect 269264 153076 269270 153128
rect 398926 152600 398932 152652
rect 398984 152640 398990 152652
rect 420178 152640 420184 152652
rect 398984 152612 420184 152640
rect 398984 152600 398990 152612
rect 420178 152600 420184 152612
rect 420236 152600 420242 152652
rect 375190 152532 375196 152584
rect 375248 152572 375254 152584
rect 418706 152572 418712 152584
rect 375248 152544 418712 152572
rect 375248 152532 375254 152544
rect 418706 152532 418712 152544
rect 418764 152532 418770 152584
rect 425790 152532 425796 152584
rect 425848 152572 425854 152584
rect 455414 152572 455420 152584
rect 425848 152544 455420 152572
rect 425848 152532 425854 152544
rect 455414 152532 455420 152544
rect 455472 152532 455478 152584
rect 257430 152464 257436 152516
rect 257488 152504 257494 152516
rect 307478 152504 307484 152516
rect 257488 152476 307484 152504
rect 257488 152464 257494 152476
rect 307478 152464 307484 152476
rect 307536 152464 307542 152516
rect 338758 152464 338764 152516
rect 338816 152504 338822 152516
rect 400214 152504 400220 152516
rect 338816 152476 400220 152504
rect 338816 152464 338822 152476
rect 400214 152464 400220 152476
rect 400272 152464 400278 152516
rect 405642 152464 405648 152516
rect 405700 152504 405706 152516
rect 456886 152504 456892 152516
rect 405700 152476 456892 152504
rect 405700 152464 405706 152476
rect 456886 152464 456892 152476
rect 456944 152464 456950 152516
rect 458818 152464 458824 152516
rect 458876 152504 458882 152516
rect 580166 152504 580172 152516
rect 458876 152476 580172 152504
rect 458876 152464 458882 152476
rect 580166 152464 580172 152476
rect 580224 152464 580230 152516
rect 204898 151920 204904 151972
rect 204956 151960 204962 151972
rect 213914 151960 213920 151972
rect 204956 151932 213920 151960
rect 204956 151920 204962 151932
rect 213914 151920 213920 151932
rect 213972 151920 213978 151972
rect 257706 151920 257712 151972
rect 257764 151960 257770 151972
rect 306558 151960 306564 151972
rect 257764 151932 306564 151960
rect 257764 151920 257770 151932
rect 306558 151920 306564 151932
rect 306616 151920 306622 151972
rect 191098 151852 191104 151904
rect 191156 151892 191162 151904
rect 214006 151892 214012 151904
rect 191156 151864 214012 151892
rect 191156 151852 191162 151864
rect 214006 151852 214012 151864
rect 214064 151852 214070 151904
rect 278130 151852 278136 151904
rect 278188 151892 278194 151904
rect 307662 151892 307668 151904
rect 278188 151864 307668 151892
rect 278188 151852 278194 151864
rect 307662 151852 307668 151864
rect 307720 151852 307726 151904
rect 189810 151784 189816 151836
rect 189868 151824 189874 151836
rect 213914 151824 213920 151836
rect 189868 151796 213920 151824
rect 189868 151784 189874 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 324314 151716 324320 151768
rect 324372 151756 324378 151768
rect 341058 151756 341064 151768
rect 324372 151728 341064 151756
rect 324372 151716 324378 151728
rect 341058 151716 341064 151728
rect 341116 151716 341122 151768
rect 343818 151716 343824 151768
rect 343876 151756 343882 151768
rect 535546 151756 535552 151768
rect 343876 151728 535552 151756
rect 343876 151716 343882 151728
rect 535546 151716 535552 151728
rect 535604 151716 535610 151768
rect 252462 151648 252468 151700
rect 252520 151688 252526 151700
rect 270494 151688 270500 151700
rect 252520 151660 270500 151688
rect 252520 151648 252526 151660
rect 270494 151648 270500 151660
rect 270552 151648 270558 151700
rect 252370 151580 252376 151632
rect 252428 151620 252434 151632
rect 273254 151620 273260 151632
rect 252428 151592 273260 151620
rect 252428 151580 252434 151592
rect 273254 151580 273260 151592
rect 273312 151580 273318 151632
rect 324314 151308 324320 151360
rect 324372 151348 324378 151360
rect 327350 151348 327356 151360
rect 324372 151320 327356 151348
rect 324372 151308 324378 151320
rect 327350 151308 327356 151320
rect 327408 151308 327414 151360
rect 365622 151104 365628 151156
rect 365680 151144 365686 151156
rect 406470 151144 406476 151156
rect 365680 151116 406476 151144
rect 365680 151104 365686 151116
rect 406470 151104 406476 151116
rect 406528 151104 406534 151156
rect 182082 151036 182088 151088
rect 182140 151076 182146 151088
rect 206278 151076 206284 151088
rect 182140 151048 206284 151076
rect 182140 151036 182146 151048
rect 206278 151036 206284 151048
rect 206336 151036 206342 151088
rect 363690 151036 363696 151088
rect 363748 151076 363754 151088
rect 412266 151076 412272 151088
rect 363748 151048 412272 151076
rect 363748 151036 363754 151048
rect 412266 151036 412272 151048
rect 412324 151036 412330 151088
rect 289354 150560 289360 150612
rect 289412 150600 289418 150612
rect 307478 150600 307484 150612
rect 289412 150572 307484 150600
rect 289412 150560 289418 150572
rect 307478 150560 307484 150572
rect 307536 150560 307542 150612
rect 196710 150492 196716 150544
rect 196768 150532 196774 150544
rect 213914 150532 213920 150544
rect 196768 150504 213920 150532
rect 196768 150492 196774 150504
rect 213914 150492 213920 150504
rect 213972 150492 213978 150544
rect 273898 150492 273904 150544
rect 273956 150532 273962 150544
rect 307294 150532 307300 150544
rect 273956 150504 307300 150532
rect 273956 150492 273962 150504
rect 307294 150492 307300 150504
rect 307352 150492 307358 150544
rect 194042 150424 194048 150476
rect 194100 150464 194106 150476
rect 214006 150464 214012 150476
rect 194100 150436 214012 150464
rect 194100 150424 194106 150436
rect 214006 150424 214012 150436
rect 214064 150424 214070 150476
rect 256142 150424 256148 150476
rect 256200 150464 256206 150476
rect 307662 150464 307668 150476
rect 256200 150436 307668 150464
rect 256200 150424 256206 150436
rect 307662 150424 307668 150436
rect 307720 150424 307726 150476
rect 211798 150356 211804 150408
rect 211856 150396 211862 150408
rect 213914 150396 213920 150408
rect 211856 150368 213920 150396
rect 211856 150356 211862 150368
rect 213914 150356 213920 150368
rect 213972 150356 213978 150408
rect 251910 150356 251916 150408
rect 251968 150396 251974 150408
rect 281626 150396 281632 150408
rect 251968 150368 281632 150396
rect 251968 150356 251974 150368
rect 281626 150356 281632 150368
rect 281684 150356 281690 150408
rect 251542 150288 251548 150340
rect 251600 150328 251606 150340
rect 255406 150328 255412 150340
rect 251600 150300 255412 150328
rect 251600 150288 251606 150300
rect 255406 150288 255412 150300
rect 255464 150288 255470 150340
rect 252646 149744 252652 149796
rect 252704 149784 252710 149796
rect 262214 149784 262220 149796
rect 252704 149756 262220 149784
rect 252704 149744 252710 149756
rect 262214 149744 262220 149756
rect 262272 149744 262278 149796
rect 379422 149744 379428 149796
rect 379480 149784 379486 149796
rect 397546 149784 397552 149796
rect 379480 149756 397552 149784
rect 379480 149744 379486 149756
rect 397546 149744 397552 149756
rect 397604 149744 397610 149796
rect 254854 149676 254860 149728
rect 254912 149716 254918 149728
rect 306650 149716 306656 149728
rect 254912 149688 306656 149716
rect 254912 149676 254918 149688
rect 306650 149676 306656 149688
rect 306708 149676 306714 149728
rect 387242 149676 387248 149728
rect 387300 149716 387306 149728
rect 454218 149716 454224 149728
rect 387300 149688 454224 149716
rect 387300 149676 387306 149688
rect 454218 149676 454224 149688
rect 454276 149676 454282 149728
rect 272610 149200 272616 149252
rect 272668 149240 272674 149252
rect 307478 149240 307484 149252
rect 272668 149212 307484 149240
rect 272668 149200 272674 149212
rect 307478 149200 307484 149212
rect 307536 149200 307542 149252
rect 296254 149132 296260 149184
rect 296312 149172 296318 149184
rect 307662 149172 307668 149184
rect 296312 149144 307668 149172
rect 296312 149132 296318 149144
rect 307662 149132 307668 149144
rect 307720 149132 307726 149184
rect 355318 149064 355324 149116
rect 355376 149104 355382 149116
rect 420270 149104 420276 149116
rect 355376 149076 420276 149104
rect 355376 149064 355382 149076
rect 420270 149064 420276 149076
rect 420328 149064 420334 149116
rect 206370 148996 206376 149048
rect 206428 149036 206434 149048
rect 213914 149036 213920 149048
rect 206428 149008 213920 149036
rect 206428 148996 206434 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 252462 148996 252468 149048
rect 252520 149036 252526 149048
rect 276014 149036 276020 149048
rect 252520 149008 276020 149036
rect 252520 148996 252526 149008
rect 276014 148996 276020 149008
rect 276072 148996 276078 149048
rect 324406 148996 324412 149048
rect 324464 149036 324470 149048
rect 352006 149036 352012 149048
rect 324464 149008 352012 149036
rect 324464 148996 324470 149008
rect 352006 148996 352012 149008
rect 352064 149036 352070 149048
rect 371878 149036 371884 149048
rect 352064 149008 371884 149036
rect 352064 148996 352070 149008
rect 371878 148996 371884 149008
rect 371936 148996 371942 149048
rect 435450 148996 435456 149048
rect 435508 149036 435514 149048
rect 442718 149036 442724 149048
rect 435508 149008 442724 149036
rect 435508 148996 435514 149008
rect 442718 148996 442724 149008
rect 442776 148996 442782 149048
rect 324314 148928 324320 148980
rect 324372 148968 324378 148980
rect 329926 148968 329932 148980
rect 324372 148940 329932 148968
rect 324372 148928 324378 148940
rect 329926 148928 329932 148940
rect 329984 148928 329990 148980
rect 431310 148724 431316 148776
rect 431368 148764 431374 148776
rect 434162 148764 434168 148776
rect 431368 148736 434168 148764
rect 431368 148724 431374 148736
rect 434162 148724 434168 148736
rect 434220 148724 434226 148776
rect 409874 148520 409880 148572
rect 409932 148560 409938 148572
rect 410702 148560 410708 148572
rect 409932 148532 410708 148560
rect 409932 148520 409938 148532
rect 410702 148520 410708 148532
rect 410760 148520 410766 148572
rect 426434 148520 426440 148572
rect 426492 148560 426498 148572
rect 427446 148560 427452 148572
rect 426492 148532 427452 148560
rect 426492 148520 426498 148532
rect 427446 148520 427452 148532
rect 427504 148520 427510 148572
rect 446490 148520 446496 148572
rect 446548 148560 446554 148572
rect 449618 148560 449624 148572
rect 446548 148532 449624 148560
rect 446548 148520 446554 148532
rect 449618 148520 449624 148532
rect 449676 148520 449682 148572
rect 419442 148492 419448 148504
rect 412606 148464 419448 148492
rect 387242 148384 387248 148436
rect 387300 148424 387306 148436
rect 412606 148424 412634 148464
rect 419442 148452 419448 148464
rect 419500 148492 419506 148504
rect 421282 148492 421288 148504
rect 419500 148464 421288 148492
rect 419500 148452 419506 148464
rect 421282 148452 421288 148464
rect 421340 148452 421346 148504
rect 387300 148396 412634 148424
rect 387300 148384 387306 148396
rect 428458 148384 428464 148436
rect 428516 148424 428522 148436
rect 435450 148424 435456 148436
rect 428516 148396 435456 148424
rect 428516 148384 428522 148396
rect 435450 148384 435456 148396
rect 435508 148384 435514 148436
rect 252002 148316 252008 148368
rect 252060 148356 252066 148368
rect 273990 148356 273996 148368
rect 252060 148328 273996 148356
rect 252060 148316 252066 148328
rect 273990 148316 273996 148328
rect 274048 148316 274054 148368
rect 360010 148316 360016 148368
rect 360068 148356 360074 148368
rect 400030 148356 400036 148368
rect 360068 148328 400036 148356
rect 360068 148316 360074 148328
rect 400030 148316 400036 148328
rect 400088 148316 400094 148368
rect 425146 148316 425152 148368
rect 425204 148356 425210 148368
rect 436738 148356 436744 148368
rect 425204 148328 436744 148356
rect 425204 148316 425210 148328
rect 436738 148316 436744 148328
rect 436796 148316 436802 148368
rect 466546 148316 466552 148368
rect 466604 148356 466610 148368
rect 522298 148356 522304 148368
rect 466604 148328 522304 148356
rect 466604 148316 466610 148328
rect 522298 148316 522304 148328
rect 522356 148316 522362 148368
rect 435542 148248 435548 148300
rect 435600 148288 435606 148300
rect 438026 148288 438032 148300
rect 435600 148260 438032 148288
rect 435600 148248 435606 148260
rect 438026 148248 438032 148260
rect 438084 148248 438090 148300
rect 436094 148180 436100 148232
rect 436152 148220 436158 148232
rect 442994 148220 443000 148232
rect 436152 148192 443000 148220
rect 436152 148180 436158 148192
rect 442994 148180 443000 148192
rect 443052 148180 443058 148232
rect 438670 148112 438676 148164
rect 438728 148152 438734 148164
rect 439590 148152 439596 148164
rect 438728 148124 439596 148152
rect 438728 148112 438734 148124
rect 439590 148112 439596 148124
rect 439648 148112 439654 148164
rect 402606 147976 402612 148028
rect 402664 148016 402670 148028
rect 403618 148016 403624 148028
rect 402664 147988 403624 148016
rect 402664 147976 402670 147988
rect 403618 147976 403624 147988
rect 403676 147976 403682 148028
rect 443638 147976 443644 148028
rect 443696 148016 443702 148028
rect 446030 148016 446036 148028
rect 443696 147988 446036 148016
rect 443696 147976 443702 147988
rect 446030 147976 446036 147988
rect 446088 147976 446094 148028
rect 274174 147772 274180 147824
rect 274232 147812 274238 147824
rect 307478 147812 307484 147824
rect 274232 147784 307484 147812
rect 274232 147772 274238 147784
rect 307478 147772 307484 147784
rect 307536 147772 307542 147824
rect 396810 147772 396816 147824
rect 396868 147812 396874 147824
rect 405826 147812 405832 147824
rect 396868 147784 405832 147812
rect 396868 147772 396874 147784
rect 405826 147772 405832 147784
rect 405884 147772 405890 147824
rect 441890 147772 441896 147824
rect 441948 147812 441954 147824
rect 442718 147812 442724 147824
rect 441948 147784 442724 147812
rect 441948 147772 441954 147784
rect 442718 147772 442724 147784
rect 442776 147812 442782 147824
rect 455966 147812 455972 147824
rect 442776 147784 455972 147812
rect 442776 147772 442782 147784
rect 455966 147772 455972 147784
rect 456024 147772 456030 147824
rect 271322 147704 271328 147756
rect 271380 147744 271386 147756
rect 307570 147744 307576 147756
rect 271380 147716 307576 147744
rect 271380 147704 271386 147716
rect 307570 147704 307576 147716
rect 307628 147704 307634 147756
rect 377398 147704 377404 147756
rect 377456 147744 377462 147756
rect 418890 147744 418896 147756
rect 377456 147716 418896 147744
rect 377456 147704 377462 147716
rect 418890 147704 418896 147716
rect 418948 147704 418954 147756
rect 448974 147704 448980 147756
rect 449032 147744 449038 147756
rect 466546 147744 466552 147756
rect 449032 147716 466552 147744
rect 449032 147704 449038 147716
rect 466546 147704 466552 147716
rect 466604 147704 466610 147756
rect 260374 147636 260380 147688
rect 260432 147676 260438 147688
rect 307662 147676 307668 147688
rect 260432 147648 307668 147676
rect 260432 147636 260438 147648
rect 307662 147636 307668 147648
rect 307720 147636 307726 147688
rect 373350 147636 373356 147688
rect 373408 147676 373414 147688
rect 416866 147676 416872 147688
rect 373408 147648 416872 147676
rect 373408 147636 373414 147648
rect 416866 147636 416872 147648
rect 416924 147636 416930 147688
rect 429102 147636 429108 147688
rect 429160 147676 429166 147688
rect 456058 147676 456064 147688
rect 429160 147648 456064 147676
rect 429160 147636 429166 147648
rect 456058 147636 456064 147648
rect 456116 147636 456122 147688
rect 339402 147568 339408 147620
rect 339460 147608 339466 147620
rect 421558 147608 421564 147620
rect 339460 147580 421564 147608
rect 339460 147568 339466 147580
rect 421558 147568 421564 147580
rect 421616 147608 421622 147620
rect 421926 147608 421932 147620
rect 421616 147580 421932 147608
rect 421616 147568 421622 147580
rect 421926 147568 421932 147580
rect 421984 147568 421990 147620
rect 446398 147568 446404 147620
rect 446456 147608 446462 147620
rect 451550 147608 451556 147620
rect 446456 147580 451556 147608
rect 446456 147568 446462 147580
rect 451550 147568 451556 147580
rect 451608 147568 451614 147620
rect 252370 147500 252376 147552
rect 252428 147540 252434 147552
rect 276106 147540 276112 147552
rect 252428 147512 276112 147540
rect 252428 147500 252434 147512
rect 276106 147500 276112 147512
rect 276164 147500 276170 147552
rect 324314 147500 324320 147552
rect 324372 147540 324378 147552
rect 345106 147540 345112 147552
rect 324372 147512 345112 147540
rect 324372 147500 324378 147512
rect 345106 147500 345112 147512
rect 345164 147500 345170 147552
rect 252462 147432 252468 147484
rect 252520 147472 252526 147484
rect 277394 147472 277400 147484
rect 252520 147444 277400 147472
rect 252520 147432 252526 147444
rect 277394 147432 277400 147444
rect 277452 147432 277458 147484
rect 251174 146956 251180 147008
rect 251232 146996 251238 147008
rect 253934 146996 253940 147008
rect 251232 146968 253940 146996
rect 251232 146956 251238 146968
rect 253934 146956 253940 146968
rect 253992 146956 253998 147008
rect 392578 146956 392584 147008
rect 392636 146996 392642 147008
rect 400122 146996 400128 147008
rect 392636 146968 400128 146996
rect 392636 146956 392642 146968
rect 400122 146956 400128 146968
rect 400180 146956 400186 147008
rect 447778 146956 447784 147008
rect 447836 146996 447842 147008
rect 459554 146996 459560 147008
rect 447836 146968 459560 146996
rect 447836 146956 447842 146968
rect 459554 146956 459560 146968
rect 459612 146956 459618 147008
rect 251542 146888 251548 146940
rect 251600 146928 251606 146940
rect 263594 146928 263600 146940
rect 251600 146900 263600 146928
rect 251600 146888 251606 146900
rect 263594 146888 263600 146900
rect 263652 146888 263658 146940
rect 327718 146888 327724 146940
rect 327776 146928 327782 146940
rect 338206 146928 338212 146940
rect 327776 146900 338212 146928
rect 327776 146888 327782 146900
rect 338206 146888 338212 146900
rect 338264 146928 338270 146940
rect 339402 146928 339408 146940
rect 338264 146900 339408 146928
rect 338264 146888 338270 146900
rect 339402 146888 339408 146900
rect 339460 146888 339466 146940
rect 395798 146888 395804 146940
rect 395856 146928 395862 146940
rect 402974 146928 402980 146940
rect 395856 146900 402980 146928
rect 395856 146888 395862 146900
rect 402974 146888 402980 146900
rect 403032 146888 403038 146940
rect 431218 146888 431224 146940
rect 431276 146928 431282 146940
rect 454310 146928 454316 146940
rect 431276 146900 454316 146928
rect 431276 146888 431282 146900
rect 454310 146888 454316 146900
rect 454368 146888 454374 146940
rect 381538 146412 381544 146464
rect 381596 146452 381602 146464
rect 407758 146452 407764 146464
rect 381596 146424 407764 146452
rect 381596 146412 381602 146424
rect 407758 146412 407764 146424
rect 407816 146412 407822 146464
rect 304534 146344 304540 146396
rect 304592 146384 304598 146396
rect 307478 146384 307484 146396
rect 304592 146356 307484 146384
rect 304592 146344 304598 146356
rect 307478 146344 307484 146356
rect 307536 146344 307542 146396
rect 331858 146344 331864 146396
rect 331916 146384 331922 146396
rect 432598 146384 432604 146396
rect 331916 146356 432604 146384
rect 331916 146344 331922 146356
rect 432598 146344 432604 146356
rect 432656 146344 432662 146396
rect 433518 146344 433524 146396
rect 433576 146384 433582 146396
rect 433978 146384 433984 146396
rect 433576 146356 433984 146384
rect 433576 146344 433582 146356
rect 433978 146344 433984 146356
rect 434036 146384 434042 146396
rect 460198 146384 460204 146396
rect 434036 146356 460204 146384
rect 434036 146344 434042 146356
rect 460198 146344 460204 146356
rect 460256 146344 460262 146396
rect 188338 146276 188344 146328
rect 188396 146316 188402 146328
rect 213914 146316 213920 146328
rect 188396 146288 213920 146316
rect 188396 146276 188402 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 254670 146276 254676 146328
rect 254728 146316 254734 146328
rect 307662 146316 307668 146328
rect 254728 146288 307668 146316
rect 254728 146276 254734 146288
rect 307662 146276 307668 146288
rect 307720 146276 307726 146328
rect 400122 146276 400128 146328
rect 400180 146316 400186 146328
rect 580350 146316 580356 146328
rect 400180 146288 580356 146316
rect 400180 146276 400186 146288
rect 580350 146276 580356 146288
rect 580408 146276 580414 146328
rect 251726 146208 251732 146260
rect 251784 146248 251790 146260
rect 259638 146248 259644 146260
rect 251784 146220 259644 146248
rect 251784 146208 251790 146220
rect 259638 146208 259644 146220
rect 259696 146208 259702 146260
rect 324314 146208 324320 146260
rect 324372 146248 324378 146260
rect 346670 146248 346676 146260
rect 324372 146220 346676 146248
rect 324372 146208 324378 146220
rect 346670 146208 346676 146220
rect 346728 146208 346734 146260
rect 251910 146140 251916 146192
rect 251968 146180 251974 146192
rect 266446 146180 266452 146192
rect 251968 146152 266452 146180
rect 251968 146140 251974 146152
rect 266446 146140 266452 146152
rect 266504 146140 266510 146192
rect 324406 146140 324412 146192
rect 324464 146180 324470 146192
rect 331306 146180 331312 146192
rect 324464 146152 331312 146180
rect 324464 146140 324470 146152
rect 331306 146140 331312 146152
rect 331364 146140 331370 146192
rect 252094 146072 252100 146124
rect 252152 146112 252158 146124
rect 270586 146112 270592 146124
rect 252152 146084 270592 146112
rect 252152 146072 252158 146084
rect 270586 146072 270592 146084
rect 270644 146072 270650 146124
rect 446766 145936 446772 145988
rect 446824 145976 446830 145988
rect 449250 145976 449256 145988
rect 446824 145948 449256 145976
rect 446824 145936 446830 145948
rect 449250 145936 449256 145948
rect 449308 145936 449314 145988
rect 252002 145596 252008 145648
rect 252060 145636 252066 145648
rect 268470 145636 268476 145648
rect 252060 145608 268476 145636
rect 252060 145596 252066 145608
rect 268470 145596 268476 145608
rect 268528 145596 268534 145648
rect 253382 145528 253388 145580
rect 253440 145568 253446 145580
rect 307018 145568 307024 145580
rect 253440 145540 307024 145568
rect 253440 145528 253446 145540
rect 307018 145528 307024 145540
rect 307076 145528 307082 145580
rect 369118 145528 369124 145580
rect 369176 145568 369182 145580
rect 423582 145568 423588 145580
rect 369176 145540 423588 145568
rect 369176 145528 369182 145540
rect 423582 145528 423588 145540
rect 423640 145528 423646 145580
rect 456058 145528 456064 145580
rect 456116 145568 456122 145580
rect 580258 145568 580264 145580
rect 456116 145540 580264 145568
rect 456116 145528 456122 145540
rect 580258 145528 580264 145540
rect 580316 145528 580322 145580
rect 399846 145392 399852 145444
rect 399904 145432 399910 145444
rect 403526 145432 403532 145444
rect 399904 145404 403532 145432
rect 399904 145392 399910 145404
rect 403526 145392 403532 145404
rect 403584 145392 403590 145444
rect 417050 145432 417056 145444
rect 412606 145404 417056 145432
rect 359458 145052 359464 145104
rect 359516 145092 359522 145104
rect 397454 145092 397460 145104
rect 359516 145064 397460 145092
rect 359516 145052 359522 145064
rect 397454 145052 397460 145064
rect 397512 145052 397518 145104
rect 399864 145064 403848 145092
rect 171778 144984 171784 145036
rect 171836 145024 171842 145036
rect 213914 145024 213920 145036
rect 171836 144996 213920 145024
rect 171836 144984 171842 144996
rect 213914 144984 213920 144996
rect 213972 144984 213978 145036
rect 287974 144984 287980 145036
rect 288032 145024 288038 145036
rect 307478 145024 307484 145036
rect 288032 144996 307484 145024
rect 288032 144984 288038 144996
rect 307478 144984 307484 144996
rect 307536 144984 307542 145036
rect 378870 144984 378876 145036
rect 378928 145024 378934 145036
rect 399864 145024 399892 145064
rect 378928 144996 399892 145024
rect 403820 145024 403848 145064
rect 412606 145024 412634 145404
rect 417050 145392 417056 145404
rect 417108 145392 417114 145444
rect 403820 144996 412634 145024
rect 378928 144984 378934 144996
rect 166258 144916 166264 144968
rect 166316 144956 166322 144968
rect 214006 144956 214012 144968
rect 166316 144928 214012 144956
rect 166316 144916 166322 144928
rect 214006 144916 214012 144928
rect 214064 144916 214070 144968
rect 268562 144916 268568 144968
rect 268620 144956 268626 144968
rect 307662 144956 307668 144968
rect 268620 144928 307668 144956
rect 268620 144916 268626 144928
rect 307662 144916 307668 144928
rect 307720 144916 307726 144968
rect 329190 144916 329196 144968
rect 329248 144956 329254 144968
rect 399846 144956 399852 144968
rect 329248 144928 399852 144956
rect 329248 144916 329254 144928
rect 399846 144916 399852 144928
rect 399904 144916 399910 144968
rect 252186 144848 252192 144900
rect 252244 144888 252250 144900
rect 267734 144888 267740 144900
rect 252244 144860 267740 144888
rect 252244 144848 252250 144860
rect 267734 144848 267740 144860
rect 267792 144848 267798 144900
rect 324406 144848 324412 144900
rect 324464 144888 324470 144900
rect 331490 144888 331496 144900
rect 324464 144860 331496 144888
rect 324464 144848 324470 144860
rect 331490 144848 331496 144860
rect 331548 144848 331554 144900
rect 452562 144848 452568 144900
rect 452620 144888 452626 144900
rect 467098 144888 467104 144900
rect 452620 144860 467104 144888
rect 452620 144848 452626 144860
rect 467098 144848 467104 144860
rect 467156 144848 467162 144900
rect 324314 144780 324320 144832
rect 324372 144820 324378 144832
rect 328546 144820 328552 144832
rect 324372 144792 328552 144820
rect 324372 144780 324378 144792
rect 328546 144780 328552 144792
rect 328604 144780 328610 144832
rect 294690 144236 294696 144288
rect 294748 144276 294754 144288
rect 307570 144276 307576 144288
rect 294748 144248 307576 144276
rect 294748 144236 294754 144248
rect 307570 144236 307576 144248
rect 307628 144236 307634 144288
rect 373258 144236 373264 144288
rect 373316 144276 373322 144288
rect 376662 144276 376668 144288
rect 373316 144248 376668 144276
rect 373316 144236 373322 144248
rect 376662 144236 376668 144248
rect 376720 144276 376726 144288
rect 397454 144276 397460 144288
rect 376720 144248 397460 144276
rect 376720 144236 376726 144248
rect 397454 144236 397460 144248
rect 397512 144236 397518 144288
rect 264514 144168 264520 144220
rect 264572 144208 264578 144220
rect 306558 144208 306564 144220
rect 264572 144180 306564 144208
rect 264572 144168 264578 144180
rect 306558 144168 306564 144180
rect 306616 144168 306622 144220
rect 340966 144168 340972 144220
rect 341024 144208 341030 144220
rect 400490 144208 400496 144220
rect 341024 144180 400496 144208
rect 341024 144168 341030 144180
rect 400490 144168 400496 144180
rect 400548 144168 400554 144220
rect 252462 144032 252468 144084
rect 252520 144072 252526 144084
rect 258074 144072 258080 144084
rect 252520 144044 258080 144072
rect 252520 144032 252526 144044
rect 258074 144032 258080 144044
rect 258132 144032 258138 144084
rect 192570 143556 192576 143608
rect 192628 143596 192634 143608
rect 213914 143596 213920 143608
rect 192628 143568 213920 143596
rect 192628 143556 192634 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 293494 143556 293500 143608
rect 293552 143596 293558 143608
rect 307478 143596 307484 143608
rect 293552 143568 307484 143596
rect 293552 143556 293558 143568
rect 307478 143556 307484 143568
rect 307536 143556 307542 143608
rect 324958 143556 324964 143608
rect 325016 143596 325022 143608
rect 327810 143596 327816 143608
rect 325016 143568 327816 143596
rect 325016 143556 325022 143568
rect 327810 143556 327816 143568
rect 327868 143556 327874 143608
rect 252462 143488 252468 143540
rect 252520 143528 252526 143540
rect 260926 143528 260932 143540
rect 252520 143500 260932 143528
rect 252520 143488 252526 143500
rect 260926 143488 260932 143500
rect 260984 143488 260990 143540
rect 324314 143488 324320 143540
rect 324372 143528 324378 143540
rect 331398 143528 331404 143540
rect 324372 143500 331404 143528
rect 324372 143488 324378 143500
rect 331398 143488 331404 143500
rect 331456 143488 331462 143540
rect 449066 143420 449072 143472
rect 449124 143460 449130 143472
rect 449526 143460 449532 143472
rect 449124 143432 449532 143460
rect 449124 143420 449130 143432
rect 449526 143420 449532 143432
rect 449584 143420 449590 143472
rect 211798 142672 211804 142724
rect 211856 142712 211862 142724
rect 213914 142712 213920 142724
rect 211856 142684 213920 142712
rect 211856 142672 211862 142684
rect 213914 142672 213920 142684
rect 213972 142672 213978 142724
rect 251818 142672 251824 142724
rect 251876 142712 251882 142724
rect 257338 142712 257344 142724
rect 251876 142684 257344 142712
rect 251876 142672 251882 142684
rect 257338 142672 257344 142684
rect 257396 142672 257402 142724
rect 279602 142196 279608 142248
rect 279660 142236 279666 142248
rect 307478 142236 307484 142248
rect 279660 142208 307484 142236
rect 279660 142196 279666 142208
rect 307478 142196 307484 142208
rect 307536 142196 307542 142248
rect 189718 142128 189724 142180
rect 189776 142168 189782 142180
rect 213914 142168 213920 142180
rect 189776 142140 213920 142168
rect 189776 142128 189782 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 255958 142128 255964 142180
rect 256016 142168 256022 142180
rect 307662 142168 307668 142180
rect 256016 142140 307668 142168
rect 256016 142128 256022 142140
rect 307662 142128 307668 142140
rect 307720 142128 307726 142180
rect 331950 142128 331956 142180
rect 332008 142168 332014 142180
rect 397546 142168 397552 142180
rect 332008 142140 397552 142168
rect 332008 142128 332014 142140
rect 397546 142128 397552 142140
rect 397604 142128 397610 142180
rect 452470 142128 452476 142180
rect 452528 142168 452534 142180
rect 498838 142168 498844 142180
rect 452528 142140 498844 142168
rect 452528 142128 452534 142140
rect 498838 142128 498844 142140
rect 498896 142128 498902 142180
rect 251726 142060 251732 142112
rect 251784 142100 251790 142112
rect 259454 142100 259460 142112
rect 251784 142072 259460 142100
rect 251784 142060 251790 142072
rect 259454 142060 259460 142072
rect 259512 142060 259518 142112
rect 324406 142060 324412 142112
rect 324464 142100 324470 142112
rect 332778 142100 332784 142112
rect 324464 142072 332784 142100
rect 324464 142060 324470 142072
rect 332778 142060 332784 142072
rect 332836 142060 332842 142112
rect 365162 142060 365168 142112
rect 365220 142100 365226 142112
rect 397454 142100 397460 142112
rect 365220 142072 397460 142100
rect 365220 142060 365226 142072
rect 397454 142060 397460 142072
rect 397512 142060 397518 142112
rect 324314 141788 324320 141840
rect 324372 141828 324378 141840
rect 327258 141828 327264 141840
rect 324372 141800 327264 141828
rect 324372 141788 324378 141800
rect 327258 141788 327264 141800
rect 327316 141788 327322 141840
rect 252370 141380 252376 141432
rect 252428 141420 252434 141432
rect 264238 141420 264244 141432
rect 252428 141392 264244 141420
rect 252428 141380 252434 141392
rect 264238 141380 264244 141392
rect 264296 141380 264302 141432
rect 301682 140904 301688 140956
rect 301740 140944 301746 140956
rect 307662 140944 307668 140956
rect 301740 140916 307668 140944
rect 301740 140904 301746 140916
rect 307662 140904 307668 140916
rect 307720 140904 307726 140956
rect 206370 140836 206376 140888
rect 206428 140876 206434 140888
rect 213914 140876 213920 140888
rect 206428 140848 213920 140876
rect 206428 140836 206434 140848
rect 213914 140836 213920 140848
rect 213972 140836 213978 140888
rect 290550 140836 290556 140888
rect 290608 140876 290614 140888
rect 307570 140876 307576 140888
rect 290608 140848 307576 140876
rect 290608 140836 290614 140848
rect 307570 140836 307576 140848
rect 307628 140836 307634 140888
rect 196618 140768 196624 140820
rect 196676 140808 196682 140820
rect 214006 140808 214012 140820
rect 196676 140780 214012 140808
rect 196676 140768 196682 140780
rect 214006 140768 214012 140780
rect 214064 140768 214070 140820
rect 257614 140768 257620 140820
rect 257672 140808 257678 140820
rect 307662 140808 307668 140820
rect 257672 140780 307668 140808
rect 257672 140768 257678 140780
rect 307662 140768 307668 140780
rect 307720 140768 307726 140820
rect 343818 140768 343824 140820
rect 343876 140808 343882 140820
rect 346394 140808 346400 140820
rect 343876 140780 346400 140808
rect 343876 140768 343882 140780
rect 346394 140768 346400 140780
rect 346452 140768 346458 140820
rect 324314 140700 324320 140752
rect 324372 140740 324378 140752
rect 337470 140740 337476 140752
rect 324372 140712 337476 140740
rect 324372 140700 324378 140712
rect 337470 140700 337476 140712
rect 337528 140700 337534 140752
rect 451918 140428 451924 140480
rect 451976 140468 451982 140480
rect 455598 140468 455604 140480
rect 451976 140440 455604 140468
rect 451976 140428 451982 140440
rect 455598 140428 455604 140440
rect 455656 140428 455662 140480
rect 194502 140020 194508 140072
rect 194560 140060 194566 140072
rect 215938 140060 215944 140072
rect 194560 140032 215944 140060
rect 194560 140020 194566 140032
rect 215938 140020 215944 140032
rect 215996 140020 216002 140072
rect 335630 140020 335636 140072
rect 335688 140060 335694 140072
rect 376662 140060 376668 140072
rect 335688 140032 376668 140060
rect 335688 140020 335694 140032
rect 376662 140020 376668 140032
rect 376720 140020 376726 140072
rect 286318 139544 286324 139596
rect 286376 139584 286382 139596
rect 306558 139584 306564 139596
rect 286376 139556 306564 139584
rect 286376 139544 286382 139556
rect 306558 139544 306564 139556
rect 306616 139544 306622 139596
rect 251726 139476 251732 139528
rect 251784 139516 251790 139528
rect 255590 139516 255596 139528
rect 251784 139488 255596 139516
rect 251784 139476 251790 139488
rect 255590 139476 255596 139488
rect 255648 139476 255654 139528
rect 256050 139476 256056 139528
rect 256108 139516 256114 139528
rect 307570 139516 307576 139528
rect 256108 139488 307576 139516
rect 256108 139476 256114 139488
rect 307570 139476 307576 139488
rect 307628 139476 307634 139528
rect 182910 139408 182916 139460
rect 182968 139448 182974 139460
rect 213914 139448 213920 139460
rect 182968 139420 213920 139448
rect 182968 139408 182974 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 250530 139408 250536 139460
rect 250588 139448 250594 139460
rect 307662 139448 307668 139460
rect 250588 139420 307668 139448
rect 250588 139408 250594 139420
rect 307662 139408 307668 139420
rect 307720 139408 307726 139460
rect 251726 139340 251732 139392
rect 251784 139380 251790 139392
rect 280154 139380 280160 139392
rect 251784 139352 280160 139380
rect 251784 139340 251790 139352
rect 280154 139340 280160 139352
rect 280212 139340 280218 139392
rect 354030 139340 354036 139392
rect 354088 139380 354094 139392
rect 354674 139380 354680 139392
rect 354088 139352 354680 139380
rect 354088 139340 354094 139352
rect 354674 139340 354680 139352
rect 354732 139380 354738 139392
rect 397454 139380 397460 139392
rect 354732 139352 397460 139380
rect 354732 139340 354738 139352
rect 397454 139340 397460 139352
rect 397512 139340 397518 139392
rect 252462 139272 252468 139324
rect 252520 139312 252526 139324
rect 260834 139312 260840 139324
rect 252520 139284 260840 139312
rect 252520 139272 252526 139284
rect 260834 139272 260840 139284
rect 260892 139272 260898 139324
rect 324314 139272 324320 139324
rect 324372 139312 324378 139324
rect 354858 139312 354864 139324
rect 324372 139284 354864 139312
rect 324372 139272 324378 139284
rect 354858 139272 354864 139284
rect 354916 139272 354922 139324
rect 452102 138864 452108 138916
rect 452160 138904 452166 138916
rect 458358 138904 458364 138916
rect 452160 138876 458364 138904
rect 452160 138864 452166 138876
rect 458358 138864 458364 138876
rect 458416 138864 458422 138916
rect 282270 138116 282276 138168
rect 282328 138156 282334 138168
rect 307662 138156 307668 138168
rect 282328 138128 307668 138156
rect 282328 138116 282334 138128
rect 307662 138116 307668 138128
rect 307720 138116 307726 138168
rect 253198 138048 253204 138100
rect 253256 138088 253262 138100
rect 307478 138088 307484 138100
rect 253256 138060 307484 138088
rect 253256 138048 253262 138060
rect 307478 138048 307484 138060
rect 307536 138048 307542 138100
rect 193950 137980 193956 138032
rect 194008 138020 194014 138032
rect 213914 138020 213920 138032
rect 194008 137992 213920 138020
rect 194008 137980 194014 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 250438 137980 250444 138032
rect 250496 138020 250502 138032
rect 307570 138020 307576 138032
rect 250496 137992 307576 138020
rect 250496 137980 250502 137992
rect 307570 137980 307576 137992
rect 307628 137980 307634 138032
rect 252462 137912 252468 137964
rect 252520 137952 252526 137964
rect 281534 137952 281540 137964
rect 252520 137924 281540 137952
rect 252520 137912 252526 137924
rect 281534 137912 281540 137924
rect 281592 137912 281598 137964
rect 324314 137912 324320 137964
rect 324372 137952 324378 137964
rect 347958 137952 347964 137964
rect 324372 137924 347964 137952
rect 324372 137912 324378 137924
rect 347958 137912 347964 137924
rect 348016 137912 348022 137964
rect 360102 137912 360108 137964
rect 360160 137952 360166 137964
rect 397546 137952 397552 137964
rect 360160 137924 397552 137952
rect 360160 137912 360166 137924
rect 397546 137912 397552 137924
rect 397604 137912 397610 137964
rect 251358 137844 251364 137896
rect 251416 137884 251422 137896
rect 269114 137884 269120 137896
rect 251416 137856 269120 137884
rect 251416 137844 251422 137856
rect 269114 137844 269120 137856
rect 269172 137844 269178 137896
rect 322934 137844 322940 137896
rect 322992 137884 322998 137896
rect 323302 137884 323308 137896
rect 322992 137856 323308 137884
rect 322992 137844 322998 137856
rect 323302 137844 323308 137856
rect 323360 137884 323366 137896
rect 330478 137884 330484 137896
rect 323360 137856 330484 137884
rect 323360 137844 323366 137856
rect 330478 137844 330484 137856
rect 330536 137844 330542 137896
rect 391842 137844 391848 137896
rect 391900 137884 391906 137896
rect 397454 137884 397460 137896
rect 391900 137856 397460 137884
rect 391900 137844 391906 137856
rect 397454 137844 397460 137856
rect 397512 137844 397518 137896
rect 256234 137232 256240 137284
rect 256292 137272 256298 137284
rect 307110 137272 307116 137284
rect 256292 137244 307116 137272
rect 256292 137232 256298 137244
rect 307110 137232 307116 137244
rect 307168 137232 307174 137284
rect 210510 136688 210516 136740
rect 210568 136728 210574 136740
rect 213914 136728 213920 136740
rect 210568 136700 213920 136728
rect 210568 136688 210574 136700
rect 213914 136688 213920 136700
rect 213972 136688 213978 136740
rect 293310 136688 293316 136740
rect 293368 136728 293374 136740
rect 306742 136728 306748 136740
rect 293368 136700 306748 136728
rect 293368 136688 293374 136700
rect 306742 136688 306748 136700
rect 306800 136688 306806 136740
rect 171870 136620 171876 136672
rect 171928 136660 171934 136672
rect 214098 136660 214104 136672
rect 171928 136632 214104 136660
rect 171928 136620 171934 136632
rect 214098 136620 214104 136632
rect 214156 136620 214162 136672
rect 276750 136620 276756 136672
rect 276808 136660 276814 136672
rect 307662 136660 307668 136672
rect 276808 136632 307668 136660
rect 276808 136620 276814 136632
rect 307662 136620 307668 136632
rect 307720 136620 307726 136672
rect 252462 136552 252468 136604
rect 252520 136592 252526 136604
rect 287698 136592 287704 136604
rect 252520 136564 287704 136592
rect 252520 136552 252526 136564
rect 287698 136552 287704 136564
rect 287756 136552 287762 136604
rect 323394 136552 323400 136604
rect 323452 136592 323458 136604
rect 343818 136592 343824 136604
rect 323452 136564 343824 136592
rect 323452 136552 323458 136564
rect 343818 136552 343824 136564
rect 343876 136552 343882 136604
rect 251726 136484 251732 136536
rect 251784 136524 251790 136536
rect 279418 136524 279424 136536
rect 251784 136496 279424 136524
rect 251784 136484 251790 136496
rect 279418 136484 279424 136496
rect 279476 136484 279482 136536
rect 324314 136484 324320 136536
rect 324372 136524 324378 136536
rect 342438 136524 342444 136536
rect 324372 136496 342444 136524
rect 324372 136484 324378 136496
rect 342438 136484 342444 136496
rect 342496 136484 342502 136536
rect 300210 135464 300216 135516
rect 300268 135504 300274 135516
rect 307662 135504 307668 135516
rect 300268 135476 307668 135504
rect 300268 135464 300274 135476
rect 307662 135464 307668 135476
rect 307720 135464 307726 135516
rect 207750 135396 207756 135448
rect 207808 135436 207814 135448
rect 214006 135436 214012 135448
rect 207808 135408 214012 135436
rect 207808 135396 207814 135408
rect 214006 135396 214012 135408
rect 214064 135396 214070 135448
rect 298738 135396 298744 135448
rect 298796 135436 298802 135448
rect 306926 135436 306932 135448
rect 298796 135408 306932 135436
rect 298796 135396 298802 135408
rect 306926 135396 306932 135408
rect 306984 135396 306990 135448
rect 202230 135328 202236 135380
rect 202288 135368 202294 135380
rect 213914 135368 213920 135380
rect 202288 135340 213920 135368
rect 202288 135328 202294 135340
rect 213914 135328 213920 135340
rect 213972 135328 213978 135380
rect 280798 135328 280804 135380
rect 280856 135368 280862 135380
rect 306558 135368 306564 135380
rect 280856 135340 306564 135368
rect 280856 135328 280862 135340
rect 306558 135328 306564 135340
rect 306616 135328 306622 135380
rect 181438 135260 181444 135312
rect 181496 135300 181502 135312
rect 214098 135300 214104 135312
rect 181496 135272 214104 135300
rect 181496 135260 181502 135272
rect 214098 135260 214104 135272
rect 214156 135260 214162 135312
rect 266998 135260 267004 135312
rect 267056 135300 267062 135312
rect 306742 135300 306748 135312
rect 267056 135272 306748 135300
rect 267056 135260 267062 135272
rect 306742 135260 306748 135272
rect 306800 135260 306806 135312
rect 390186 135260 390192 135312
rect 390244 135300 390250 135312
rect 391934 135300 391940 135312
rect 390244 135272 391940 135300
rect 390244 135260 390250 135272
rect 391934 135260 391940 135272
rect 391992 135300 391998 135312
rect 397454 135300 397460 135312
rect 391992 135272 397460 135300
rect 391992 135260 391998 135272
rect 397454 135260 397460 135272
rect 397512 135260 397518 135312
rect 251450 135192 251456 135244
rect 251508 135232 251514 135244
rect 287790 135232 287796 135244
rect 251508 135204 287796 135232
rect 251508 135192 251514 135204
rect 287790 135192 287796 135204
rect 287848 135192 287854 135244
rect 324406 135192 324412 135244
rect 324464 135232 324470 135244
rect 335446 135232 335452 135244
rect 324464 135204 335452 135232
rect 324464 135192 324470 135204
rect 335446 135192 335452 135204
rect 335504 135192 335510 135244
rect 451918 135192 451924 135244
rect 451976 135232 451982 135244
rect 454310 135232 454316 135244
rect 451976 135204 454316 135232
rect 451976 135192 451982 135204
rect 454310 135192 454316 135204
rect 454368 135192 454374 135244
rect 252462 135124 252468 135176
rect 252520 135164 252526 135176
rect 271230 135164 271236 135176
rect 252520 135136 271236 135164
rect 252520 135124 252526 135136
rect 271230 135124 271236 135136
rect 271288 135124 271294 135176
rect 324314 135124 324320 135176
rect 324372 135164 324378 135176
rect 332686 135164 332692 135176
rect 324372 135136 332692 135164
rect 324372 135124 324378 135136
rect 332686 135124 332692 135136
rect 332744 135124 332750 135176
rect 394050 134648 394056 134700
rect 394108 134688 394114 134700
rect 396074 134688 396080 134700
rect 394108 134660 396080 134688
rect 394108 134648 394114 134660
rect 396074 134648 396080 134660
rect 396132 134688 396138 134700
rect 397454 134688 397460 134700
rect 396132 134660 397460 134688
rect 396132 134648 396138 134660
rect 397454 134648 397460 134660
rect 397512 134648 397518 134700
rect 327074 134512 327080 134564
rect 327132 134552 327138 134564
rect 367094 134552 367100 134564
rect 327132 134524 367100 134552
rect 327132 134512 327138 134524
rect 367094 134512 367100 134524
rect 367152 134512 367158 134564
rect 387150 134512 387156 134564
rect 387208 134552 387214 134564
rect 399018 134552 399024 134564
rect 387208 134524 399024 134552
rect 387208 134512 387214 134524
rect 399018 134512 399024 134524
rect 399076 134512 399082 134564
rect 296070 134036 296076 134088
rect 296128 134076 296134 134088
rect 307662 134076 307668 134088
rect 296128 134048 307668 134076
rect 296128 134036 296134 134048
rect 307662 134036 307668 134048
rect 307720 134036 307726 134088
rect 174630 133968 174636 134020
rect 174688 134008 174694 134020
rect 214006 134008 214012 134020
rect 174688 133980 214012 134008
rect 174688 133968 174694 133980
rect 214006 133968 214012 133980
rect 214064 133968 214070 134020
rect 290458 133968 290464 134020
rect 290516 134008 290522 134020
rect 307478 134008 307484 134020
rect 290516 133980 307484 134008
rect 290516 133968 290522 133980
rect 307478 133968 307484 133980
rect 307536 133968 307542 134020
rect 170398 133900 170404 133952
rect 170456 133940 170462 133952
rect 213914 133940 213920 133952
rect 170456 133912 213920 133940
rect 170456 133900 170462 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 289262 133900 289268 133952
rect 289320 133940 289326 133952
rect 307570 133940 307576 133952
rect 289320 133912 307576 133940
rect 289320 133900 289326 133912
rect 307570 133900 307576 133912
rect 307628 133900 307634 133952
rect 251358 133832 251364 133884
rect 251416 133872 251422 133884
rect 290642 133872 290648 133884
rect 251416 133844 290648 133872
rect 251416 133832 251422 133844
rect 290642 133832 290648 133844
rect 290700 133832 290706 133884
rect 324314 133832 324320 133884
rect 324372 133872 324378 133884
rect 357526 133872 357532 133884
rect 324372 133844 357532 133872
rect 324372 133832 324378 133844
rect 357526 133832 357532 133844
rect 357584 133832 357590 133884
rect 452194 133832 452200 133884
rect 452252 133872 452258 133884
rect 482278 133872 482284 133884
rect 452252 133844 482284 133872
rect 452252 133832 452258 133844
rect 482278 133832 482284 133844
rect 482336 133832 482342 133884
rect 252370 133764 252376 133816
rect 252428 133804 252434 133816
rect 282362 133804 282368 133816
rect 252428 133776 282368 133804
rect 252428 133764 252434 133776
rect 282362 133764 282368 133776
rect 282420 133764 282426 133816
rect 252462 133696 252468 133748
rect 252520 133736 252526 133748
rect 269942 133736 269948 133748
rect 252520 133708 269948 133736
rect 252520 133696 252526 133708
rect 269942 133696 269948 133708
rect 270000 133696 270006 133748
rect 321646 133152 321652 133204
rect 321704 133192 321710 133204
rect 357434 133192 357440 133204
rect 321704 133164 357440 133192
rect 321704 133152 321710 133164
rect 357434 133152 357440 133164
rect 357492 133152 357498 133204
rect 297450 132608 297456 132660
rect 297508 132648 297514 132660
rect 307662 132648 307668 132660
rect 297508 132620 307668 132648
rect 297508 132608 297514 132620
rect 307662 132608 307668 132620
rect 307720 132608 307726 132660
rect 207658 132540 207664 132592
rect 207716 132580 207722 132592
rect 214006 132580 214012 132592
rect 207716 132552 214012 132580
rect 207716 132540 207722 132552
rect 214006 132540 214012 132552
rect 214064 132540 214070 132592
rect 282454 132540 282460 132592
rect 282512 132580 282518 132592
rect 307478 132580 307484 132592
rect 282512 132552 307484 132580
rect 282512 132540 282518 132552
rect 307478 132540 307484 132552
rect 307536 132540 307542 132592
rect 391290 132540 391296 132592
rect 391348 132580 391354 132592
rect 394602 132580 394608 132592
rect 391348 132552 394608 132580
rect 391348 132540 391354 132552
rect 394602 132540 394608 132552
rect 394660 132580 394666 132592
rect 397546 132580 397552 132592
rect 394660 132552 397552 132580
rect 394660 132540 394666 132552
rect 397546 132540 397552 132552
rect 397604 132540 397610 132592
rect 173158 132472 173164 132524
rect 173216 132512 173222 132524
rect 213914 132512 213920 132524
rect 173216 132484 213920 132512
rect 173216 132472 173222 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 269850 132472 269856 132524
rect 269908 132512 269914 132524
rect 307570 132512 307576 132524
rect 269908 132484 307576 132512
rect 269908 132472 269914 132484
rect 307570 132472 307576 132484
rect 307628 132472 307634 132524
rect 392578 132472 392584 132524
rect 392636 132512 392642 132524
rect 397454 132512 397460 132524
rect 392636 132484 397460 132512
rect 392636 132472 392642 132484
rect 397454 132472 397460 132484
rect 397512 132472 397518 132524
rect 252462 132404 252468 132456
rect 252520 132444 252526 132456
rect 300118 132444 300124 132456
rect 252520 132416 300124 132444
rect 252520 132404 252526 132416
rect 300118 132404 300124 132416
rect 300176 132404 300182 132456
rect 449986 132404 449992 132456
rect 450044 132444 450050 132456
rect 472618 132444 472624 132456
rect 450044 132416 472624 132444
rect 450044 132404 450050 132416
rect 472618 132404 472624 132416
rect 472676 132404 472682 132456
rect 251542 132336 251548 132388
rect 251600 132376 251606 132388
rect 265618 132376 265624 132388
rect 251600 132348 265624 132376
rect 251600 132336 251606 132348
rect 265618 132336 265624 132348
rect 265676 132336 265682 132388
rect 252002 131792 252008 131844
rect 252060 131832 252066 131844
rect 279510 131832 279516 131844
rect 252060 131804 279516 131832
rect 252060 131792 252066 131804
rect 279510 131792 279516 131804
rect 279568 131792 279574 131844
rect 265710 131724 265716 131776
rect 265768 131764 265774 131776
rect 301498 131764 301504 131776
rect 265768 131736 301504 131764
rect 265768 131724 265774 131736
rect 301498 131724 301504 131736
rect 301556 131724 301562 131776
rect 337470 131724 337476 131776
rect 337528 131764 337534 131776
rect 398742 131764 398748 131776
rect 337528 131736 398748 131764
rect 337528 131724 337534 131736
rect 398742 131724 398748 131736
rect 398800 131724 398806 131776
rect 303062 131248 303068 131300
rect 303120 131288 303126 131300
rect 307478 131288 307484 131300
rect 303120 131260 307484 131288
rect 303120 131248 303126 131260
rect 307478 131248 307484 131260
rect 307536 131248 307542 131300
rect 287698 131180 287704 131232
rect 287756 131220 287762 131232
rect 307570 131220 307576 131232
rect 287756 131192 307576 131220
rect 287756 131180 287762 131192
rect 307570 131180 307576 131192
rect 307628 131180 307634 131232
rect 264422 131112 264428 131164
rect 264480 131152 264486 131164
rect 307662 131152 307668 131164
rect 264480 131124 307668 131152
rect 264480 131112 264486 131124
rect 307662 131112 307668 131124
rect 307720 131112 307726 131164
rect 252370 131044 252376 131096
rect 252428 131084 252434 131096
rect 304258 131084 304264 131096
rect 252428 131056 304264 131084
rect 252428 131044 252434 131056
rect 304258 131044 304264 131056
rect 304316 131044 304322 131096
rect 324406 131044 324412 131096
rect 324464 131084 324470 131096
rect 356238 131084 356244 131096
rect 324464 131056 356244 131084
rect 324464 131044 324470 131056
rect 356238 131044 356244 131056
rect 356296 131084 356302 131096
rect 360838 131084 360844 131096
rect 356296 131056 360844 131084
rect 356296 131044 356302 131056
rect 360838 131044 360844 131056
rect 360896 131044 360902 131096
rect 252462 130976 252468 131028
rect 252520 131016 252526 131028
rect 274082 131016 274088 131028
rect 252520 130988 274088 131016
rect 252520 130976 252526 130988
rect 274082 130976 274088 130988
rect 274140 130976 274146 131028
rect 324314 130976 324320 131028
rect 324372 131016 324378 131028
rect 339586 131016 339592 131028
rect 324372 130988 339592 131016
rect 324372 130976 324378 130988
rect 339586 130976 339592 130988
rect 339644 130976 339650 131028
rect 252462 130500 252468 130552
rect 252520 130540 252526 130552
rect 257522 130540 257528 130552
rect 252520 130512 257528 130540
rect 252520 130500 252526 130512
rect 257522 130500 257528 130512
rect 257580 130500 257586 130552
rect 449158 130024 449164 130076
rect 449216 130064 449222 130076
rect 449434 130064 449440 130076
rect 449216 130036 449440 130064
rect 449216 130024 449222 130036
rect 449434 130024 449440 130036
rect 449492 130024 449498 130076
rect 257338 129956 257344 130008
rect 257396 129996 257402 130008
rect 307570 129996 307576 130008
rect 257396 129968 307576 129996
rect 257396 129956 257402 129968
rect 307570 129956 307576 129968
rect 307628 129956 307634 130008
rect 292022 129888 292028 129940
rect 292080 129928 292086 129940
rect 307662 129928 307668 129940
rect 292080 129900 307668 129928
rect 292080 129888 292086 129900
rect 307662 129888 307668 129900
rect 307720 129888 307726 129940
rect 273990 129820 273996 129872
rect 274048 129860 274054 129872
rect 307478 129860 307484 129872
rect 274048 129832 307484 129860
rect 274048 129820 274054 129832
rect 307478 129820 307484 129832
rect 307536 129820 307542 129872
rect 395890 129820 395896 129872
rect 395948 129860 395954 129872
rect 398282 129860 398288 129872
rect 395948 129832 398288 129860
rect 395948 129820 395954 129832
rect 398282 129820 398288 129832
rect 398340 129820 398346 129872
rect 184198 129752 184204 129804
rect 184256 129792 184262 129804
rect 213914 129792 213920 129804
rect 184256 129764 213920 129792
rect 184256 129752 184262 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 304350 129752 304356 129804
rect 304408 129792 304414 129804
rect 307110 129792 307116 129804
rect 304408 129764 307116 129792
rect 304408 129752 304414 129764
rect 307110 129752 307116 129764
rect 307168 129752 307174 129804
rect 360930 129752 360936 129804
rect 360988 129792 360994 129804
rect 397546 129792 397552 129804
rect 360988 129764 397552 129792
rect 360988 129752 360994 129764
rect 397546 129752 397552 129764
rect 397604 129752 397610 129804
rect 252462 129684 252468 129736
rect 252520 129724 252526 129736
rect 284938 129724 284944 129736
rect 252520 129696 284944 129724
rect 252520 129684 252526 129696
rect 284938 129684 284944 129696
rect 284996 129684 285002 129736
rect 324406 129684 324412 129736
rect 324464 129724 324470 129736
rect 343726 129724 343732 129736
rect 324464 129696 343732 129724
rect 324464 129684 324470 129696
rect 343726 129684 343732 129696
rect 343784 129724 343790 129736
rect 362218 129724 362224 129736
rect 343784 129696 362224 129724
rect 343784 129684 343790 129696
rect 362218 129684 362224 129696
rect 362276 129684 362282 129736
rect 385678 129684 385684 129736
rect 385736 129724 385742 129736
rect 397454 129724 397460 129736
rect 385736 129696 397460 129724
rect 385736 129684 385742 129696
rect 397454 129684 397460 129696
rect 397512 129684 397518 129736
rect 452562 129684 452568 129736
rect 452620 129724 452626 129736
rect 465074 129724 465080 129736
rect 452620 129696 465080 129724
rect 452620 129684 452626 129696
rect 465074 129684 465080 129696
rect 465132 129684 465138 129736
rect 251450 129616 251456 129668
rect 251508 129656 251514 129668
rect 268378 129656 268384 129668
rect 251508 129628 268384 129656
rect 251508 129616 251514 129628
rect 268378 129616 268384 129628
rect 268436 129616 268442 129668
rect 252370 129548 252376 129600
rect 252428 129588 252434 129600
rect 267090 129588 267096 129600
rect 252428 129560 267096 129588
rect 252428 129548 252434 129560
rect 267090 129548 267096 129560
rect 267148 129548 267154 129600
rect 324314 129412 324320 129464
rect 324372 129452 324378 129464
rect 327074 129452 327080 129464
rect 324372 129424 327080 129452
rect 324372 129412 324378 129424
rect 327074 129412 327080 129424
rect 327132 129412 327138 129464
rect 285030 128392 285036 128444
rect 285088 128432 285094 128444
rect 306558 128432 306564 128444
rect 285088 128404 306564 128432
rect 285088 128392 285094 128404
rect 306558 128392 306564 128404
rect 306616 128392 306622 128444
rect 186958 128324 186964 128376
rect 187016 128364 187022 128376
rect 213914 128364 213920 128376
rect 187016 128336 213920 128364
rect 187016 128324 187022 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 268470 128324 268476 128376
rect 268528 128364 268534 128376
rect 307110 128364 307116 128376
rect 268528 128336 307116 128364
rect 268528 128324 268534 128336
rect 307110 128324 307116 128336
rect 307168 128324 307174 128376
rect 251634 128256 251640 128308
rect 251692 128296 251698 128308
rect 295978 128296 295984 128308
rect 251692 128268 295984 128296
rect 251692 128256 251698 128268
rect 295978 128256 295984 128268
rect 296036 128256 296042 128308
rect 324314 128256 324320 128308
rect 324372 128296 324378 128308
rect 349338 128296 349344 128308
rect 324372 128268 349344 128296
rect 324372 128256 324378 128268
rect 349338 128256 349344 128268
rect 349396 128296 349402 128308
rect 392670 128296 392676 128308
rect 349396 128268 392676 128296
rect 349396 128256 349402 128268
rect 392670 128256 392676 128268
rect 392728 128256 392734 128308
rect 452102 128256 452108 128308
rect 452160 128296 452166 128308
rect 458266 128296 458272 128308
rect 452160 128268 458272 128296
rect 452160 128256 452166 128268
rect 458266 128256 458272 128268
rect 458324 128256 458330 128308
rect 252462 128188 252468 128240
rect 252520 128228 252526 128240
rect 264330 128228 264336 128240
rect 252520 128200 264336 128228
rect 252520 128188 252526 128200
rect 264330 128188 264336 128200
rect 264388 128188 264394 128240
rect 324406 128188 324412 128240
rect 324464 128228 324470 128240
rect 329834 128228 329840 128240
rect 324464 128200 329840 128228
rect 324464 128188 324470 128200
rect 329834 128188 329840 128200
rect 329892 128188 329898 128240
rect 385678 127576 385684 127628
rect 385736 127616 385742 127628
rect 397454 127616 397460 127628
rect 385736 127588 397460 127616
rect 385736 127576 385742 127588
rect 397454 127576 397460 127588
rect 397512 127576 397518 127628
rect 252186 127440 252192 127492
rect 252244 127480 252250 127492
rect 257706 127480 257712 127492
rect 252244 127452 257712 127480
rect 252244 127440 252250 127452
rect 257706 127440 257712 127452
rect 257764 127440 257770 127492
rect 297542 127100 297548 127152
rect 297600 127140 297606 127152
rect 307110 127140 307116 127152
rect 297600 127112 307116 127140
rect 297600 127100 297606 127112
rect 307110 127100 307116 127112
rect 307168 127100 307174 127152
rect 264238 127032 264244 127084
rect 264296 127072 264302 127084
rect 307662 127072 307668 127084
rect 264296 127044 307668 127072
rect 264296 127032 264302 127044
rect 307662 127032 307668 127044
rect 307720 127032 307726 127084
rect 170490 126964 170496 127016
rect 170548 127004 170554 127016
rect 213914 127004 213920 127016
rect 170548 126976 213920 127004
rect 170548 126964 170554 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 260190 126964 260196 127016
rect 260248 127004 260254 127016
rect 306742 127004 306748 127016
rect 260248 126976 306748 127004
rect 260248 126964 260254 126976
rect 306742 126964 306748 126976
rect 306800 126964 306806 127016
rect 252462 126896 252468 126948
rect 252520 126936 252526 126948
rect 293218 126936 293224 126948
rect 252520 126908 293224 126936
rect 252520 126896 252526 126908
rect 293218 126896 293224 126908
rect 293276 126896 293282 126948
rect 342990 126896 342996 126948
rect 343048 126936 343054 126948
rect 343634 126936 343640 126948
rect 343048 126908 343640 126936
rect 343048 126896 343054 126908
rect 343634 126896 343640 126908
rect 343692 126936 343698 126948
rect 397546 126936 397552 126948
rect 343692 126908 397552 126936
rect 343692 126896 343698 126908
rect 397546 126896 397552 126908
rect 397604 126896 397610 126948
rect 452562 126896 452568 126948
rect 452620 126936 452626 126948
rect 476206 126936 476212 126948
rect 452620 126908 476212 126936
rect 452620 126896 452626 126908
rect 476206 126896 476212 126908
rect 476264 126896 476270 126948
rect 252094 126828 252100 126880
rect 252152 126868 252158 126880
rect 275370 126868 275376 126880
rect 252152 126840 275376 126868
rect 252152 126828 252158 126840
rect 275370 126828 275376 126840
rect 275428 126828 275434 126880
rect 377950 126828 377956 126880
rect 378008 126868 378014 126880
rect 397454 126868 397460 126880
rect 378008 126840 397460 126868
rect 378008 126828 378014 126840
rect 397454 126828 397460 126840
rect 397512 126828 397518 126880
rect 251358 126216 251364 126268
rect 251416 126256 251422 126268
rect 300302 126256 300308 126268
rect 251416 126228 300308 126256
rect 251416 126216 251422 126228
rect 300302 126216 300308 126228
rect 300360 126216 300366 126268
rect 203610 125672 203616 125724
rect 203668 125712 203674 125724
rect 213914 125712 213920 125724
rect 203668 125684 213920 125712
rect 203668 125672 203674 125684
rect 213914 125672 213920 125684
rect 213972 125672 213978 125724
rect 284938 125672 284944 125724
rect 284996 125712 285002 125724
rect 307662 125712 307668 125724
rect 284996 125684 307668 125712
rect 284996 125672 285002 125684
rect 307662 125672 307668 125684
rect 307720 125672 307726 125724
rect 200758 125604 200764 125656
rect 200816 125644 200822 125656
rect 214006 125644 214012 125656
rect 200816 125616 214012 125644
rect 200816 125604 200822 125616
rect 214006 125604 214012 125616
rect 214064 125604 214070 125656
rect 275278 125604 275284 125656
rect 275336 125644 275342 125656
rect 306742 125644 306748 125656
rect 275336 125616 306748 125644
rect 275336 125604 275342 125616
rect 306742 125604 306748 125616
rect 306800 125604 306806 125656
rect 324314 125536 324320 125588
rect 324372 125576 324378 125588
rect 347866 125576 347872 125588
rect 324372 125548 347872 125576
rect 324372 125536 324378 125548
rect 347866 125536 347872 125548
rect 347924 125536 347930 125588
rect 353938 125536 353944 125588
rect 353996 125576 354002 125588
rect 397454 125576 397460 125588
rect 353996 125548 397460 125576
rect 353996 125536 354002 125548
rect 397454 125536 397460 125548
rect 397512 125536 397518 125588
rect 452562 125536 452568 125588
rect 452620 125576 452626 125588
rect 464338 125576 464344 125588
rect 452620 125548 464344 125576
rect 452620 125536 452626 125548
rect 464338 125536 464344 125548
rect 464396 125536 464402 125588
rect 251910 125332 251916 125384
rect 251968 125372 251974 125384
rect 256234 125372 256240 125384
rect 251968 125344 256240 125372
rect 251968 125332 251974 125344
rect 256234 125332 256240 125344
rect 256292 125332 256298 125384
rect 252462 124992 252468 125044
rect 252520 125032 252526 125044
rect 258902 125032 258908 125044
rect 252520 125004 258908 125032
rect 252520 124992 252526 125004
rect 258902 124992 258908 125004
rect 258960 124992 258966 125044
rect 252278 124856 252284 124908
rect 252336 124896 252342 124908
rect 302970 124896 302976 124908
rect 252336 124868 302976 124896
rect 252336 124856 252342 124868
rect 302970 124856 302976 124868
rect 303028 124856 303034 124908
rect 451274 124720 451280 124772
rect 451332 124760 451338 124772
rect 454218 124760 454224 124772
rect 451332 124732 454224 124760
rect 451332 124720 451338 124732
rect 454218 124720 454224 124732
rect 454276 124720 454282 124772
rect 302878 124312 302884 124364
rect 302936 124352 302942 124364
rect 307662 124352 307668 124364
rect 302936 124324 307668 124352
rect 302936 124312 302942 124324
rect 307662 124312 307668 124324
rect 307720 124312 307726 124364
rect 171962 124244 171968 124296
rect 172020 124284 172026 124296
rect 214006 124284 214012 124296
rect 172020 124256 214012 124284
rect 172020 124244 172026 124256
rect 214006 124244 214012 124256
rect 214064 124244 214070 124296
rect 291930 124244 291936 124296
rect 291988 124284 291994 124296
rect 306742 124284 306748 124296
rect 291988 124256 306748 124284
rect 291988 124244 291994 124256
rect 306742 124244 306748 124256
rect 306800 124244 306806 124296
rect 167638 124176 167644 124228
rect 167696 124216 167702 124228
rect 213914 124216 213920 124228
rect 167696 124188 213920 124216
rect 167696 124176 167702 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 258718 124176 258724 124228
rect 258776 124216 258782 124228
rect 307110 124216 307116 124228
rect 258776 124188 307116 124216
rect 258776 124176 258782 124188
rect 307110 124176 307116 124188
rect 307168 124176 307174 124228
rect 252370 124108 252376 124160
rect 252428 124148 252434 124160
rect 283558 124148 283564 124160
rect 252428 124120 283564 124148
rect 252428 124108 252434 124120
rect 283558 124108 283564 124120
rect 283616 124108 283622 124160
rect 252462 124040 252468 124092
rect 252520 124080 252526 124092
rect 263042 124080 263048 124092
rect 252520 124052 263048 124080
rect 252520 124040 252526 124052
rect 263042 124040 263048 124052
rect 263100 124040 263106 124092
rect 251174 123496 251180 123548
rect 251232 123536 251238 123548
rect 253290 123536 253296 123548
rect 251232 123508 253296 123536
rect 251232 123496 251238 123508
rect 253290 123496 253296 123508
rect 253348 123496 253354 123548
rect 338206 123428 338212 123480
rect 338264 123468 338270 123480
rect 397362 123468 397368 123480
rect 338264 123440 397368 123468
rect 338264 123428 338270 123440
rect 397362 123428 397368 123440
rect 397420 123428 397426 123480
rect 395430 123224 395436 123276
rect 395488 123264 395494 123276
rect 397454 123264 397460 123276
rect 395488 123236 397460 123264
rect 395488 123224 395494 123236
rect 397454 123224 397460 123236
rect 397512 123224 397518 123276
rect 300118 122952 300124 123004
rect 300176 122992 300182 123004
rect 307110 122992 307116 123004
rect 300176 122964 307116 122992
rect 300176 122952 300182 122964
rect 307110 122952 307116 122964
rect 307168 122952 307174 123004
rect 183002 122884 183008 122936
rect 183060 122924 183066 122936
rect 214006 122924 214012 122936
rect 183060 122896 214012 122924
rect 183060 122884 183066 122896
rect 214006 122884 214012 122896
rect 214064 122884 214070 122936
rect 289170 122884 289176 122936
rect 289228 122924 289234 122936
rect 306558 122924 306564 122936
rect 289228 122896 306564 122924
rect 289228 122884 289234 122896
rect 306558 122884 306564 122896
rect 306616 122884 306622 122936
rect 166350 122816 166356 122868
rect 166408 122856 166414 122868
rect 213914 122856 213920 122868
rect 166408 122828 213920 122856
rect 166408 122816 166414 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 260098 122816 260104 122868
rect 260156 122856 260162 122868
rect 307662 122856 307668 122868
rect 260156 122828 307668 122856
rect 260156 122816 260162 122828
rect 307662 122816 307668 122828
rect 307720 122816 307726 122868
rect 252462 122748 252468 122800
rect 252520 122788 252526 122800
rect 287882 122788 287888 122800
rect 252520 122760 287888 122788
rect 252520 122748 252526 122760
rect 287882 122748 287888 122760
rect 287940 122748 287946 122800
rect 324314 122748 324320 122800
rect 324372 122788 324378 122800
rect 345014 122788 345020 122800
rect 324372 122760 345020 122788
rect 324372 122748 324378 122760
rect 345014 122748 345020 122760
rect 345072 122748 345078 122800
rect 252002 122680 252008 122732
rect 252060 122720 252066 122732
rect 264606 122720 264612 122732
rect 252060 122692 264612 122720
rect 252060 122680 252066 122692
rect 264606 122680 264612 122692
rect 264664 122680 264670 122732
rect 452562 122612 452568 122664
rect 452620 122652 452626 122664
rect 459554 122652 459560 122664
rect 452620 122624 459560 122652
rect 452620 122612 452626 122624
rect 459554 122612 459560 122624
rect 459612 122612 459618 122664
rect 251358 122476 251364 122528
rect 251416 122516 251422 122528
rect 254578 122516 254584 122528
rect 251416 122488 254584 122516
rect 251416 122476 251422 122488
rect 254578 122476 254584 122488
rect 254636 122476 254642 122528
rect 395338 122272 395344 122324
rect 395396 122312 395402 122324
rect 397454 122312 397460 122324
rect 395396 122284 397460 122312
rect 395396 122272 395402 122284
rect 397454 122272 397460 122284
rect 397512 122272 397518 122324
rect 287790 121592 287796 121644
rect 287848 121632 287854 121644
rect 307662 121632 307668 121644
rect 287848 121604 307668 121632
rect 287848 121592 287854 121604
rect 307662 121592 307668 121604
rect 307720 121592 307726 121644
rect 189902 121524 189908 121576
rect 189960 121564 189966 121576
rect 213914 121564 213920 121576
rect 189960 121536 213920 121564
rect 189960 121524 189966 121536
rect 213914 121524 213920 121536
rect 213972 121524 213978 121576
rect 283558 121524 283564 121576
rect 283616 121564 283622 121576
rect 307478 121564 307484 121576
rect 283616 121536 307484 121564
rect 283616 121524 283622 121536
rect 307478 121524 307484 121536
rect 307536 121524 307542 121576
rect 169018 121456 169024 121508
rect 169076 121496 169082 121508
rect 214006 121496 214012 121508
rect 169076 121468 214012 121496
rect 169076 121456 169082 121468
rect 214006 121456 214012 121468
rect 214064 121456 214070 121508
rect 264330 121456 264336 121508
rect 264388 121496 264394 121508
rect 307570 121496 307576 121508
rect 264388 121468 307576 121496
rect 264388 121456 264394 121468
rect 307570 121456 307576 121468
rect 307628 121456 307634 121508
rect 252462 121388 252468 121440
rect 252520 121428 252526 121440
rect 280890 121428 280896 121440
rect 252520 121400 280896 121428
rect 252520 121388 252526 121400
rect 280890 121388 280896 121400
rect 280948 121388 280954 121440
rect 324314 121388 324320 121440
rect 324372 121428 324378 121440
rect 324372 121400 345014 121428
rect 324372 121388 324378 121400
rect 251818 121320 251824 121372
rect 251876 121360 251882 121372
rect 261570 121360 261576 121372
rect 251876 121332 261576 121360
rect 251876 121320 251882 121332
rect 261570 121320 261576 121332
rect 261628 121320 261634 121372
rect 324406 121320 324412 121372
rect 324464 121360 324470 121372
rect 338114 121360 338120 121372
rect 324464 121332 338120 121360
rect 324464 121320 324470 121332
rect 338114 121320 338120 121332
rect 338172 121320 338178 121372
rect 344986 121360 345014 121400
rect 367002 121388 367008 121440
rect 367060 121428 367066 121440
rect 397454 121428 397460 121440
rect 367060 121400 397460 121428
rect 367060 121388 367066 121400
rect 397454 121388 397460 121400
rect 397512 121388 397518 121440
rect 346578 121360 346584 121372
rect 344986 121332 346584 121360
rect 346578 121320 346584 121332
rect 346636 121360 346642 121372
rect 370498 121360 370504 121372
rect 346636 121332 370504 121360
rect 346636 121320 346642 121332
rect 370498 121320 370504 121332
rect 370556 121320 370562 121372
rect 252370 120232 252376 120284
rect 252428 120272 252434 120284
rect 258994 120272 259000 120284
rect 252428 120244 259000 120272
rect 252428 120232 252434 120244
rect 258994 120232 259000 120244
rect 259052 120232 259058 120284
rect 301498 120232 301504 120284
rect 301556 120272 301562 120284
rect 306742 120272 306748 120284
rect 301556 120244 306748 120272
rect 301556 120232 301562 120244
rect 306742 120232 306748 120244
rect 306800 120232 306806 120284
rect 206462 120164 206468 120216
rect 206520 120204 206526 120216
rect 214006 120204 214012 120216
rect 206520 120176 214012 120204
rect 206520 120164 206526 120176
rect 214006 120164 214012 120176
rect 214064 120164 214070 120216
rect 279510 120164 279516 120216
rect 279568 120204 279574 120216
rect 307570 120204 307576 120216
rect 279568 120176 307576 120204
rect 279568 120164 279574 120176
rect 307570 120164 307576 120176
rect 307628 120164 307634 120216
rect 169294 120096 169300 120148
rect 169352 120136 169358 120148
rect 213914 120136 213920 120148
rect 169352 120108 213920 120136
rect 169352 120096 169358 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 261478 120096 261484 120148
rect 261536 120136 261542 120148
rect 307662 120136 307668 120148
rect 261536 120108 307668 120136
rect 261536 120096 261542 120108
rect 307662 120096 307668 120108
rect 307720 120096 307726 120148
rect 252462 120028 252468 120080
rect 252520 120068 252526 120080
rect 292206 120068 292212 120080
rect 252520 120040 292212 120068
rect 252520 120028 252526 120040
rect 292206 120028 292212 120040
rect 292264 120028 292270 120080
rect 324314 120028 324320 120080
rect 324372 120068 324378 120080
rect 346486 120068 346492 120080
rect 324372 120040 346492 120068
rect 324372 120028 324378 120040
rect 346486 120028 346492 120040
rect 346544 120028 346550 120080
rect 383010 120028 383016 120080
rect 383068 120068 383074 120080
rect 397454 120068 397460 120080
rect 383068 120040 397460 120068
rect 383068 120028 383074 120040
rect 397454 120028 397460 120040
rect 397512 120028 397518 120080
rect 251358 119960 251364 120012
rect 251416 120000 251422 120012
rect 272518 120000 272524 120012
rect 251416 119972 272524 120000
rect 251416 119960 251422 119972
rect 272518 119960 272524 119972
rect 272576 119960 272582 120012
rect 271414 119348 271420 119400
rect 271472 119388 271478 119400
rect 307294 119388 307300 119400
rect 271472 119360 307300 119388
rect 271472 119348 271478 119360
rect 307294 119348 307300 119360
rect 307352 119348 307358 119400
rect 325050 119348 325056 119400
rect 325108 119388 325114 119400
rect 333974 119388 333980 119400
rect 325108 119360 333980 119388
rect 325108 119348 325114 119360
rect 333974 119348 333980 119360
rect 334032 119348 334038 119400
rect 252278 119280 252284 119332
rect 252336 119320 252342 119332
rect 260282 119320 260288 119332
rect 252336 119292 260288 119320
rect 252336 119280 252342 119292
rect 260282 119280 260288 119292
rect 260340 119280 260346 119332
rect 211890 118804 211896 118856
rect 211948 118844 211954 118856
rect 214098 118844 214104 118856
rect 211948 118816 214104 118844
rect 211948 118804 211954 118816
rect 214098 118804 214104 118816
rect 214156 118804 214162 118856
rect 302970 118804 302976 118856
rect 303028 118844 303034 118856
rect 307662 118844 307668 118856
rect 303028 118816 307668 118844
rect 303028 118804 303034 118816
rect 307662 118804 307668 118816
rect 307720 118804 307726 118856
rect 173342 118736 173348 118788
rect 173400 118776 173406 118788
rect 213914 118776 213920 118788
rect 173400 118748 213920 118776
rect 173400 118736 173406 118748
rect 213914 118736 213920 118748
rect 213972 118736 213978 118788
rect 292114 118736 292120 118788
rect 292172 118776 292178 118788
rect 307570 118776 307576 118788
rect 292172 118748 307576 118776
rect 292172 118736 292178 118748
rect 307570 118736 307576 118748
rect 307628 118736 307634 118788
rect 167730 118668 167736 118720
rect 167788 118708 167794 118720
rect 214006 118708 214012 118720
rect 167788 118680 214012 118708
rect 167788 118668 167794 118680
rect 214006 118668 214012 118680
rect 214064 118668 214070 118720
rect 282362 118668 282368 118720
rect 282420 118708 282426 118720
rect 307478 118708 307484 118720
rect 282420 118680 307484 118708
rect 282420 118668 282426 118680
rect 307478 118668 307484 118680
rect 307536 118668 307542 118720
rect 251818 118600 251824 118652
rect 251876 118640 251882 118652
rect 293402 118640 293408 118652
rect 251876 118612 293408 118640
rect 251876 118600 251882 118612
rect 293402 118600 293408 118612
rect 293460 118600 293466 118652
rect 324314 118600 324320 118652
rect 324372 118640 324378 118652
rect 354766 118640 354772 118652
rect 324372 118612 354772 118640
rect 324372 118600 324378 118612
rect 354766 118600 354772 118612
rect 354824 118600 354830 118652
rect 452470 118600 452476 118652
rect 452528 118640 452534 118652
rect 484394 118640 484400 118652
rect 452528 118612 484400 118640
rect 452528 118600 452534 118612
rect 484394 118600 484400 118612
rect 484452 118600 484458 118652
rect 252462 118532 252468 118584
rect 252520 118572 252526 118584
rect 262858 118572 262864 118584
rect 252520 118544 262864 118572
rect 252520 118532 252526 118544
rect 262858 118532 262864 118544
rect 262916 118532 262922 118584
rect 254578 117512 254584 117564
rect 254636 117552 254642 117564
rect 307662 117552 307668 117564
rect 254636 117524 307668 117552
rect 254636 117512 254642 117524
rect 307662 117512 307668 117524
rect 307720 117512 307726 117564
rect 298830 117444 298836 117496
rect 298888 117484 298894 117496
rect 306558 117484 306564 117496
rect 298888 117456 306564 117484
rect 298888 117444 298894 117456
rect 306558 117444 306564 117456
rect 306616 117444 306622 117496
rect 188430 117376 188436 117428
rect 188488 117416 188494 117428
rect 214006 117416 214012 117428
rect 188488 117388 214012 117416
rect 188488 117376 188494 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 293218 117376 293224 117428
rect 293276 117416 293282 117428
rect 307662 117416 307668 117428
rect 293276 117388 307668 117416
rect 293276 117376 293282 117388
rect 307662 117376 307668 117388
rect 307720 117376 307726 117428
rect 169202 117308 169208 117360
rect 169260 117348 169266 117360
rect 213914 117348 213920 117360
rect 169260 117320 213920 117348
rect 169260 117308 169266 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 304442 117308 304448 117360
rect 304500 117348 304506 117360
rect 307570 117348 307576 117360
rect 304500 117320 307576 117348
rect 304500 117308 304506 117320
rect 307570 117308 307576 117320
rect 307628 117308 307634 117360
rect 251358 117240 251364 117292
rect 251416 117280 251422 117292
rect 261662 117280 261668 117292
rect 251416 117252 261668 117280
rect 251416 117240 251422 117252
rect 261662 117240 261668 117252
rect 261720 117240 261726 117292
rect 347222 117240 347228 117292
rect 347280 117280 347286 117292
rect 365070 117280 365076 117292
rect 347280 117252 365076 117280
rect 347280 117240 347286 117252
rect 365070 117240 365076 117252
rect 365128 117240 365134 117292
rect 380158 117240 380164 117292
rect 380216 117280 380222 117292
rect 397454 117280 397460 117292
rect 380216 117252 397460 117280
rect 380216 117240 380222 117252
rect 397454 117240 397460 117252
rect 397512 117240 397518 117292
rect 449342 117240 449348 117292
rect 449400 117280 449406 117292
rect 503714 117280 503720 117292
rect 449400 117252 503720 117280
rect 449400 117240 449406 117252
rect 503714 117240 503720 117252
rect 503772 117240 503778 117292
rect 252462 117172 252468 117224
rect 252520 117212 252526 117224
rect 258810 117212 258816 117224
rect 252520 117184 258816 117212
rect 252520 117172 252526 117184
rect 258810 117172 258816 117184
rect 258868 117172 258874 117224
rect 252002 116560 252008 116612
rect 252060 116600 252066 116612
rect 305730 116600 305736 116612
rect 252060 116572 305736 116600
rect 252060 116560 252066 116572
rect 305730 116560 305736 116572
rect 305788 116560 305794 116612
rect 324314 116560 324320 116612
rect 324372 116600 324378 116612
rect 347222 116600 347228 116612
rect 324372 116572 347228 116600
rect 324372 116560 324378 116572
rect 347222 116560 347228 116572
rect 347280 116560 347286 116612
rect 185670 116016 185676 116068
rect 185728 116056 185734 116068
rect 213914 116056 213920 116068
rect 185728 116028 213920 116056
rect 185728 116016 185734 116028
rect 213914 116016 213920 116028
rect 213972 116016 213978 116068
rect 272518 116016 272524 116068
rect 272576 116056 272582 116068
rect 306742 116056 306748 116068
rect 272576 116028 306748 116056
rect 272576 116016 272582 116028
rect 306742 116016 306748 116028
rect 306800 116016 306806 116068
rect 181530 115948 181536 116000
rect 181588 115988 181594 116000
rect 214006 115988 214012 116000
rect 181588 115960 214012 115988
rect 181588 115948 181594 115960
rect 214006 115948 214012 115960
rect 214064 115948 214070 116000
rect 262858 115948 262864 116000
rect 262916 115988 262922 116000
rect 307478 115988 307484 116000
rect 262916 115960 307484 115988
rect 262916 115948 262922 115960
rect 307478 115948 307484 115960
rect 307536 115948 307542 116000
rect 252278 115880 252284 115932
rect 252336 115920 252342 115932
rect 285122 115920 285128 115932
rect 252336 115892 285128 115920
rect 252336 115880 252342 115892
rect 285122 115880 285128 115892
rect 285180 115880 285186 115932
rect 324314 115880 324320 115932
rect 324372 115920 324378 115932
rect 342346 115920 342352 115932
rect 324372 115892 342352 115920
rect 324372 115880 324378 115892
rect 342346 115880 342352 115892
rect 342404 115880 342410 115932
rect 354582 115880 354588 115932
rect 354640 115920 354646 115932
rect 397454 115920 397460 115932
rect 354640 115892 397460 115920
rect 354640 115880 354646 115892
rect 397454 115880 397460 115892
rect 397512 115880 397518 115932
rect 251910 115812 251916 115864
rect 251968 115852 251974 115864
rect 262950 115852 262956 115864
rect 251968 115824 262956 115852
rect 251968 115812 251974 115824
rect 262950 115812 262956 115824
rect 263008 115812 263014 115864
rect 451550 115812 451556 115864
rect 451608 115852 451614 115864
rect 455506 115852 455512 115864
rect 451608 115824 455512 115852
rect 451608 115812 451614 115824
rect 455506 115812 455512 115824
rect 455564 115812 455570 115864
rect 324958 115268 324964 115320
rect 325016 115308 325022 115320
rect 332594 115308 332600 115320
rect 325016 115280 332600 115308
rect 325016 115268 325022 115280
rect 332594 115268 332600 115280
rect 332652 115268 332658 115320
rect 251818 115200 251824 115252
rect 251876 115240 251882 115252
rect 268562 115240 268568 115252
rect 251876 115212 268568 115240
rect 251876 115200 251882 115212
rect 268562 115200 268568 115212
rect 268620 115200 268626 115252
rect 286410 115200 286416 115252
rect 286468 115240 286474 115252
rect 307386 115240 307392 115252
rect 286468 115212 307392 115240
rect 286468 115200 286474 115212
rect 307386 115200 307392 115212
rect 307444 115200 307450 115252
rect 323578 115200 323584 115252
rect 323636 115240 323642 115252
rect 337378 115240 337384 115252
rect 323636 115212 337384 115240
rect 323636 115200 323642 115212
rect 337378 115200 337384 115212
rect 337436 115200 337442 115252
rect 203702 114588 203708 114640
rect 203760 114628 203766 114640
rect 214006 114628 214012 114640
rect 203760 114600 214012 114628
rect 203760 114588 203766 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 294598 114588 294604 114640
rect 294656 114628 294662 114640
rect 307570 114628 307576 114640
rect 294656 114600 307576 114628
rect 294656 114588 294662 114600
rect 307570 114588 307576 114600
rect 307628 114588 307634 114640
rect 184290 114520 184296 114572
rect 184348 114560 184354 114572
rect 213914 114560 213920 114572
rect 184348 114532 213920 114560
rect 184348 114520 184354 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 265618 114520 265624 114572
rect 265676 114560 265682 114572
rect 307662 114560 307668 114572
rect 265676 114532 307668 114560
rect 265676 114520 265682 114532
rect 307662 114520 307668 114532
rect 307720 114520 307726 114572
rect 251358 114452 251364 114504
rect 251416 114492 251422 114504
rect 265710 114492 265716 114504
rect 251416 114464 265716 114492
rect 251416 114452 251422 114464
rect 265710 114452 265716 114464
rect 265768 114452 265774 114504
rect 324314 114452 324320 114504
rect 324372 114492 324378 114504
rect 358814 114492 358820 114504
rect 324372 114464 358820 114492
rect 324372 114452 324378 114464
rect 358814 114452 358820 114464
rect 358872 114452 358878 114504
rect 362862 114452 362868 114504
rect 362920 114492 362926 114504
rect 397454 114492 397460 114504
rect 362920 114464 397460 114492
rect 362920 114452 362926 114464
rect 397454 114452 397460 114464
rect 397512 114452 397518 114504
rect 452470 114452 452476 114504
rect 452528 114492 452534 114504
rect 485774 114492 485780 114504
rect 452528 114464 485780 114492
rect 452528 114452 452534 114464
rect 485774 114452 485780 114464
rect 485832 114452 485838 114504
rect 324406 114384 324412 114436
rect 324464 114424 324470 114436
rect 351914 114424 351920 114436
rect 324464 114396 351920 114424
rect 324464 114384 324470 114396
rect 351914 114384 351920 114396
rect 351972 114424 351978 114436
rect 363598 114424 363604 114436
rect 351972 114396 363604 114424
rect 351972 114384 351978 114396
rect 363598 114384 363604 114396
rect 363656 114384 363662 114436
rect 251634 114180 251640 114232
rect 251692 114220 251698 114232
rect 254762 114220 254768 114232
rect 251692 114192 254768 114220
rect 251692 114180 251698 114192
rect 254762 114180 254768 114192
rect 254820 114180 254826 114232
rect 252462 113772 252468 113824
rect 252520 113812 252526 113824
rect 271138 113812 271144 113824
rect 252520 113784 271144 113812
rect 252520 113772 252526 113784
rect 271138 113772 271144 113784
rect 271196 113772 271202 113824
rect 360194 113772 360200 113824
rect 360252 113812 360258 113824
rect 387150 113812 387156 113824
rect 360252 113784 387156 113812
rect 360252 113772 360258 113784
rect 387150 113772 387156 113784
rect 387208 113772 387214 113824
rect 295978 113296 295984 113348
rect 296036 113336 296042 113348
rect 306558 113336 306564 113348
rect 296036 113308 306564 113336
rect 296036 113296 296042 113308
rect 306558 113296 306564 113308
rect 306616 113296 306622 113348
rect 198090 113228 198096 113280
rect 198148 113268 198154 113280
rect 214006 113268 214012 113280
rect 198148 113240 214012 113268
rect 198148 113228 198154 113240
rect 214006 113228 214012 113240
rect 214064 113228 214070 113280
rect 279418 113228 279424 113280
rect 279476 113268 279482 113280
rect 306926 113268 306932 113280
rect 279476 113240 306932 113268
rect 279476 113228 279482 113240
rect 306926 113228 306932 113240
rect 306984 113228 306990 113280
rect 173250 113160 173256 113212
rect 173308 113200 173314 113212
rect 213914 113200 213920 113212
rect 173308 113172 213920 113200
rect 173308 113160 173314 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 268378 113160 268384 113212
rect 268436 113200 268442 113212
rect 307662 113200 307668 113212
rect 268436 113172 307668 113200
rect 268436 113160 268442 113172
rect 307662 113160 307668 113172
rect 307720 113160 307726 113212
rect 395982 113092 395988 113144
rect 396040 113132 396046 113144
rect 397454 113132 397460 113144
rect 396040 113104 397460 113132
rect 396040 113092 396046 113104
rect 397454 113092 397460 113104
rect 397512 113092 397518 113144
rect 456058 113092 456064 113144
rect 456116 113132 456122 113144
rect 580166 113132 580172 113144
rect 456116 113104 580172 113132
rect 456116 113092 456122 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 252462 112820 252468 112872
rect 252520 112860 252526 112872
rect 257430 112860 257436 112872
rect 252520 112832 257436 112860
rect 252520 112820 252526 112832
rect 257430 112820 257436 112832
rect 257488 112820 257494 112872
rect 252186 112480 252192 112532
rect 252244 112520 252250 112532
rect 271322 112520 271328 112532
rect 252244 112492 271328 112520
rect 252244 112480 252250 112492
rect 271322 112480 271328 112492
rect 271380 112480 271386 112532
rect 257522 112412 257528 112464
rect 257580 112452 257586 112464
rect 307202 112452 307208 112464
rect 257580 112424 307208 112452
rect 257580 112412 257586 112424
rect 307202 112412 307208 112424
rect 307260 112412 307266 112464
rect 251634 112208 251640 112260
rect 251692 112248 251698 112260
rect 254854 112248 254860 112260
rect 251692 112220 254860 112248
rect 251692 112208 251698 112220
rect 254854 112208 254860 112220
rect 254912 112208 254918 112260
rect 202322 111868 202328 111920
rect 202380 111908 202386 111920
rect 214006 111908 214012 111920
rect 202380 111880 214012 111908
rect 202380 111868 202386 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 301590 111868 301596 111920
rect 301648 111908 301654 111920
rect 307662 111908 307668 111920
rect 301648 111880 307668 111908
rect 301648 111868 301654 111880
rect 307662 111868 307668 111880
rect 307720 111868 307726 111920
rect 169110 111800 169116 111852
rect 169168 111840 169174 111852
rect 213914 111840 213920 111852
rect 169168 111812 213920 111840
rect 169168 111800 169174 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 271230 111800 271236 111852
rect 271288 111840 271294 111852
rect 307478 111840 307484 111852
rect 271288 111812 307484 111840
rect 271288 111800 271294 111812
rect 307478 111800 307484 111812
rect 307536 111800 307542 111852
rect 168282 111732 168288 111784
rect 168340 111772 168346 111784
rect 196710 111772 196716 111784
rect 168340 111744 196716 111772
rect 168340 111732 168346 111744
rect 196710 111732 196716 111744
rect 196768 111732 196774 111784
rect 387058 111732 387064 111784
rect 387116 111772 387122 111784
rect 397454 111772 397460 111784
rect 387116 111744 397460 111772
rect 387116 111732 387122 111744
rect 397454 111732 397460 111744
rect 397512 111732 397518 111784
rect 452470 111732 452476 111784
rect 452528 111772 452534 111784
rect 469214 111772 469220 111784
rect 452528 111744 469220 111772
rect 452528 111732 452534 111744
rect 469214 111732 469220 111744
rect 469272 111732 469278 111784
rect 390462 111664 390468 111716
rect 390520 111704 390526 111716
rect 399570 111704 399576 111716
rect 390520 111676 399576 111704
rect 390520 111664 390526 111676
rect 399570 111664 399576 111676
rect 399628 111664 399634 111716
rect 452562 111664 452568 111716
rect 452620 111704 452626 111716
rect 466454 111704 466460 111716
rect 452620 111676 466460 111704
rect 452620 111664 452626 111676
rect 466454 111664 466460 111676
rect 466512 111664 466518 111716
rect 251818 111256 251824 111308
rect 251876 111296 251882 111308
rect 260374 111296 260380 111308
rect 251876 111268 260380 111296
rect 251876 111256 251882 111268
rect 260374 111256 260380 111268
rect 260432 111256 260438 111308
rect 252278 111052 252284 111104
rect 252336 111092 252342 111104
rect 305638 111092 305644 111104
rect 252336 111064 305644 111092
rect 252336 111052 252342 111064
rect 305638 111052 305644 111064
rect 305696 111052 305702 111104
rect 345658 111052 345664 111104
rect 345716 111092 345722 111104
rect 397546 111092 397552 111104
rect 345716 111064 397552 111092
rect 345716 111052 345722 111064
rect 397546 111052 397552 111064
rect 397604 111052 397610 111104
rect 304258 110576 304264 110628
rect 304316 110616 304322 110628
rect 307478 110616 307484 110628
rect 304316 110588 307484 110616
rect 304316 110576 304322 110588
rect 307478 110576 307484 110588
rect 307536 110576 307542 110628
rect 263042 110508 263048 110560
rect 263100 110548 263106 110560
rect 307570 110548 307576 110560
rect 263100 110520 307576 110548
rect 263100 110508 263106 110520
rect 307570 110508 307576 110520
rect 307628 110508 307634 110560
rect 173434 110440 173440 110492
rect 173492 110480 173498 110492
rect 213914 110480 213920 110492
rect 173492 110452 213920 110480
rect 173492 110440 173498 110452
rect 213914 110440 213920 110452
rect 213972 110440 213978 110492
rect 253290 110440 253296 110492
rect 253348 110480 253354 110492
rect 307662 110480 307668 110492
rect 253348 110452 307668 110480
rect 253348 110440 253354 110452
rect 307662 110440 307668 110452
rect 307720 110440 307726 110492
rect 167822 110372 167828 110424
rect 167880 110412 167886 110424
rect 194042 110412 194048 110424
rect 167880 110384 194048 110412
rect 167880 110372 167886 110384
rect 194042 110372 194048 110384
rect 194100 110372 194106 110424
rect 251910 110372 251916 110424
rect 251968 110412 251974 110424
rect 289354 110412 289360 110424
rect 251968 110384 289360 110412
rect 251968 110372 251974 110384
rect 289354 110372 289360 110384
rect 289412 110372 289418 110424
rect 324314 110372 324320 110424
rect 324372 110412 324378 110424
rect 347774 110412 347780 110424
rect 324372 110384 347780 110412
rect 324372 110372 324378 110384
rect 347774 110372 347780 110384
rect 347832 110372 347838 110424
rect 378778 110372 378784 110424
rect 378836 110412 378842 110424
rect 397454 110412 397460 110424
rect 378836 110384 397460 110412
rect 378836 110372 378842 110384
rect 397454 110372 397460 110384
rect 397512 110372 397518 110424
rect 252462 110304 252468 110356
rect 252520 110344 252526 110356
rect 273898 110344 273904 110356
rect 252520 110316 273904 110344
rect 252520 110304 252526 110316
rect 273898 110304 273904 110316
rect 273956 110304 273962 110356
rect 452102 110304 452108 110356
rect 452160 110344 452166 110356
rect 456886 110344 456892 110356
rect 452160 110316 456892 110344
rect 452160 110304 452166 110316
rect 456886 110304 456892 110316
rect 456944 110304 456950 110356
rect 252094 110236 252100 110288
rect 252152 110276 252158 110288
rect 256142 110276 256148 110288
rect 252152 110248 256148 110276
rect 252152 110236 252158 110248
rect 256142 110236 256148 110248
rect 256200 110236 256206 110288
rect 300394 109148 300400 109200
rect 300452 109188 300458 109200
rect 307478 109188 307484 109200
rect 300452 109160 307484 109188
rect 300452 109148 300458 109160
rect 307478 109148 307484 109160
rect 307536 109148 307542 109200
rect 174722 109080 174728 109132
rect 174780 109120 174786 109132
rect 214006 109120 214012 109132
rect 174780 109092 214012 109120
rect 174780 109080 174786 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 275370 109080 275376 109132
rect 275428 109120 275434 109132
rect 307570 109120 307576 109132
rect 275428 109092 307576 109120
rect 275428 109080 275434 109092
rect 307570 109080 307576 109092
rect 307628 109080 307634 109132
rect 170582 109012 170588 109064
rect 170640 109052 170646 109064
rect 213914 109052 213920 109064
rect 170640 109024 213920 109052
rect 170640 109012 170646 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 258810 109012 258816 109064
rect 258868 109052 258874 109064
rect 307662 109052 307668 109064
rect 258868 109024 307668 109052
rect 258868 109012 258874 109024
rect 307662 109012 307668 109024
rect 307720 109012 307726 109064
rect 395338 109012 395344 109064
rect 395396 109052 395402 109064
rect 397730 109052 397736 109064
rect 395396 109024 397736 109052
rect 395396 109012 395402 109024
rect 397730 109012 397736 109024
rect 397788 109012 397794 109064
rect 168098 108944 168104 108996
rect 168156 108984 168162 108996
rect 189810 108984 189816 108996
rect 168156 108956 189816 108984
rect 168156 108944 168162 108956
rect 189810 108944 189816 108956
rect 189868 108944 189874 108996
rect 252370 108944 252376 108996
rect 252428 108984 252434 108996
rect 296254 108984 296260 108996
rect 252428 108956 296260 108984
rect 252428 108944 252434 108956
rect 296254 108944 296260 108956
rect 296312 108944 296318 108996
rect 324406 108944 324412 108996
rect 324464 108984 324470 108996
rect 366358 108984 366364 108996
rect 324464 108956 366364 108984
rect 324464 108944 324470 108956
rect 366358 108944 366364 108956
rect 366416 108944 366422 108996
rect 252462 108876 252468 108928
rect 252520 108916 252526 108928
rect 272610 108916 272616 108928
rect 252520 108888 272616 108916
rect 252520 108876 252526 108888
rect 272610 108876 272616 108888
rect 272668 108876 272674 108928
rect 324314 108876 324320 108928
rect 324372 108916 324378 108928
rect 340138 108916 340144 108928
rect 324372 108888 340144 108916
rect 324372 108876 324378 108888
rect 340138 108876 340144 108888
rect 340196 108876 340202 108928
rect 249150 107856 249156 107908
rect 249208 107896 249214 107908
rect 307662 107896 307668 107908
rect 249208 107868 307668 107896
rect 249208 107856 249214 107868
rect 307662 107856 307668 107868
rect 307720 107856 307726 107908
rect 296162 107788 296168 107840
rect 296220 107828 296226 107840
rect 307570 107828 307576 107840
rect 296220 107800 307576 107828
rect 296220 107788 296226 107800
rect 307570 107788 307576 107800
rect 307628 107788 307634 107840
rect 170674 107720 170680 107772
rect 170732 107760 170738 107772
rect 214006 107760 214012 107772
rect 170732 107732 214012 107760
rect 170732 107720 170738 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 273898 107720 273904 107772
rect 273956 107760 273962 107772
rect 307662 107760 307668 107772
rect 273956 107732 307668 107760
rect 273956 107720 273962 107732
rect 307662 107720 307668 107732
rect 307720 107720 307726 107772
rect 166442 107652 166448 107704
rect 166500 107692 166506 107704
rect 213914 107692 213920 107704
rect 166500 107664 213920 107692
rect 166500 107652 166506 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 363598 107652 363604 107704
rect 363656 107692 363662 107704
rect 397454 107692 397460 107704
rect 363656 107664 397460 107692
rect 363656 107652 363662 107664
rect 397454 107652 397460 107664
rect 397512 107652 397518 107704
rect 252094 107584 252100 107636
rect 252152 107624 252158 107636
rect 274174 107624 274180 107636
rect 252152 107596 274180 107624
rect 252152 107584 252158 107596
rect 274174 107584 274180 107596
rect 274232 107584 274238 107636
rect 323302 107584 323308 107636
rect 323360 107624 323366 107636
rect 367738 107624 367744 107636
rect 323360 107596 367744 107624
rect 323360 107584 323366 107596
rect 367738 107584 367744 107596
rect 367796 107584 367802 107636
rect 252002 106904 252008 106956
rect 252060 106944 252066 106956
rect 308398 106944 308404 106956
rect 252060 106916 308404 106944
rect 252060 106904 252066 106916
rect 308398 106904 308404 106916
rect 308456 106904 308462 106956
rect 376018 106904 376024 106956
rect 376076 106944 376082 106956
rect 397638 106944 397644 106956
rect 376076 106916 397644 106944
rect 376076 106904 376082 106916
rect 397638 106904 397644 106916
rect 397696 106904 397702 106956
rect 274082 106428 274088 106480
rect 274140 106468 274146 106480
rect 307662 106468 307668 106480
rect 274140 106440 307668 106468
rect 274140 106428 274146 106440
rect 307662 106428 307668 106440
rect 307720 106428 307726 106480
rect 204990 106360 204996 106412
rect 205048 106400 205054 106412
rect 214006 106400 214012 106412
rect 205048 106372 214012 106400
rect 205048 106360 205054 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 285122 106360 285128 106412
rect 285180 106400 285186 106412
rect 307570 106400 307576 106412
rect 285180 106372 307576 106400
rect 285180 106360 285186 106372
rect 307570 106360 307576 106372
rect 307628 106360 307634 106412
rect 194042 106292 194048 106344
rect 194100 106332 194106 106344
rect 213914 106332 213920 106344
rect 194100 106304 213920 106332
rect 194100 106292 194106 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 252462 106224 252468 106276
rect 252520 106264 252526 106276
rect 304534 106264 304540 106276
rect 252520 106236 304540 106264
rect 252520 106224 252526 106236
rect 304534 106224 304540 106236
rect 304592 106224 304598 106276
rect 324314 106224 324320 106276
rect 324372 106264 324378 106276
rect 356146 106264 356152 106276
rect 324372 106236 356152 106264
rect 324372 106224 324378 106236
rect 356146 106224 356152 106236
rect 356204 106264 356210 106276
rect 363782 106264 363788 106276
rect 356204 106236 363788 106264
rect 356204 106224 356210 106236
rect 363782 106224 363788 106236
rect 363840 106224 363846 106276
rect 251910 106156 251916 106208
rect 251968 106196 251974 106208
rect 294690 106196 294696 106208
rect 251968 106168 294696 106196
rect 251968 106156 251974 106168
rect 294690 106156 294696 106168
rect 294748 106156 294754 106208
rect 251358 106088 251364 106140
rect 251416 106128 251422 106140
rect 254670 106128 254676 106140
rect 251416 106100 254676 106128
rect 251416 106088 251422 106100
rect 254670 106088 254676 106100
rect 254728 106088 254734 106140
rect 182818 105544 182824 105596
rect 182876 105584 182882 105596
rect 216030 105584 216036 105596
rect 182876 105556 216036 105584
rect 182876 105544 182882 105556
rect 216030 105544 216036 105556
rect 216088 105544 216094 105596
rect 365070 105544 365076 105596
rect 365128 105584 365134 105596
rect 397454 105584 397460 105596
rect 365128 105556 397460 105584
rect 365128 105544 365134 105556
rect 397454 105544 397460 105556
rect 397512 105544 397518 105596
rect 211982 105000 211988 105052
rect 212040 105040 212046 105052
rect 213914 105040 213920 105052
rect 212040 105012 213920 105040
rect 212040 105000 212046 105012
rect 213914 105000 213920 105012
rect 213972 105000 213978 105052
rect 294782 105000 294788 105052
rect 294840 105040 294846 105052
rect 307662 105040 307668 105052
rect 294840 105012 307668 105040
rect 294840 105000 294846 105012
rect 307662 105000 307668 105012
rect 307720 105000 307726 105052
rect 198182 104932 198188 104984
rect 198240 104972 198246 104984
rect 214006 104972 214012 104984
rect 198240 104944 214012 104972
rect 198240 104932 198246 104944
rect 214006 104932 214012 104944
rect 214064 104932 214070 104984
rect 196802 104864 196808 104916
rect 196860 104904 196866 104916
rect 213914 104904 213920 104916
rect 196860 104876 213920 104904
rect 196860 104864 196866 104876
rect 213914 104864 213920 104876
rect 213972 104864 213978 104916
rect 304626 104864 304632 104916
rect 304684 104904 304690 104916
rect 307570 104904 307576 104916
rect 304684 104876 307576 104904
rect 304684 104864 304690 104876
rect 307570 104864 307576 104876
rect 307628 104864 307634 104916
rect 452562 104864 452568 104916
rect 452620 104904 452626 104916
rect 454218 104904 454224 104916
rect 452620 104876 454224 104904
rect 452620 104864 452626 104876
rect 454218 104864 454224 104876
rect 454276 104864 454282 104916
rect 251910 104796 251916 104848
rect 251968 104836 251974 104848
rect 308490 104836 308496 104848
rect 251968 104808 308496 104836
rect 251968 104796 251974 104808
rect 308490 104796 308496 104808
rect 308548 104796 308554 104848
rect 324314 104796 324320 104848
rect 324372 104836 324378 104848
rect 335538 104836 335544 104848
rect 324372 104808 335544 104836
rect 324372 104796 324378 104808
rect 335538 104796 335544 104808
rect 335596 104796 335602 104848
rect 378962 104796 378968 104848
rect 379020 104836 379026 104848
rect 397546 104836 397552 104848
rect 379020 104808 397552 104836
rect 379020 104796 379026 104808
rect 397546 104796 397552 104808
rect 397604 104796 397610 104848
rect 252462 104728 252468 104780
rect 252520 104768 252526 104780
rect 287974 104768 287980 104780
rect 252520 104740 287980 104768
rect 252520 104728 252526 104740
rect 287974 104728 287980 104740
rect 288032 104728 288038 104780
rect 252278 104116 252284 104168
rect 252336 104156 252342 104168
rect 293494 104156 293500 104168
rect 252336 104128 293500 104156
rect 252336 104116 252342 104128
rect 293494 104116 293500 104128
rect 293552 104116 293558 104168
rect 324498 104116 324504 104168
rect 324556 104156 324562 104168
rect 329098 104156 329104 104168
rect 324556 104128 329104 104156
rect 324556 104116 324562 104128
rect 329098 104116 329104 104128
rect 329156 104116 329162 104168
rect 293402 103640 293408 103692
rect 293460 103680 293466 103692
rect 307662 103680 307668 103692
rect 293460 103652 307668 103680
rect 293460 103640 293466 103652
rect 307662 103640 307668 103652
rect 307720 103640 307726 103692
rect 195330 103572 195336 103624
rect 195388 103612 195394 103624
rect 214006 103612 214012 103624
rect 195388 103584 214012 103612
rect 195388 103572 195394 103584
rect 214006 103572 214012 103584
rect 214064 103572 214070 103624
rect 287882 103572 287888 103624
rect 287940 103612 287946 103624
rect 307478 103612 307484 103624
rect 287940 103584 307484 103612
rect 287940 103572 287946 103584
rect 307478 103572 307484 103584
rect 307536 103572 307542 103624
rect 191190 103504 191196 103556
rect 191248 103544 191254 103556
rect 213914 103544 213920 103556
rect 191248 103516 213920 103544
rect 191248 103504 191254 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 262950 103504 262956 103556
rect 263008 103544 263014 103556
rect 307570 103544 307576 103556
rect 263008 103516 307576 103544
rect 263008 103504 263014 103516
rect 307570 103504 307576 103516
rect 307628 103504 307634 103556
rect 252462 103436 252468 103488
rect 252520 103476 252526 103488
rect 286410 103476 286416 103488
rect 252520 103448 286416 103476
rect 252520 103436 252526 103448
rect 286410 103436 286416 103448
rect 286468 103436 286474 103488
rect 321646 103436 321652 103488
rect 321704 103476 321710 103488
rect 374638 103476 374644 103488
rect 321704 103448 374644 103476
rect 321704 103436 321710 103448
rect 374638 103436 374644 103448
rect 374696 103436 374702 103488
rect 382090 103436 382096 103488
rect 382148 103476 382154 103488
rect 397546 103476 397552 103488
rect 382148 103448 397552 103476
rect 382148 103436 382154 103448
rect 397546 103436 397552 103448
rect 397604 103436 397610 103488
rect 252002 103368 252008 103420
rect 252060 103408 252066 103420
rect 264514 103408 264520 103420
rect 252060 103380 264520 103408
rect 252060 103368 252066 103380
rect 264514 103368 264520 103380
rect 264572 103368 264578 103420
rect 452562 103028 452568 103080
rect 452620 103068 452626 103080
rect 454126 103068 454132 103080
rect 452620 103040 454132 103068
rect 452620 103028 452626 103040
rect 454126 103028 454132 103040
rect 454184 103028 454190 103080
rect 252370 102960 252376 103012
rect 252428 103000 252434 103012
rect 257522 103000 257528 103012
rect 252428 102972 257528 103000
rect 252428 102960 252434 102972
rect 257522 102960 257528 102972
rect 257580 102960 257586 103012
rect 167914 102756 167920 102808
rect 167972 102796 167978 102808
rect 214650 102796 214656 102808
rect 167972 102768 214656 102796
rect 167972 102756 167978 102768
rect 214650 102756 214656 102768
rect 214708 102756 214714 102808
rect 303522 102348 303528 102400
rect 303580 102388 303586 102400
rect 308398 102388 308404 102400
rect 303580 102360 308404 102388
rect 303580 102348 303586 102360
rect 308398 102348 308404 102360
rect 308456 102348 308462 102400
rect 294690 102280 294696 102332
rect 294748 102320 294754 102332
rect 307662 102320 307668 102332
rect 294748 102292 307668 102320
rect 294748 102280 294754 102292
rect 307662 102280 307668 102292
rect 307720 102280 307726 102332
rect 209038 102212 209044 102264
rect 209096 102252 209102 102264
rect 214006 102252 214012 102264
rect 209096 102224 214012 102252
rect 209096 102212 209102 102224
rect 214006 102212 214012 102224
rect 214064 102212 214070 102264
rect 287974 102212 287980 102264
rect 288032 102252 288038 102264
rect 307478 102252 307484 102264
rect 288032 102224 307484 102252
rect 288032 102212 288038 102224
rect 307478 102212 307484 102224
rect 307536 102212 307542 102264
rect 189810 102144 189816 102196
rect 189868 102184 189874 102196
rect 213914 102184 213920 102196
rect 189868 102156 213920 102184
rect 189868 102144 189874 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 257430 102144 257436 102196
rect 257488 102184 257494 102196
rect 307570 102184 307576 102196
rect 257488 102156 307576 102184
rect 257488 102144 257494 102156
rect 307570 102144 307576 102156
rect 307628 102144 307634 102196
rect 252462 102076 252468 102128
rect 252520 102116 252526 102128
rect 271414 102116 271420 102128
rect 252520 102088 271420 102116
rect 252520 102076 252526 102088
rect 271414 102076 271420 102088
rect 271472 102076 271478 102128
rect 324314 102076 324320 102128
rect 324372 102116 324378 102128
rect 351362 102116 351368 102128
rect 324372 102088 351368 102116
rect 324372 102076 324378 102088
rect 351362 102076 351368 102088
rect 351420 102076 351426 102128
rect 388438 102076 388444 102128
rect 388496 102116 388502 102128
rect 397546 102116 397552 102128
rect 388496 102088 397552 102116
rect 388496 102076 388502 102088
rect 397546 102076 397552 102088
rect 397604 102076 397610 102128
rect 324406 102008 324412 102060
rect 324464 102048 324470 102060
rect 335354 102048 335360 102060
rect 324464 102020 335360 102048
rect 324464 102008 324470 102020
rect 335354 102008 335360 102020
rect 335412 102008 335418 102060
rect 393222 102008 393228 102060
rect 393280 102048 393286 102060
rect 397638 102048 397644 102060
rect 393280 102020 397644 102048
rect 393280 102008 393286 102020
rect 397638 102008 397644 102020
rect 397696 102008 397702 102060
rect 166534 101396 166540 101448
rect 166592 101436 166598 101448
rect 214558 101436 214564 101448
rect 166592 101408 214564 101436
rect 166592 101396 166598 101408
rect 214558 101396 214564 101408
rect 214616 101396 214622 101448
rect 252094 101396 252100 101448
rect 252152 101436 252158 101448
rect 297358 101436 297364 101448
rect 252152 101408 297364 101436
rect 252152 101396 252158 101408
rect 297358 101396 297364 101408
rect 297416 101396 297422 101448
rect 327074 101396 327080 101448
rect 327132 101436 327138 101448
rect 394050 101436 394056 101448
rect 327132 101408 394056 101436
rect 327132 101396 327138 101408
rect 394050 101396 394056 101408
rect 394108 101396 394114 101448
rect 257522 100920 257528 100972
rect 257580 100960 257586 100972
rect 307662 100960 307668 100972
rect 257580 100932 307668 100960
rect 257580 100920 257586 100932
rect 307662 100920 307668 100932
rect 307720 100920 307726 100972
rect 252002 100852 252008 100904
rect 252060 100892 252066 100904
rect 255958 100892 255964 100904
rect 252060 100864 255964 100892
rect 252060 100852 252066 100864
rect 255958 100852 255964 100864
rect 256016 100852 256022 100904
rect 296254 100784 296260 100836
rect 296312 100824 296318 100836
rect 307570 100824 307576 100836
rect 296312 100796 307576 100824
rect 296312 100784 296318 100796
rect 307570 100784 307576 100796
rect 307628 100784 307634 100836
rect 196710 100716 196716 100768
rect 196768 100756 196774 100768
rect 213914 100756 213920 100768
rect 196768 100728 213920 100756
rect 196768 100716 196774 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 301774 100716 301780 100768
rect 301832 100756 301838 100768
rect 306742 100756 306748 100768
rect 301832 100728 306748 100756
rect 301832 100716 301838 100728
rect 306742 100716 306748 100728
rect 306800 100716 306806 100768
rect 251726 100648 251732 100700
rect 251784 100688 251790 100700
rect 301682 100688 301688 100700
rect 251784 100660 301688 100688
rect 251784 100648 251790 100660
rect 301682 100648 301688 100660
rect 301740 100648 301746 100700
rect 324314 100648 324320 100700
rect 324372 100688 324378 100700
rect 345750 100688 345756 100700
rect 324372 100660 345756 100688
rect 324372 100648 324378 100660
rect 345750 100648 345756 100660
rect 345808 100648 345814 100700
rect 452562 100648 452568 100700
rect 452620 100688 452626 100700
rect 477494 100688 477500 100700
rect 452620 100660 477500 100688
rect 452620 100648 452626 100660
rect 477494 100648 477500 100660
rect 477552 100648 477558 100700
rect 252462 100580 252468 100632
rect 252520 100620 252526 100632
rect 279602 100620 279608 100632
rect 252520 100592 279608 100620
rect 252520 100580 252526 100592
rect 279602 100580 279608 100592
rect 279660 100580 279666 100632
rect 252370 100512 252376 100564
rect 252428 100552 252434 100564
rect 270034 100552 270040 100564
rect 252428 100524 270040 100552
rect 252428 100512 252434 100524
rect 270034 100512 270040 100524
rect 270092 100512 270098 100564
rect 374638 99968 374644 100020
rect 374696 100008 374702 100020
rect 397546 100008 397552 100020
rect 374696 99980 397552 100008
rect 374696 99968 374702 99980
rect 397546 99968 397552 99980
rect 397604 99968 397610 100020
rect 192662 99424 192668 99476
rect 192720 99464 192726 99476
rect 213914 99464 213920 99476
rect 192720 99436 213920 99464
rect 192720 99424 192726 99436
rect 213914 99424 213920 99436
rect 213972 99424 213978 99476
rect 303154 99424 303160 99476
rect 303212 99464 303218 99476
rect 307662 99464 307668 99476
rect 303212 99436 307668 99464
rect 303212 99424 303218 99436
rect 307662 99424 307668 99436
rect 307720 99424 307726 99476
rect 167822 99356 167828 99408
rect 167880 99396 167886 99408
rect 214006 99396 214012 99408
rect 167880 99368 214012 99396
rect 167880 99356 167886 99368
rect 214006 99356 214012 99368
rect 214064 99356 214070 99408
rect 297358 99356 297364 99408
rect 297416 99396 297422 99408
rect 307570 99396 307576 99408
rect 297416 99368 307576 99396
rect 297416 99356 297422 99368
rect 307570 99356 307576 99368
rect 307628 99356 307634 99408
rect 576118 99356 576124 99408
rect 576176 99396 576182 99408
rect 580166 99396 580172 99408
rect 576176 99368 580172 99396
rect 576176 99356 576182 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 251542 99288 251548 99340
rect 251600 99328 251606 99340
rect 257614 99328 257620 99340
rect 251600 99300 257620 99328
rect 251600 99288 251606 99300
rect 257614 99288 257620 99300
rect 257672 99288 257678 99340
rect 251818 99152 251824 99204
rect 251876 99192 251882 99204
rect 290550 99192 290556 99204
rect 251876 99164 290556 99192
rect 251876 99152 251882 99164
rect 290550 99152 290556 99164
rect 290608 99152 290614 99204
rect 251174 99084 251180 99136
rect 251232 99124 251238 99136
rect 253382 99124 253388 99136
rect 251232 99096 253388 99124
rect 251232 99084 251238 99096
rect 253382 99084 253388 99096
rect 253440 99084 253446 99136
rect 452286 98880 452292 98932
rect 452344 98920 452350 98932
rect 454034 98920 454040 98932
rect 452344 98892 454040 98920
rect 452344 98880 452350 98892
rect 454034 98880 454040 98892
rect 454092 98880 454098 98932
rect 332594 98608 332600 98660
rect 332652 98648 332658 98660
rect 391934 98648 391940 98660
rect 332652 98620 391940 98648
rect 332652 98608 332658 98620
rect 391934 98608 391940 98620
rect 391992 98608 391998 98660
rect 172054 98064 172060 98116
rect 172112 98104 172118 98116
rect 214006 98104 214012 98116
rect 172112 98076 214012 98104
rect 172112 98064 172118 98076
rect 214006 98064 214012 98076
rect 214064 98064 214070 98116
rect 300302 98064 300308 98116
rect 300360 98104 300366 98116
rect 307570 98104 307576 98116
rect 300360 98076 307576 98104
rect 300360 98064 300366 98076
rect 307570 98064 307576 98076
rect 307628 98064 307634 98116
rect 164878 97996 164884 98048
rect 164936 98036 164942 98048
rect 213914 98036 213920 98048
rect 164936 98008 213920 98036
rect 164936 97996 164942 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 283650 97996 283656 98048
rect 283708 98036 283714 98048
rect 307662 98036 307668 98048
rect 283708 98008 307668 98036
rect 283708 97996 283714 98008
rect 307662 97996 307668 98008
rect 307720 97996 307726 98048
rect 399018 97792 399024 97844
rect 399076 97832 399082 97844
rect 399662 97832 399668 97844
rect 399076 97804 399668 97832
rect 399076 97792 399082 97804
rect 399662 97792 399668 97804
rect 399720 97792 399726 97844
rect 252186 97588 252192 97640
rect 252244 97628 252250 97640
rect 256050 97628 256056 97640
rect 252244 97600 256056 97628
rect 252244 97588 252250 97600
rect 256050 97588 256056 97600
rect 256108 97588 256114 97640
rect 453298 97248 453304 97300
rect 453356 97288 453362 97300
rect 467834 97288 467840 97300
rect 453356 97260 467840 97288
rect 453356 97248 453362 97260
rect 467834 97248 467840 97260
rect 467892 97248 467898 97300
rect 255958 96772 255964 96824
rect 256016 96812 256022 96824
rect 307662 96812 307668 96824
rect 256016 96784 307668 96812
rect 256016 96772 256022 96784
rect 307662 96772 307668 96784
rect 307720 96772 307726 96824
rect 251910 96704 251916 96756
rect 251968 96744 251974 96756
rect 307570 96744 307576 96756
rect 251968 96716 307576 96744
rect 251968 96704 251974 96716
rect 307570 96704 307576 96716
rect 307628 96704 307634 96756
rect 209130 96636 209136 96688
rect 209188 96676 209194 96688
rect 213914 96676 213920 96688
rect 209188 96648 213920 96676
rect 209188 96636 209194 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 249058 96636 249064 96688
rect 249116 96676 249122 96688
rect 307662 96676 307668 96688
rect 249116 96648 307668 96676
rect 249116 96636 249122 96648
rect 307662 96636 307668 96648
rect 307720 96636 307726 96688
rect 356790 96636 356796 96688
rect 356848 96676 356854 96688
rect 397546 96676 397552 96688
rect 356848 96648 397552 96676
rect 356848 96636 356854 96648
rect 397546 96636 397552 96648
rect 397604 96636 397610 96688
rect 174538 96568 174544 96620
rect 174596 96608 174602 96620
rect 321462 96608 321468 96620
rect 174596 96580 321468 96608
rect 174596 96568 174602 96580
rect 321462 96568 321468 96580
rect 321520 96568 321526 96620
rect 299290 95888 299296 95940
rect 299348 95928 299354 95940
rect 314654 95928 314660 95940
rect 299348 95900 314660 95928
rect 299348 95888 299354 95900
rect 314654 95888 314660 95900
rect 314712 95888 314718 95940
rect 378042 95276 378048 95328
rect 378100 95316 378106 95328
rect 419350 95316 419356 95328
rect 378100 95288 419356 95316
rect 378100 95276 378106 95288
rect 419350 95276 419356 95288
rect 419408 95276 419414 95328
rect 441890 95276 441896 95328
rect 441948 95316 441954 95328
rect 460934 95316 460940 95328
rect 441948 95288 460940 95316
rect 441948 95276 441954 95288
rect 460934 95276 460940 95288
rect 460992 95276 460998 95328
rect 211154 95208 211160 95260
rect 211212 95248 211218 95260
rect 213914 95248 213920 95260
rect 211212 95220 213920 95248
rect 211212 95208 211218 95220
rect 213914 95208 213920 95220
rect 213972 95208 213978 95260
rect 298922 95208 298928 95260
rect 298980 95248 298986 95260
rect 307662 95248 307668 95260
rect 298980 95220 307668 95248
rect 298980 95208 298986 95220
rect 307662 95208 307668 95220
rect 307720 95208 307726 95260
rect 342898 95208 342904 95260
rect 342956 95248 342962 95260
rect 400674 95248 400680 95260
rect 342956 95220 400680 95248
rect 342956 95208 342962 95220
rect 400674 95208 400680 95220
rect 400732 95208 400738 95260
rect 448974 95208 448980 95260
rect 449032 95248 449038 95260
rect 480346 95248 480352 95260
rect 449032 95220 480352 95248
rect 449032 95208 449038 95220
rect 480346 95208 480352 95220
rect 480404 95208 480410 95260
rect 193858 95140 193864 95192
rect 193916 95180 193922 95192
rect 322934 95180 322940 95192
rect 193916 95152 322940 95180
rect 193916 95140 193922 95152
rect 322934 95140 322940 95152
rect 322992 95140 322998 95192
rect 356698 95140 356704 95192
rect 356756 95180 356762 95192
rect 422570 95180 422576 95192
rect 356756 95152 422576 95180
rect 356756 95140 356762 95152
rect 422570 95140 422576 95152
rect 422628 95140 422634 95192
rect 438670 95140 438676 95192
rect 438728 95180 438734 95192
rect 525058 95180 525064 95192
rect 438728 95152 525064 95180
rect 438728 95140 438734 95152
rect 525058 95140 525064 95152
rect 525116 95140 525122 95192
rect 202138 95072 202144 95124
rect 202196 95112 202202 95124
rect 321646 95112 321652 95124
rect 202196 95084 321652 95112
rect 202196 95072 202202 95084
rect 321646 95072 321652 95084
rect 321704 95072 321710 95124
rect 368290 95072 368296 95124
rect 368348 95112 368354 95124
rect 447042 95112 447048 95124
rect 368348 95084 447048 95112
rect 368348 95072 368354 95084
rect 447042 95072 447048 95084
rect 447100 95072 447106 95124
rect 63402 95004 63408 95056
rect 63460 95044 63466 95056
rect 196802 95044 196808 95056
rect 63460 95016 196808 95044
rect 63460 95004 63466 95016
rect 196802 95004 196808 95016
rect 196860 95004 196866 95056
rect 276658 95004 276664 95056
rect 276716 95044 276722 95056
rect 325694 95044 325700 95056
rect 276716 95016 325700 95044
rect 276716 95004 276722 95016
rect 325694 95004 325700 95016
rect 325752 95044 325758 95056
rect 326338 95044 326344 95056
rect 325752 95016 326344 95044
rect 325752 95004 325758 95016
rect 326338 95004 326344 95016
rect 326396 95004 326402 95056
rect 371970 95004 371976 95056
rect 372028 95044 372034 95056
rect 430942 95044 430948 95056
rect 372028 95016 430948 95044
rect 372028 95004 372034 95016
rect 430942 95004 430948 95016
rect 431000 95004 431006 95056
rect 438118 95004 438124 95056
rect 438176 95044 438182 95056
rect 438670 95044 438676 95056
rect 438176 95016 438676 95044
rect 438176 95004 438182 95016
rect 438670 95004 438676 95016
rect 438728 95004 438734 95056
rect 438762 95004 438768 95056
rect 438820 95044 438826 95056
rect 459646 95044 459652 95056
rect 438820 95016 459652 95044
rect 438820 95004 438826 95016
rect 459646 95004 459652 95016
rect 459704 95004 459710 95056
rect 436738 94936 436744 94988
rect 436796 94976 436802 94988
rect 463694 94976 463700 94988
rect 436796 94948 463700 94976
rect 436796 94936 436802 94948
rect 463694 94936 463700 94948
rect 463752 94936 463758 94988
rect 425790 94868 425796 94920
rect 425848 94908 425854 94920
rect 458818 94908 458824 94920
rect 425848 94880 458824 94908
rect 425848 94868 425854 94880
rect 458818 94868 458824 94880
rect 458876 94868 458882 94920
rect 395798 94800 395804 94852
rect 395856 94840 395862 94852
rect 395856 94812 431954 94840
rect 395856 94800 395862 94812
rect 431926 94772 431954 94812
rect 432230 94800 432236 94852
rect 432288 94840 432294 94852
rect 438762 94840 438768 94852
rect 432288 94812 438768 94840
rect 432288 94800 432294 94812
rect 438762 94800 438768 94812
rect 438820 94800 438826 94852
rect 441246 94772 441252 94784
rect 431926 94744 441252 94772
rect 441246 94732 441252 94744
rect 441304 94732 441310 94784
rect 317414 94460 317420 94512
rect 317472 94500 317478 94512
rect 344278 94500 344284 94512
rect 317472 94472 344284 94500
rect 317472 94460 317478 94472
rect 344278 94460 344284 94472
rect 344336 94460 344342 94512
rect 115842 94052 115848 94104
rect 115900 94092 115906 94104
rect 169294 94092 169300 94104
rect 115900 94064 169300 94092
rect 115900 94052 115906 94064
rect 169294 94052 169300 94064
rect 169352 94052 169358 94104
rect 113174 93984 113180 94036
rect 113232 94024 113238 94036
rect 181438 94024 181444 94036
rect 113232 93996 181444 94024
rect 113232 93984 113238 93996
rect 181438 93984 181444 93996
rect 181496 93984 181502 94036
rect 126514 93916 126520 93968
rect 126572 93956 126578 93968
rect 200758 93956 200764 93968
rect 126572 93928 200764 93956
rect 126572 93916 126578 93928
rect 200758 93916 200764 93928
rect 200816 93916 200822 93968
rect 94958 93848 94964 93900
rect 95016 93888 95022 93900
rect 170674 93888 170680 93900
rect 95016 93860 170680 93888
rect 95016 93848 95022 93860
rect 170674 93848 170680 93860
rect 170732 93848 170738 93900
rect 66162 93780 66168 93832
rect 66220 93820 66226 93832
rect 198182 93820 198188 93832
rect 66220 93792 198188 93820
rect 66220 93780 66226 93792
rect 198182 93780 198188 93792
rect 198240 93780 198246 93832
rect 308398 93780 308404 93832
rect 308456 93820 308462 93832
rect 321738 93820 321744 93832
rect 308456 93792 321744 93820
rect 308456 93780 308462 93792
rect 321738 93780 321744 93792
rect 321796 93780 321802 93832
rect 353294 93780 353300 93832
rect 353352 93820 353358 93832
rect 387242 93820 387248 93832
rect 353352 93792 387248 93820
rect 353352 93780 353358 93792
rect 387242 93780 387248 93792
rect 387300 93780 387306 93832
rect 399478 93780 399484 93832
rect 399536 93820 399542 93832
rect 405182 93820 405188 93832
rect 399536 93792 405188 93820
rect 399536 93780 399542 93792
rect 405182 93780 405188 93792
rect 405240 93780 405246 93832
rect 447686 93780 447692 93832
rect 447744 93820 447750 93832
rect 476114 93820 476120 93832
rect 447744 93792 476120 93820
rect 447744 93780 447750 93792
rect 476114 93780 476120 93792
rect 476172 93780 476178 93832
rect 387150 93712 387156 93764
rect 387208 93752 387214 93764
rect 416774 93752 416780 93764
rect 387208 93724 416780 93752
rect 387208 93712 387214 93724
rect 416774 93712 416780 93724
rect 416832 93712 416838 93764
rect 417418 93712 417424 93764
rect 417476 93752 417482 93764
rect 458174 93752 458180 93764
rect 417476 93724 458180 93752
rect 417476 93712 417482 93724
rect 458174 93712 458180 93724
rect 458232 93712 458238 93764
rect 391198 93644 391204 93696
rect 391256 93684 391262 93696
rect 407114 93684 407120 93696
rect 391256 93656 407120 93684
rect 391256 93644 391262 93656
rect 407114 93644 407120 93656
rect 407172 93644 407178 93696
rect 423858 93644 423864 93696
rect 423916 93684 423922 93696
rect 456794 93684 456800 93696
rect 423916 93656 456800 93684
rect 423916 93644 423922 93656
rect 456794 93644 456800 93656
rect 456852 93644 456858 93696
rect 393958 93576 393964 93628
rect 394016 93616 394022 93628
rect 403250 93616 403256 93628
rect 394016 93588 403256 93616
rect 394016 93576 394022 93588
rect 403250 93576 403256 93588
rect 403308 93576 403314 93628
rect 435358 93576 435364 93628
rect 435416 93616 435422 93628
rect 457438 93616 457444 93628
rect 435416 93588 457444 93616
rect 435416 93576 435422 93588
rect 457438 93576 457444 93588
rect 457496 93576 457502 93628
rect 382918 93508 382924 93560
rect 382976 93548 382982 93560
rect 440602 93548 440608 93560
rect 382976 93520 440608 93548
rect 382976 93508 382982 93520
rect 440602 93508 440608 93520
rect 440660 93508 440666 93560
rect 443178 93508 443184 93560
rect 443236 93548 443242 93560
rect 459738 93548 459744 93560
rect 443236 93520 459744 93548
rect 443236 93508 443242 93520
rect 459738 93508 459744 93520
rect 459796 93508 459802 93560
rect 130746 93372 130752 93424
rect 130804 93412 130810 93424
rect 171778 93412 171784 93424
rect 130804 93384 171784 93412
rect 130804 93372 130810 93384
rect 171778 93372 171784 93384
rect 171836 93372 171842 93424
rect 151722 93304 151728 93356
rect 151780 93344 151786 93356
rect 195238 93344 195244 93356
rect 151780 93316 195244 93344
rect 151780 93304 151786 93316
rect 195238 93304 195244 93316
rect 195296 93304 195302 93356
rect 113818 93236 113824 93288
rect 113876 93276 113882 93288
rect 173342 93276 173348 93288
rect 113876 93248 173348 93276
rect 113876 93236 113882 93248
rect 173342 93236 173348 93248
rect 173400 93236 173406 93288
rect 97258 93168 97264 93220
rect 97316 93208 97322 93220
rect 174722 93208 174728 93220
rect 97316 93180 174728 93208
rect 97316 93168 97322 93180
rect 174722 93168 174728 93180
rect 174780 93168 174786 93220
rect 121454 93100 121460 93152
rect 121512 93140 121518 93152
rect 214926 93140 214932 93152
rect 121512 93112 214932 93140
rect 121512 93100 121518 93112
rect 214926 93100 214932 93112
rect 214984 93100 214990 93152
rect 318794 93100 318800 93152
rect 318852 93140 318858 93152
rect 353294 93140 353300 93152
rect 318852 93112 353300 93140
rect 318852 93100 318858 93112
rect 353294 93100 353300 93112
rect 353352 93100 353358 93152
rect 416774 92828 416780 92880
rect 416832 92868 416838 92880
rect 418062 92868 418068 92880
rect 416832 92840 418068 92868
rect 416832 92828 416838 92840
rect 418062 92828 418068 92840
rect 418120 92828 418126 92880
rect 418890 92488 418896 92540
rect 418948 92528 418954 92540
rect 420638 92528 420644 92540
rect 418948 92500 420644 92528
rect 418948 92488 418954 92500
rect 420638 92488 420644 92500
rect 420696 92488 420702 92540
rect 422938 92488 422944 92540
rect 422996 92528 423002 92540
rect 424502 92528 424508 92540
rect 422996 92500 424508 92528
rect 422996 92488 423002 92500
rect 424502 92488 424508 92500
rect 424560 92488 424566 92540
rect 447778 92488 447784 92540
rect 447836 92528 447842 92540
rect 449618 92528 449624 92540
rect 447836 92500 449624 92528
rect 447836 92488 447842 92500
rect 449618 92488 449624 92500
rect 449676 92488 449682 92540
rect 98178 92420 98184 92472
rect 98236 92460 98242 92472
rect 121454 92460 121460 92472
rect 98236 92432 121460 92460
rect 98236 92420 98242 92432
rect 121454 92420 121460 92432
rect 121512 92420 121518 92472
rect 125778 92420 125784 92472
rect 125836 92460 125842 92472
rect 189718 92460 189724 92472
rect 125836 92432 189724 92460
rect 125836 92420 125842 92432
rect 189718 92420 189724 92432
rect 189776 92420 189782 92472
rect 192478 92420 192484 92472
rect 192536 92460 192542 92472
rect 321554 92460 321560 92472
rect 192536 92432 321560 92460
rect 192536 92420 192542 92432
rect 321554 92420 321560 92432
rect 321612 92420 321618 92472
rect 382182 92420 382188 92472
rect 382240 92460 382246 92472
rect 410978 92460 410984 92472
rect 382240 92432 410984 92460
rect 382240 92420 382246 92432
rect 410978 92420 410984 92432
rect 411036 92420 411042 92472
rect 120350 92352 120356 92404
rect 120408 92392 120414 92404
rect 182910 92392 182916 92404
rect 120408 92364 182916 92392
rect 120408 92352 120414 92364
rect 182910 92352 182916 92364
rect 182968 92352 182974 92404
rect 404538 92352 404544 92404
rect 404596 92392 404602 92404
rect 462314 92392 462320 92404
rect 404596 92364 462320 92392
rect 404596 92352 404602 92364
rect 462314 92352 462320 92364
rect 462372 92352 462378 92404
rect 116762 92284 116768 92336
rect 116820 92324 116826 92336
rect 171870 92324 171876 92336
rect 116820 92296 171876 92324
rect 116820 92284 116826 92296
rect 171870 92284 171876 92296
rect 171928 92284 171934 92336
rect 375282 92284 375288 92336
rect 375340 92324 375346 92336
rect 416130 92324 416136 92336
rect 375340 92296 416136 92324
rect 375340 92284 375346 92296
rect 416130 92284 416136 92296
rect 416188 92284 416194 92336
rect 432874 92284 432880 92336
rect 432932 92324 432938 92336
rect 461026 92324 461032 92336
rect 432932 92296 461032 92324
rect 432932 92284 432938 92296
rect 461026 92284 461032 92296
rect 461084 92284 461090 92336
rect 152090 92216 152096 92268
rect 152148 92256 152154 92268
rect 191098 92256 191104 92268
rect 152148 92228 191104 92256
rect 152148 92216 152154 92228
rect 191098 92216 191104 92228
rect 191156 92216 191162 92268
rect 386322 92216 386328 92268
rect 386380 92256 386386 92268
rect 405734 92256 405740 92268
rect 386380 92228 405740 92256
rect 386380 92216 386386 92228
rect 405734 92216 405740 92228
rect 405792 92216 405798 92268
rect 407114 92216 407120 92268
rect 407172 92256 407178 92268
rect 576118 92256 576124 92268
rect 407172 92228 576124 92256
rect 407172 92216 407178 92228
rect 576118 92216 576124 92228
rect 576176 92216 576182 92268
rect 133138 92148 133144 92200
rect 133196 92188 133202 92200
rect 167914 92188 167920 92200
rect 133196 92160 167920 92188
rect 133196 92148 133202 92160
rect 167914 92148 167920 92160
rect 167972 92148 167978 92200
rect 135714 92080 135720 92132
rect 135772 92120 135778 92132
rect 166534 92120 166540 92132
rect 135772 92092 166540 92120
rect 135772 92080 135778 92092
rect 166534 92080 166540 92092
rect 166592 92080 166598 92132
rect 405734 91740 405740 91792
rect 405792 91780 405798 91792
rect 406470 91780 406476 91792
rect 405792 91752 406476 91780
rect 405792 91740 405798 91752
rect 406470 91740 406476 91752
rect 406528 91740 406534 91792
rect 107378 91196 107384 91248
rect 107436 91236 107442 91248
rect 119338 91236 119344 91248
rect 107436 91208 119344 91236
rect 107436 91196 107442 91208
rect 119338 91196 119344 91208
rect 119396 91196 119402 91248
rect 98638 91128 98644 91180
rect 98696 91168 98702 91180
rect 116578 91168 116584 91180
rect 98696 91140 116584 91168
rect 98696 91128 98702 91140
rect 116578 91128 116584 91140
rect 116636 91128 116642 91180
rect 87138 91060 87144 91112
rect 87196 91100 87202 91112
rect 134518 91100 134524 91112
rect 87196 91072 134524 91100
rect 87196 91060 87202 91072
rect 134518 91060 134524 91072
rect 134576 91060 134582 91112
rect 416130 91060 416136 91112
rect 416188 91100 416194 91112
rect 418982 91100 418988 91112
rect 416188 91072 418988 91100
rect 416188 91060 416194 91072
rect 418982 91060 418988 91072
rect 419040 91060 419046 91112
rect 67266 90992 67272 91044
rect 67324 91032 67330 91044
rect 214558 91032 214564 91044
rect 67324 91004 214564 91032
rect 67324 90992 67330 91004
rect 214558 90992 214564 91004
rect 214616 90992 214622 91044
rect 369762 90992 369768 91044
rect 369820 91032 369826 91044
rect 437382 91032 437388 91044
rect 369820 91004 437388 91032
rect 369820 90992 369826 91004
rect 437382 90992 437388 91004
rect 437440 90992 437446 91044
rect 67450 90924 67456 90976
rect 67508 90964 67514 90976
rect 209038 90964 209044 90976
rect 67508 90936 209044 90964
rect 67508 90924 67514 90936
rect 209038 90924 209044 90936
rect 209096 90924 209102 90976
rect 340874 90924 340880 90976
rect 340932 90964 340938 90976
rect 398190 90964 398196 90976
rect 340932 90936 398196 90964
rect 340932 90924 340938 90936
rect 398190 90924 398196 90936
rect 398248 90924 398254 90976
rect 415486 90924 415492 90976
rect 415544 90964 415550 90976
rect 416682 90964 416688 90976
rect 415544 90936 416688 90964
rect 415544 90924 415550 90936
rect 416682 90924 416688 90936
rect 416740 90964 416746 90976
rect 462406 90964 462412 90976
rect 416740 90936 462412 90964
rect 416740 90924 416746 90936
rect 462406 90924 462412 90936
rect 462464 90924 462470 90976
rect 129458 90856 129464 90908
rect 129516 90896 129522 90908
rect 192570 90896 192576 90908
rect 129516 90868 192576 90896
rect 129516 90856 129522 90868
rect 192570 90856 192576 90868
rect 192628 90856 192634 90908
rect 426434 90856 426440 90908
rect 426492 90896 426498 90908
rect 427722 90896 427728 90908
rect 426492 90868 427728 90896
rect 426492 90856 426498 90868
rect 427722 90856 427728 90868
rect 427780 90896 427786 90908
rect 470686 90896 470692 90908
rect 427780 90868 470692 90896
rect 427780 90856 427786 90868
rect 470686 90856 470692 90868
rect 470744 90856 470750 90908
rect 110138 90788 110144 90840
rect 110196 90828 110202 90840
rect 169202 90828 169208 90840
rect 110196 90800 169208 90828
rect 110196 90788 110202 90800
rect 169202 90788 169208 90800
rect 169260 90788 169266 90840
rect 124030 90720 124036 90772
rect 124088 90760 124094 90772
rect 171962 90760 171968 90772
rect 124088 90732 171968 90760
rect 124088 90720 124094 90732
rect 171962 90720 171968 90732
rect 172020 90720 172026 90772
rect 151538 90652 151544 90704
rect 151596 90692 151602 90704
rect 185578 90692 185584 90704
rect 151596 90664 185584 90692
rect 151596 90652 151602 90664
rect 185578 90652 185584 90664
rect 185636 90652 185642 90704
rect 216582 90380 216588 90432
rect 216640 90420 216646 90432
rect 317506 90420 317512 90432
rect 216640 90392 317512 90420
rect 216640 90380 216646 90392
rect 317506 90380 317512 90392
rect 317564 90380 317570 90432
rect 192478 90312 192484 90364
rect 192536 90352 192542 90364
rect 307294 90352 307300 90364
rect 192536 90324 307300 90352
rect 192536 90312 192542 90324
rect 307294 90312 307300 90324
rect 307352 90312 307358 90364
rect 311158 90312 311164 90364
rect 311216 90352 311222 90364
rect 340874 90352 340880 90364
rect 311216 90324 340880 90352
rect 311216 90312 311222 90324
rect 340874 90312 340880 90324
rect 340932 90312 340938 90364
rect 403618 90312 403624 90364
rect 403676 90352 403682 90364
rect 428366 90352 428372 90364
rect 403676 90324 428372 90352
rect 403676 90312 403682 90324
rect 428366 90312 428372 90324
rect 428424 90312 428430 90364
rect 66070 89632 66076 89684
rect 66128 89672 66134 89684
rect 209130 89672 209136 89684
rect 66128 89644 209136 89672
rect 66128 89632 66134 89644
rect 209130 89632 209136 89644
rect 209188 89632 209194 89684
rect 409138 89632 409144 89684
rect 409196 89672 409202 89684
rect 500218 89672 500224 89684
rect 409196 89644 500224 89672
rect 409196 89632 409202 89644
rect 500218 89632 500224 89644
rect 500276 89632 500282 89684
rect 117130 89564 117136 89616
rect 117188 89604 117194 89616
rect 206462 89604 206468 89616
rect 117188 89576 206468 89604
rect 117188 89564 117194 89576
rect 206462 89564 206468 89576
rect 206520 89564 206526 89616
rect 413554 89564 413560 89616
rect 413612 89604 413618 89616
rect 467926 89604 467932 89616
rect 413612 89576 467932 89604
rect 413612 89564 413618 89576
rect 467926 89564 467932 89576
rect 467984 89564 467990 89616
rect 99742 89496 99748 89548
rect 99800 89536 99806 89548
rect 173434 89536 173440 89548
rect 99800 89508 173440 89536
rect 99800 89496 99806 89508
rect 173434 89496 173440 89508
rect 173492 89496 173498 89548
rect 110322 89428 110328 89480
rect 110380 89468 110386 89480
rect 181530 89468 181536 89480
rect 110380 89440 181536 89468
rect 110380 89428 110386 89440
rect 181530 89428 181536 89440
rect 181588 89428 181594 89480
rect 151354 89360 151360 89412
rect 151412 89400 151418 89412
rect 204898 89400 204904 89412
rect 151412 89372 204904 89400
rect 151412 89360 151418 89372
rect 204898 89360 204904 89372
rect 204956 89360 204962 89412
rect 132218 89292 132224 89344
rect 132276 89332 132282 89344
rect 166258 89332 166264 89344
rect 132276 89304 166264 89332
rect 132276 89292 132282 89304
rect 166258 89292 166264 89304
rect 166316 89292 166322 89344
rect 310514 88952 310520 89004
rect 310572 88992 310578 89004
rect 397454 88992 397460 89004
rect 310572 88964 397460 88992
rect 310572 88952 310578 88964
rect 397454 88952 397460 88964
rect 397512 88952 397518 89004
rect 408494 88952 408500 89004
rect 408552 88992 408558 89004
rect 409690 88992 409696 89004
rect 408552 88964 409696 88992
rect 408552 88952 408558 88964
rect 409690 88952 409696 88964
rect 409748 88952 409754 89004
rect 427814 88952 427820 89004
rect 427872 88992 427878 89004
rect 429010 88992 429016 89004
rect 427872 88964 429016 88992
rect 427872 88952 427878 88964
rect 429010 88952 429016 88964
rect 429068 88952 429074 89004
rect 75362 88272 75368 88324
rect 75420 88312 75426 88324
rect 211154 88312 211160 88324
rect 75420 88284 211160 88312
rect 75420 88272 75426 88284
rect 211154 88272 211160 88284
rect 211212 88272 211218 88324
rect 401594 88272 401600 88324
rect 401652 88312 401658 88324
rect 402606 88312 402612 88324
rect 401652 88284 402612 88312
rect 401652 88272 401658 88284
rect 402606 88272 402612 88284
rect 402664 88312 402670 88324
rect 549254 88312 549260 88324
rect 402664 88284 549260 88312
rect 402664 88272 402670 88284
rect 549254 88272 549260 88284
rect 549312 88272 549318 88324
rect 86402 88204 86408 88256
rect 86460 88244 86466 88256
rect 164878 88244 164884 88256
rect 86460 88216 164884 88244
rect 86460 88204 86466 88216
rect 164878 88204 164884 88216
rect 164936 88204 164942 88256
rect 316034 88204 316040 88256
rect 316092 88244 316098 88256
rect 454218 88244 454224 88256
rect 316092 88216 454224 88244
rect 316092 88204 316098 88216
rect 454218 88204 454224 88216
rect 454276 88204 454282 88256
rect 105722 88136 105728 88188
rect 105780 88176 105786 88188
rect 184290 88176 184296 88188
rect 105780 88148 184296 88176
rect 105780 88136 105786 88148
rect 184290 88136 184296 88148
rect 184348 88136 184354 88188
rect 400858 88136 400864 88188
rect 400916 88176 400922 88188
rect 401318 88176 401324 88188
rect 400916 88148 401324 88176
rect 400916 88136 400922 88148
rect 401318 88136 401324 88148
rect 401376 88176 401382 88188
rect 494054 88176 494060 88188
rect 401376 88148 494060 88176
rect 401376 88136 401382 88148
rect 494054 88136 494060 88148
rect 494112 88136 494118 88188
rect 134794 88068 134800 88120
rect 134852 88108 134858 88120
rect 188338 88108 188344 88120
rect 134852 88080 188344 88108
rect 134852 88068 134858 88080
rect 188338 88068 188344 88080
rect 188396 88068 188402 88120
rect 119890 88000 119896 88052
rect 119948 88040 119954 88052
rect 169018 88040 169024 88052
rect 119948 88012 169024 88040
rect 119948 88000 119954 88012
rect 169018 88000 169024 88012
rect 169076 88000 169082 88052
rect 121362 87932 121368 87984
rect 121420 87972 121426 87984
rect 166350 87972 166356 87984
rect 121420 87944 166356 87972
rect 121420 87932 121426 87944
rect 166350 87932 166356 87944
rect 166408 87932 166414 87984
rect 179230 87592 179236 87644
rect 179288 87632 179294 87644
rect 267826 87632 267832 87644
rect 179288 87604 267832 87632
rect 179288 87592 179294 87604
rect 267826 87592 267832 87604
rect 267884 87632 267890 87644
rect 355318 87632 355324 87644
rect 267884 87604 355324 87632
rect 267884 87592 267890 87604
rect 355318 87592 355324 87604
rect 355376 87592 355382 87644
rect 62022 86912 62028 86964
rect 62080 86952 62086 86964
rect 189810 86952 189816 86964
rect 62080 86924 189816 86952
rect 62080 86912 62086 86924
rect 189810 86912 189816 86924
rect 189868 86912 189874 86964
rect 416682 86912 416688 86964
rect 416740 86952 416746 86964
rect 418798 86952 418804 86964
rect 416740 86924 418804 86952
rect 416740 86912 416746 86924
rect 418798 86912 418804 86924
rect 418856 86912 418862 86964
rect 418982 86912 418988 86964
rect 419040 86952 419046 86964
rect 580166 86952 580172 86964
rect 419040 86924 580172 86952
rect 419040 86912 419046 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 112438 86844 112444 86896
rect 112496 86884 112502 86896
rect 211890 86884 211896 86896
rect 112496 86856 211896 86884
rect 112496 86844 112502 86856
rect 211890 86844 211896 86856
rect 211948 86844 211954 86896
rect 103330 86776 103336 86828
rect 103388 86816 103394 86828
rect 184198 86816 184204 86828
rect 103388 86788 184204 86816
rect 103388 86776 103394 86788
rect 184198 86776 184204 86788
rect 184256 86776 184262 86828
rect 118050 86708 118056 86760
rect 118108 86748 118114 86760
rect 193950 86748 193956 86760
rect 118108 86720 193956 86748
rect 118108 86708 118114 86720
rect 193950 86708 193956 86720
rect 194008 86708 194014 86760
rect 102962 86640 102968 86692
rect 103020 86680 103026 86692
rect 173250 86680 173256 86692
rect 103020 86652 173256 86680
rect 103020 86640 103026 86652
rect 173250 86640 173256 86652
rect 173308 86640 173314 86692
rect 122834 86572 122840 86624
rect 122892 86612 122898 86624
rect 167638 86612 167644 86624
rect 122892 86584 167644 86612
rect 122892 86572 122898 86584
rect 167638 86572 167644 86584
rect 167696 86572 167702 86624
rect 299382 86300 299388 86352
rect 299440 86340 299446 86352
rect 320818 86340 320824 86352
rect 299440 86312 320824 86340
rect 299440 86300 299446 86312
rect 320818 86300 320824 86312
rect 320876 86300 320882 86352
rect 328454 86300 328460 86352
rect 328512 86340 328518 86352
rect 374638 86340 374644 86352
rect 328512 86312 374644 86340
rect 328512 86300 328518 86312
rect 374638 86300 374644 86312
rect 374696 86300 374702 86352
rect 242894 86232 242900 86284
rect 242952 86272 242958 86284
rect 294046 86272 294052 86284
rect 242952 86244 294052 86272
rect 242952 86232 242958 86244
rect 294046 86232 294052 86244
rect 294104 86232 294110 86284
rect 312538 86232 312544 86284
rect 312596 86272 312602 86284
rect 401594 86272 401600 86284
rect 312596 86244 401600 86272
rect 312596 86232 312602 86244
rect 401594 86232 401600 86244
rect 401652 86232 401658 86284
rect 67542 85484 67548 85536
rect 67600 85524 67606 85536
rect 191190 85524 191196 85536
rect 67600 85496 191196 85524
rect 67600 85484 67606 85496
rect 191190 85484 191196 85496
rect 191248 85484 191254 85536
rect 90634 85416 90640 85468
rect 90692 85456 90698 85468
rect 211982 85456 211988 85468
rect 90692 85428 211988 85456
rect 90692 85416 90698 85428
rect 211982 85416 211988 85428
rect 212040 85416 212046 85468
rect 111058 85348 111064 85400
rect 111116 85388 111122 85400
rect 174630 85388 174636 85400
rect 111116 85360 174636 85388
rect 111116 85348 111122 85360
rect 174630 85348 174636 85360
rect 174688 85348 174694 85400
rect 121914 85280 121920 85332
rect 121972 85320 121978 85332
rect 183002 85320 183008 85332
rect 121972 85292 183008 85320
rect 121972 85280 121978 85292
rect 183002 85280 183008 85292
rect 183060 85280 183066 85332
rect 2774 85212 2780 85264
rect 2832 85252 2838 85264
rect 4798 85252 4804 85264
rect 2832 85224 4804 85252
rect 2832 85212 2838 85224
rect 4798 85212 4804 85224
rect 4856 85212 4862 85264
rect 115290 85212 115296 85264
rect 115348 85252 115354 85264
rect 167730 85252 167736 85264
rect 115348 85224 167736 85252
rect 115348 85212 115354 85224
rect 167730 85212 167736 85224
rect 167788 85212 167794 85264
rect 104710 84124 104716 84176
rect 104768 84164 104774 84176
rect 213270 84164 213276 84176
rect 104768 84136 213276 84164
rect 104768 84124 104774 84136
rect 213270 84124 213276 84136
rect 213328 84124 213334 84176
rect 313734 84124 313740 84176
rect 313792 84164 313798 84176
rect 466546 84164 466552 84176
rect 313792 84136 466552 84164
rect 313792 84124 313798 84136
rect 466546 84124 466552 84136
rect 466604 84124 466610 84176
rect 101950 84056 101956 84108
rect 102008 84096 102014 84108
rect 202322 84096 202328 84108
rect 102008 84068 202328 84096
rect 102008 84056 102014 84068
rect 202322 84056 202328 84068
rect 202380 84056 202386 84108
rect 96522 83988 96528 84040
rect 96580 84028 96586 84040
rect 170582 84028 170588 84040
rect 96580 84000 170588 84028
rect 96580 83988 96586 84000
rect 170582 83988 170588 84000
rect 170640 83988 170646 84040
rect 95142 83920 95148 83972
rect 95200 83960 95206 83972
rect 166442 83960 166448 83972
rect 95200 83932 166448 83960
rect 95200 83920 95206 83932
rect 166442 83920 166448 83932
rect 166500 83920 166506 83972
rect 118602 83852 118608 83904
rect 118660 83892 118666 83904
rect 189902 83892 189908 83904
rect 118660 83864 189908 83892
rect 118660 83852 118666 83864
rect 189902 83852 189908 83864
rect 189960 83852 189966 83904
rect 125410 83784 125416 83836
rect 125468 83824 125474 83836
rect 196618 83824 196624 83836
rect 125468 83796 196624 83824
rect 125468 83784 125474 83796
rect 196618 83784 196624 83796
rect 196676 83784 196682 83836
rect 238018 83512 238024 83564
rect 238076 83552 238082 83564
rect 251266 83552 251272 83564
rect 238076 83524 251272 83552
rect 238076 83512 238082 83524
rect 251266 83512 251272 83524
rect 251324 83512 251330 83564
rect 199378 83444 199384 83496
rect 199436 83484 199442 83496
rect 271138 83484 271144 83496
rect 199436 83456 271144 83484
rect 199436 83444 199442 83456
rect 271138 83444 271144 83456
rect 271196 83444 271202 83496
rect 313274 82832 313280 82884
rect 313332 82872 313338 82884
rect 313734 82872 313740 82884
rect 313332 82844 313740 82872
rect 313332 82832 313338 82844
rect 313734 82832 313740 82844
rect 313792 82832 313798 82884
rect 64782 82764 64788 82816
rect 64840 82804 64846 82816
rect 308398 82804 308404 82816
rect 64840 82776 308404 82804
rect 64840 82764 64846 82776
rect 308398 82764 308404 82776
rect 308456 82764 308462 82816
rect 108850 82696 108856 82748
rect 108908 82736 108914 82748
rect 207658 82736 207664 82748
rect 108908 82708 207664 82736
rect 108908 82696 108914 82708
rect 207658 82696 207664 82708
rect 207716 82696 207722 82748
rect 238754 82696 238760 82748
rect 238812 82736 238818 82748
rect 295334 82736 295340 82748
rect 238812 82708 295340 82736
rect 238812 82696 238818 82708
rect 295334 82696 295340 82708
rect 295392 82736 295398 82748
rect 450170 82736 450176 82748
rect 295392 82708 450176 82736
rect 295392 82696 295398 82708
rect 450170 82696 450176 82708
rect 450228 82696 450234 82748
rect 125502 82628 125508 82680
rect 125560 82668 125566 82680
rect 203610 82668 203616 82680
rect 125560 82640 203616 82668
rect 125560 82628 125566 82640
rect 203610 82628 203616 82640
rect 203668 82628 203674 82680
rect 108942 82560 108948 82612
rect 109000 82600 109006 82612
rect 185670 82600 185676 82612
rect 109000 82572 185676 82600
rect 109000 82560 109006 82572
rect 185670 82560 185676 82572
rect 185728 82560 185734 82612
rect 97902 82492 97908 82544
rect 97960 82532 97966 82544
rect 170490 82532 170496 82544
rect 97960 82504 170496 82532
rect 97960 82492 97966 82504
rect 170490 82492 170496 82504
rect 170548 82492 170554 82544
rect 93762 81336 93768 81388
rect 93820 81376 93826 81388
rect 204990 81376 204996 81388
rect 93820 81348 204996 81376
rect 93820 81336 93826 81348
rect 204990 81336 204996 81348
rect 205048 81336 205054 81388
rect 126882 81268 126888 81320
rect 126940 81308 126946 81320
rect 211798 81308 211804 81320
rect 126940 81280 211804 81308
rect 126940 81268 126946 81280
rect 211798 81268 211804 81280
rect 211856 81268 211862 81320
rect 111702 81200 111708 81252
rect 111760 81240 111766 81252
rect 188430 81240 188436 81252
rect 111760 81212 188436 81240
rect 111760 81200 111766 81212
rect 188430 81200 188436 81212
rect 188488 81200 188494 81252
rect 100662 81132 100668 81184
rect 100720 81172 100726 81184
rect 169110 81172 169116 81184
rect 100720 81144 169116 81172
rect 100720 81132 100726 81144
rect 169110 81132 169116 81144
rect 169168 81132 169174 81184
rect 107470 81064 107476 81116
rect 107528 81104 107534 81116
rect 173158 81104 173164 81116
rect 107528 81076 173164 81104
rect 107528 81064 107534 81076
rect 173158 81064 173164 81076
rect 173216 81064 173222 81116
rect 185578 80656 185584 80708
rect 185636 80696 185642 80708
rect 307202 80696 307208 80708
rect 185636 80668 307208 80696
rect 185636 80656 185642 80668
rect 307202 80656 307208 80668
rect 307260 80656 307266 80708
rect 336826 80656 336832 80708
rect 336884 80696 336890 80708
rect 427814 80696 427820 80708
rect 336884 80668 427820 80696
rect 336884 80656 336890 80668
rect 427814 80656 427820 80668
rect 427872 80656 427878 80708
rect 92382 79976 92388 80028
rect 92440 80016 92446 80028
rect 194042 80016 194048 80028
rect 92440 79988 194048 80016
rect 92440 79976 92446 79988
rect 194042 79976 194048 79988
rect 194100 79976 194106 80028
rect 309778 79976 309784 80028
rect 309836 80016 309842 80028
rect 310422 80016 310428 80028
rect 309836 79988 310428 80016
rect 309836 79976 309842 79988
rect 310422 79976 310428 79988
rect 310480 80016 310486 80028
rect 419626 80016 419632 80028
rect 310480 79988 419632 80016
rect 310480 79976 310486 79988
rect 419626 79976 419632 79988
rect 419684 79976 419690 80028
rect 115842 79908 115848 79960
rect 115900 79948 115906 79960
rect 210510 79948 210516 79960
rect 115900 79920 210516 79948
rect 115900 79908 115906 79920
rect 210510 79908 210516 79920
rect 210568 79908 210574 79960
rect 122742 79840 122748 79892
rect 122800 79880 122806 79892
rect 213178 79880 213184 79892
rect 122800 79852 213184 79880
rect 122800 79840 122806 79852
rect 213178 79840 213184 79852
rect 213236 79840 213242 79892
rect 89622 79772 89628 79824
rect 89680 79812 89686 79824
rect 167822 79812 167828 79824
rect 89680 79784 167828 79812
rect 89680 79772 89686 79784
rect 167822 79772 167828 79784
rect 167880 79772 167886 79824
rect 276658 79296 276664 79348
rect 276716 79336 276722 79348
rect 310422 79336 310428 79348
rect 276716 79308 310428 79336
rect 276716 79296 276722 79308
rect 310422 79296 310428 79308
rect 310480 79296 310486 79348
rect 99282 78616 99288 78668
rect 99340 78656 99346 78668
rect 186958 78656 186964 78668
rect 99340 78628 186964 78656
rect 99340 78616 99346 78628
rect 186958 78616 186964 78628
rect 187016 78616 187022 78668
rect 245654 78616 245660 78668
rect 245712 78656 245718 78668
rect 411254 78656 411260 78668
rect 245712 78628 411260 78656
rect 245712 78616 245718 78628
rect 411254 78616 411260 78628
rect 411312 78616 411318 78668
rect 86862 78548 86868 78600
rect 86920 78588 86926 78600
rect 172054 78588 172060 78600
rect 86920 78560 172060 78588
rect 86920 78548 86926 78560
rect 172054 78548 172060 78560
rect 172112 78548 172118 78600
rect 124122 78480 124128 78532
rect 124180 78520 124186 78532
rect 206370 78520 206376 78532
rect 124180 78492 206376 78520
rect 124180 78480 124186 78492
rect 206370 78480 206376 78492
rect 206428 78480 206434 78532
rect 134518 78412 134524 78464
rect 134576 78452 134582 78464
rect 192662 78452 192668 78464
rect 134576 78424 192668 78452
rect 134576 78412 134582 78424
rect 192662 78412 192668 78424
rect 192720 78412 192726 78464
rect 334710 77256 334716 77308
rect 334768 77296 334774 77308
rect 336826 77296 336832 77308
rect 334768 77268 336832 77296
rect 334768 77256 334774 77268
rect 336826 77256 336832 77268
rect 336884 77256 336890 77308
rect 116578 77188 116584 77240
rect 116636 77228 116642 77240
rect 214742 77228 214748 77240
rect 116636 77200 214748 77228
rect 116636 77188 116642 77200
rect 214742 77188 214748 77200
rect 214800 77188 214806 77240
rect 285582 77188 285588 77240
rect 285640 77228 285646 77240
rect 286870 77228 286876 77240
rect 285640 77200 286876 77228
rect 285640 77188 285646 77200
rect 286870 77188 286876 77200
rect 286928 77228 286934 77240
rect 433334 77228 433340 77240
rect 286928 77200 433340 77228
rect 286928 77188 286934 77200
rect 433334 77188 433340 77200
rect 433392 77188 433398 77240
rect 113082 77120 113088 77172
rect 113140 77160 113146 77172
rect 202230 77160 202236 77172
rect 113140 77132 202236 77160
rect 113140 77120 113146 77132
rect 202230 77120 202236 77132
rect 202288 77120 202294 77172
rect 75914 76576 75920 76628
rect 75972 76616 75978 76628
rect 285122 76616 285128 76628
rect 75972 76588 285128 76616
rect 75972 76576 75978 76588
rect 285122 76576 285128 76588
rect 285180 76576 285186 76628
rect 63494 76508 63500 76560
rect 63552 76548 63558 76560
rect 303062 76548 303068 76560
rect 63552 76520 303068 76548
rect 63552 76508 63558 76520
rect 303062 76508 303068 76520
rect 303120 76508 303126 76560
rect 85482 75828 85488 75880
rect 85540 75868 85546 75880
rect 196710 75868 196716 75880
rect 85540 75840 196716 75868
rect 85540 75828 85546 75840
rect 196710 75828 196716 75840
rect 196768 75828 196774 75880
rect 119338 75760 119344 75812
rect 119396 75800 119402 75812
rect 203702 75800 203708 75812
rect 119396 75772 203708 75800
rect 119396 75760 119402 75772
rect 203702 75760 203708 75772
rect 203760 75760 203766 75812
rect 139394 75216 139400 75268
rect 139452 75256 139458 75268
rect 323578 75256 323584 75268
rect 139452 75228 323584 75256
rect 139452 75216 139458 75228
rect 323578 75216 323584 75228
rect 323636 75216 323642 75268
rect 23474 75148 23480 75200
rect 23532 75188 23538 75200
rect 297542 75188 297548 75200
rect 23532 75160 297548 75188
rect 23532 75148 23538 75160
rect 297542 75148 297548 75160
rect 297600 75148 297606 75200
rect 67634 74468 67640 74520
rect 67692 74508 67698 74520
rect 195330 74508 195336 74520
rect 67692 74480 195336 74508
rect 67692 74468 67698 74480
rect 195330 74468 195336 74480
rect 195388 74468 195394 74520
rect 177758 73924 177764 73976
rect 177816 73964 177822 73976
rect 347038 73964 347044 73976
rect 177816 73936 347044 73964
rect 177816 73924 177822 73936
rect 347038 73924 347044 73936
rect 347096 73924 347102 73976
rect 35894 73856 35900 73908
rect 35952 73896 35958 73908
rect 268470 73896 268476 73908
rect 35952 73868 268476 73896
rect 35952 73856 35958 73868
rect 268470 73856 268476 73868
rect 268528 73856 268534 73908
rect 20714 73788 20720 73840
rect 20772 73828 20778 73840
rect 297358 73828 297364 73840
rect 20772 73800 297364 73828
rect 20772 73788 20778 73800
rect 297358 73788 297364 73800
rect 297416 73788 297422 73840
rect 346394 73788 346400 73840
rect 346452 73828 346458 73840
rect 451550 73828 451556 73840
rect 346452 73800 451556 73828
rect 346452 73788 346458 73800
rect 451550 73788 451556 73800
rect 451608 73788 451614 73840
rect 104802 73108 104808 73160
rect 104860 73148 104866 73160
rect 198090 73148 198096 73160
rect 104860 73120 198096 73148
rect 104860 73108 104866 73120
rect 198090 73108 198096 73120
rect 198148 73108 198154 73160
rect 438854 73108 438860 73160
rect 438912 73148 438918 73160
rect 471974 73148 471980 73160
rect 438912 73120 471980 73148
rect 438912 73108 438918 73120
rect 471974 73108 471980 73120
rect 472032 73148 472038 73160
rect 580166 73148 580172 73160
rect 472032 73120 580172 73148
rect 472032 73108 472038 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 124214 72496 124220 72548
rect 124272 72536 124278 72548
rect 250530 72536 250536 72548
rect 124272 72508 250536 72536
rect 124272 72496 124278 72508
rect 250530 72496 250536 72508
rect 250588 72496 250594 72548
rect 247678 72428 247684 72480
rect 247736 72468 247742 72480
rect 418890 72468 418896 72480
rect 247736 72440 418896 72468
rect 247736 72428 247742 72440
rect 418890 72428 418896 72440
rect 418948 72428 418954 72480
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 44818 71720 44824 71732
rect 3476 71692 44824 71720
rect 3476 71680 3482 71692
rect 44818 71680 44824 71692
rect 44876 71680 44882 71732
rect 88334 71068 88340 71120
rect 88392 71108 88398 71120
rect 300210 71108 300216 71120
rect 88392 71080 300216 71108
rect 88392 71068 88398 71080
rect 300210 71068 300216 71080
rect 300268 71068 300274 71120
rect 303614 71068 303620 71120
rect 303672 71108 303678 71120
rect 396810 71108 396816 71120
rect 303672 71080 396816 71108
rect 303672 71068 303678 71080
rect 396810 71068 396816 71080
rect 396868 71068 396874 71120
rect 69014 71000 69020 71052
rect 69072 71040 69078 71052
rect 304626 71040 304632 71052
rect 69072 71012 304632 71040
rect 69072 71000 69078 71012
rect 304626 71000 304632 71012
rect 304684 71000 304690 71052
rect 271138 69776 271144 69828
rect 271196 69816 271202 69828
rect 451734 69816 451740 69828
rect 271196 69788 451740 69816
rect 271196 69776 271202 69788
rect 451734 69776 451740 69788
rect 451792 69776 451798 69828
rect 74534 69708 74540 69760
rect 74592 69748 74598 69760
rect 282454 69748 282460 69760
rect 74592 69720 282460 69748
rect 74592 69708 74598 69720
rect 282454 69708 282460 69720
rect 282512 69708 282518 69760
rect 64874 69640 64880 69692
rect 64932 69680 64938 69692
rect 305914 69680 305920 69692
rect 64932 69652 305920 69680
rect 64932 69640 64938 69652
rect 305914 69640 305920 69652
rect 305972 69640 305978 69692
rect 89714 68280 89720 68332
rect 89772 68320 89778 68332
rect 249150 68320 249156 68332
rect 89772 68292 249156 68320
rect 89772 68280 89778 68292
rect 249150 68280 249156 68292
rect 249208 68280 249214 68332
rect 184934 66988 184940 67040
rect 184992 67028 184998 67040
rect 315298 67028 315304 67040
rect 184992 67000 315304 67028
rect 184992 66988 184998 67000
rect 315298 66988 315304 67000
rect 315356 66988 315362 67040
rect 100754 66920 100760 66972
rect 100812 66960 100818 66972
rect 275370 66960 275376 66972
rect 100812 66932 275376 66960
rect 100812 66920 100818 66932
rect 275370 66920 275376 66932
rect 275428 66920 275434 66972
rect 62114 66852 62120 66904
rect 62172 66892 62178 66904
rect 304442 66892 304448 66904
rect 62172 66864 304448 66892
rect 62172 66852 62178 66864
rect 304442 66852 304448 66864
rect 304500 66852 304506 66904
rect 324958 66852 324964 66904
rect 325016 66892 325022 66904
rect 451366 66892 451372 66904
rect 325016 66864 451372 66892
rect 325016 66852 325022 66864
rect 451366 66852 451372 66864
rect 451424 66852 451430 66904
rect 110414 65560 110420 65612
rect 110472 65600 110478 65612
rect 263042 65600 263048 65612
rect 110472 65572 263048 65600
rect 110472 65560 110478 65572
rect 263042 65560 263048 65572
rect 263100 65560 263106 65612
rect 80054 65492 80060 65544
rect 80112 65532 80118 65544
rect 279510 65532 279516 65544
rect 80112 65504 279516 65532
rect 80112 65492 80118 65504
rect 279510 65492 279516 65504
rect 279568 65492 279574 65544
rect 284202 64812 284208 64864
rect 284260 64852 284266 64864
rect 447778 64852 447784 64864
rect 284260 64824 447784 64852
rect 284260 64812 284266 64824
rect 447778 64812 447784 64824
rect 447836 64812 447842 64864
rect 241514 64268 241520 64320
rect 241572 64308 241578 64320
rect 284202 64308 284208 64320
rect 241572 64280 284208 64308
rect 241572 64268 241578 64280
rect 284202 64268 284208 64280
rect 284260 64268 284266 64320
rect 38654 64200 38660 64252
rect 38712 64240 38718 64252
rect 285030 64240 285036 64252
rect 38712 64212 285036 64240
rect 38712 64200 38718 64212
rect 285030 64200 285036 64212
rect 285088 64200 285094 64252
rect 33134 64132 33140 64184
rect 33192 64172 33198 64184
rect 301774 64172 301780 64184
rect 33192 64144 301780 64172
rect 33192 64132 33198 64144
rect 301774 64132 301780 64144
rect 301832 64132 301838 64184
rect 70394 62840 70400 62892
rect 70452 62880 70458 62892
rect 269850 62880 269856 62892
rect 70452 62852 269856 62880
rect 70452 62840 70458 62852
rect 269850 62840 269856 62852
rect 269908 62840 269914 62892
rect 53834 62772 53840 62824
rect 53892 62812 53898 62824
rect 293402 62812 293408 62824
rect 53892 62784 293408 62812
rect 53892 62772 53898 62784
rect 293402 62772 293408 62784
rect 293460 62772 293466 62824
rect 197998 61480 198004 61532
rect 198056 61520 198062 61532
rect 273254 61520 273260 61532
rect 198056 61492 273260 61520
rect 198056 61480 198062 61492
rect 273254 61480 273260 61492
rect 273312 61520 273318 61532
rect 354030 61520 354036 61532
rect 273312 61492 354036 61520
rect 273312 61480 273318 61492
rect 354030 61480 354036 61492
rect 354088 61480 354094 61532
rect 95234 61412 95240 61464
rect 95292 61452 95298 61464
rect 280798 61452 280804 61464
rect 95292 61424 280804 61452
rect 95292 61412 95298 61424
rect 280798 61412 280804 61424
rect 280856 61412 280862 61464
rect 71774 61344 71780 61396
rect 71832 61384 71838 61396
rect 274082 61384 274088 61396
rect 71832 61356 274088 61384
rect 71832 61344 71838 61356
rect 274082 61344 274088 61356
rect 274140 61344 274146 61396
rect 345014 61344 345020 61396
rect 345072 61384 345078 61396
rect 408494 61384 408500 61396
rect 345072 61356 408500 61384
rect 345072 61344 345078 61356
rect 408494 61344 408500 61356
rect 408552 61344 408558 61396
rect 460198 60664 460204 60716
rect 460256 60704 460262 60716
rect 580166 60704 580172 60716
rect 460256 60676 580172 60704
rect 460256 60664 460262 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 99374 60052 99380 60104
rect 99432 60092 99438 60104
rect 266998 60092 267004 60104
rect 99432 60064 267004 60092
rect 99432 60052 99438 60064
rect 266998 60052 267004 60064
rect 267056 60052 267062 60104
rect 269114 60052 269120 60104
rect 269172 60092 269178 60104
rect 363598 60092 363604 60104
rect 269172 60064 363604 60092
rect 269172 60052 269178 60064
rect 363598 60052 363604 60064
rect 363656 60052 363662 60104
rect 11054 59984 11060 60036
rect 11112 60024 11118 60036
rect 303154 60024 303160 60036
rect 11112 59996 303160 60024
rect 11112 59984 11118 59996
rect 303154 59984 303160 59996
rect 303212 59984 303218 60036
rect 355318 59984 355324 60036
rect 355376 60024 355382 60036
rect 416774 60024 416780 60036
rect 355376 59996 416780 60024
rect 355376 59984 355382 59996
rect 416774 59984 416780 59996
rect 416832 59984 416838 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 62758 59344 62764 59356
rect 3108 59316 62764 59344
rect 3108 59304 3114 59316
rect 62758 59304 62764 59316
rect 62816 59304 62822 59356
rect 350534 59304 350540 59356
rect 350592 59344 350598 59356
rect 434714 59344 434720 59356
rect 350592 59316 434720 59344
rect 350592 59304 350598 59316
rect 434714 59304 434720 59316
rect 434772 59304 434778 59356
rect 266446 58760 266452 58812
rect 266504 58800 266510 58812
rect 350534 58800 350540 58812
rect 266504 58772 350540 58800
rect 266504 58760 266510 58772
rect 350534 58760 350540 58772
rect 350592 58760 350598 58812
rect 106274 58692 106280 58744
rect 106332 58732 106338 58744
rect 276750 58732 276756 58744
rect 106332 58704 276756 58732
rect 106332 58692 106338 58704
rect 276750 58692 276756 58704
rect 276808 58692 276814 58744
rect 85574 58624 85580 58676
rect 85632 58664 85638 58676
rect 296162 58664 296168 58676
rect 85632 58636 296168 58664
rect 85632 58624 85638 58636
rect 296162 58624 296168 58636
rect 296220 58624 296226 58676
rect 341518 57944 341524 57996
rect 341576 57984 341582 57996
rect 345014 57984 345020 57996
rect 341576 57956 345020 57984
rect 341576 57944 341582 57956
rect 345014 57944 345020 57956
rect 345072 57944 345078 57996
rect 103514 57264 103520 57316
rect 103572 57304 103578 57316
rect 300394 57304 300400 57316
rect 103572 57276 300400 57304
rect 103572 57264 103578 57276
rect 300394 57264 300400 57276
rect 300452 57264 300458 57316
rect 13814 57196 13820 57248
rect 13872 57236 13878 57248
rect 284938 57236 284944 57248
rect 13872 57208 284944 57236
rect 13872 57196 13878 57208
rect 284938 57196 284944 57208
rect 284996 57196 285002 57248
rect 296162 57196 296168 57248
rect 296220 57236 296226 57248
rect 435358 57236 435364 57248
rect 296220 57208 435364 57236
rect 296220 57196 296226 57208
rect 435358 57196 435364 57208
rect 435416 57196 435422 57248
rect 255314 55972 255320 56024
rect 255372 56012 255378 56024
rect 269758 56012 269764 56024
rect 255372 55984 269764 56012
rect 255372 55972 255378 55984
rect 269758 55972 269764 55984
rect 269816 55972 269822 56024
rect 110506 55904 110512 55956
rect 110564 55944 110570 55956
rect 293310 55944 293316 55956
rect 110564 55916 293316 55944
rect 110564 55904 110570 55916
rect 293310 55904 293316 55916
rect 293368 55904 293374 55956
rect 19334 55836 19340 55888
rect 19392 55876 19398 55888
rect 260190 55876 260196 55888
rect 19392 55848 260196 55876
rect 19392 55836 19398 55848
rect 260190 55836 260196 55848
rect 260248 55836 260254 55888
rect 4062 55156 4068 55208
rect 4120 55196 4126 55208
rect 251174 55196 251180 55208
rect 4120 55168 251180 55196
rect 4120 55156 4126 55168
rect 251174 55156 251180 55168
rect 251232 55156 251238 55208
rect 262122 54544 262128 54596
rect 262180 54584 262186 54596
rect 381538 54584 381544 54596
rect 262180 54556 381544 54584
rect 262180 54544 262186 54556
rect 381538 54544 381544 54556
rect 381596 54544 381602 54596
rect 56594 54476 56600 54528
rect 56652 54516 56658 54528
rect 264422 54516 264428 54528
rect 56652 54488 264428 54516
rect 56652 54476 56658 54488
rect 264422 54476 264428 54488
rect 264480 54476 264486 54528
rect 3418 53796 3424 53848
rect 3476 53836 3482 53848
rect 4062 53836 4068 53848
rect 3476 53808 4068 53836
rect 3476 53796 3482 53808
rect 4062 53796 4068 53808
rect 4120 53796 4126 53848
rect 281442 53728 281448 53780
rect 281500 53768 281506 53780
rect 395430 53768 395436 53780
rect 281500 53740 395436 53768
rect 281500 53728 281506 53740
rect 395430 53728 395436 53740
rect 395488 53728 395494 53780
rect 73154 53116 73160 53168
rect 73212 53156 73218 53168
rect 292114 53156 292120 53168
rect 73212 53128 292120 53156
rect 73212 53116 73218 53128
rect 292114 53116 292120 53128
rect 292172 53116 292178 53168
rect 19426 53048 19432 53100
rect 19484 53088 19490 53100
rect 283650 53088 283656 53100
rect 19484 53060 283656 53088
rect 19484 53048 19490 53060
rect 283650 53048 283656 53060
rect 283708 53048 283714 53100
rect 280154 52436 280160 52488
rect 280212 52476 280218 52488
rect 281442 52476 281448 52488
rect 280212 52448 281448 52476
rect 280212 52436 280218 52448
rect 281442 52436 281448 52448
rect 281500 52436 281506 52488
rect 244918 51824 244924 51876
rect 244976 51864 244982 51876
rect 409138 51864 409144 51876
rect 244976 51836 409144 51864
rect 244976 51824 244982 51836
rect 409138 51824 409144 51836
rect 409196 51824 409202 51876
rect 45554 51756 45560 51808
rect 45612 51796 45618 51808
rect 273990 51796 273996 51808
rect 45612 51768 273996 51796
rect 45612 51756 45618 51768
rect 273990 51756 273996 51768
rect 274048 51756 274054 51808
rect 28994 51688 29000 51740
rect 29052 51728 29058 51740
rect 296254 51728 296260 51740
rect 29052 51700 296260 51728
rect 29052 51688 29058 51700
rect 296254 51688 296260 51700
rect 296312 51688 296318 51740
rect 51074 50396 51080 50448
rect 51132 50436 51138 50448
rect 262950 50436 262956 50448
rect 51132 50408 262956 50436
rect 51132 50396 51138 50408
rect 262950 50396 262956 50408
rect 263008 50396 263014 50448
rect 284938 50396 284944 50448
rect 284996 50436 285002 50448
rect 342990 50436 342996 50448
rect 284996 50408 342996 50436
rect 284996 50396 285002 50408
rect 342990 50396 342996 50408
rect 343048 50396 343054 50448
rect 67634 50328 67640 50380
rect 67692 50368 67698 50380
rect 297450 50368 297456 50380
rect 67692 50340 297456 50368
rect 67692 50328 67698 50340
rect 297450 50328 297456 50340
rect 297508 50328 297514 50380
rect 342346 50328 342352 50380
rect 342404 50368 342410 50380
rect 405734 50368 405740 50380
rect 342404 50340 405740 50368
rect 342404 50328 342410 50340
rect 405734 50328 405740 50340
rect 405792 50328 405798 50380
rect 77294 49036 77300 49088
rect 77352 49076 77358 49088
rect 296070 49076 296076 49088
rect 77352 49048 296076 49076
rect 77352 49036 77358 49048
rect 296070 49036 296076 49048
rect 296128 49036 296134 49088
rect 2774 48968 2780 49020
rect 2832 49008 2838 49020
rect 286318 49008 286324 49020
rect 2832 48980 286324 49008
rect 2832 48968 2838 48980
rect 286318 48968 286324 48980
rect 286376 48968 286382 49020
rect 298094 48968 298100 49020
rect 298152 49008 298158 49020
rect 337470 49008 337476 49020
rect 298152 48980 337476 49008
rect 298152 48968 298158 48980
rect 337470 48968 337476 48980
rect 337528 48968 337534 49020
rect 342898 48968 342904 49020
rect 342956 49008 342962 49020
rect 444374 49008 444380 49020
rect 342956 48980 444380 49008
rect 342956 48968 342962 48980
rect 444374 48968 444380 48980
rect 444432 48968 444438 49020
rect 291838 48288 291844 48340
rect 291896 48328 291902 48340
rect 298094 48328 298100 48340
rect 291896 48300 298100 48328
rect 291896 48288 291902 48300
rect 298094 48288 298100 48300
rect 298152 48288 298158 48340
rect 216030 47676 216036 47728
rect 216088 47716 216094 47728
rect 292574 47716 292580 47728
rect 216088 47688 292580 47716
rect 216088 47676 216094 47688
rect 292574 47676 292580 47688
rect 292632 47716 292638 47728
rect 373350 47716 373356 47728
rect 292632 47688 373356 47716
rect 292632 47676 292638 47688
rect 373350 47676 373356 47688
rect 373408 47676 373414 47728
rect 92474 47608 92480 47660
rect 92532 47648 92538 47660
rect 298738 47648 298744 47660
rect 92532 47620 298744 47648
rect 92532 47608 92538 47620
rect 298738 47608 298744 47620
rect 298796 47608 298802 47660
rect 60734 47540 60740 47592
rect 60792 47580 60798 47592
rect 294782 47580 294788 47592
rect 60792 47552 294788 47580
rect 60792 47540 60798 47552
rect 294782 47540 294788 47552
rect 294840 47540 294846 47592
rect 271690 46860 271696 46912
rect 271748 46900 271754 46912
rect 398098 46900 398104 46912
rect 271748 46872 398104 46900
rect 271748 46860 271754 46872
rect 398098 46860 398104 46872
rect 398156 46860 398162 46912
rect 399570 46860 399576 46912
rect 399628 46900 399634 46912
rect 580166 46900 580172 46912
rect 399628 46872 580172 46900
rect 399628 46860 399634 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 26234 46248 26240 46300
rect 26292 46288 26298 46300
rect 257522 46288 257528 46300
rect 26292 46260 257528 46288
rect 26292 46248 26298 46260
rect 257522 46248 257528 46260
rect 257580 46248 257586 46300
rect 42794 46180 42800 46232
rect 42852 46220 42858 46232
rect 292022 46220 292028 46232
rect 42852 46192 292028 46220
rect 42852 46180 42858 46192
rect 292022 46180 292028 46192
rect 292080 46180 292086 46232
rect 248414 45568 248420 45620
rect 248472 45608 248478 45620
rect 271690 45608 271696 45620
rect 248472 45580 271696 45608
rect 248472 45568 248478 45580
rect 271690 45568 271696 45580
rect 271748 45568 271754 45620
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 48958 45540 48964 45552
rect 3568 45512 48964 45540
rect 3568 45500 3574 45512
rect 48958 45500 48964 45512
rect 49016 45500 49022 45552
rect 59354 44888 59360 44940
rect 59412 44928 59418 44940
rect 298830 44928 298836 44940
rect 59412 44900 298836 44928
rect 59412 44888 59418 44900
rect 298830 44888 298836 44900
rect 298888 44888 298894 44940
rect 44174 44820 44180 44872
rect 44232 44860 44238 44872
rect 287974 44860 287980 44872
rect 44232 44832 287980 44860
rect 44232 44820 44238 44832
rect 287974 44820 287980 44832
rect 288032 44820 288038 44872
rect 81434 43460 81440 43512
rect 81492 43500 81498 43512
rect 289262 43500 289268 43512
rect 81492 43472 289268 43500
rect 81492 43460 81498 43472
rect 289262 43460 289268 43472
rect 289320 43460 289326 43512
rect 295334 43460 295340 43512
rect 295392 43500 295398 43512
rect 329282 43500 329288 43512
rect 295392 43472 329288 43500
rect 295392 43460 295398 43472
rect 329282 43460 329288 43472
rect 329340 43460 329346 43512
rect 6914 43392 6920 43444
rect 6972 43432 6978 43444
rect 300302 43432 300308 43444
rect 6972 43404 300308 43432
rect 6972 43392 6978 43404
rect 300302 43392 300308 43404
rect 300360 43392 300366 43444
rect 177850 42168 177856 42220
rect 177908 42208 177914 42220
rect 337470 42208 337476 42220
rect 177908 42180 337476 42208
rect 177908 42168 177914 42180
rect 337470 42168 337476 42180
rect 337528 42168 337534 42220
rect 118694 42100 118700 42152
rect 118752 42140 118758 42152
rect 301590 42140 301596 42152
rect 118752 42112 301596 42140
rect 118752 42100 118758 42112
rect 301590 42100 301596 42112
rect 301648 42100 301654 42152
rect 44266 42032 44272 42084
rect 44324 42072 44330 42084
rect 262858 42072 262864 42084
rect 44324 42044 262864 42072
rect 44324 42032 44330 42044
rect 262858 42032 262864 42044
rect 262916 42032 262922 42084
rect 342254 41352 342260 41404
rect 342312 41392 342318 41404
rect 422938 41392 422944 41404
rect 342312 41364 422944 41392
rect 342312 41352 342318 41364
rect 422938 41352 422944 41364
rect 422996 41352 423002 41404
rect 338022 41284 338028 41336
rect 338080 41324 338086 41336
rect 359458 41324 359464 41336
rect 338080 41296 359464 41324
rect 338080 41284 338086 41296
rect 359458 41284 359464 41296
rect 359516 41284 359522 41336
rect 85666 40740 85672 40792
rect 85724 40780 85730 40792
rect 290458 40780 290464 40792
rect 85724 40752 290464 40780
rect 85724 40740 85730 40752
rect 290458 40740 290464 40752
rect 290516 40740 290522 40792
rect 322934 40740 322940 40792
rect 322992 40780 322998 40792
rect 342254 40780 342260 40792
rect 322992 40752 342260 40780
rect 322992 40740 322998 40752
rect 342254 40740 342260 40752
rect 342312 40740 342318 40792
rect 46934 40672 46940 40724
rect 46992 40712 46998 40724
rect 257430 40712 257436 40724
rect 46992 40684 257436 40712
rect 46992 40672 46998 40684
rect 257430 40672 257436 40684
rect 257488 40672 257494 40724
rect 259454 40672 259460 40724
rect 259512 40712 259518 40724
rect 336734 40712 336740 40724
rect 259512 40684 336740 40712
rect 259512 40672 259518 40684
rect 336734 40672 336740 40684
rect 336792 40712 336798 40724
rect 338022 40712 338028 40724
rect 336792 40684 338028 40712
rect 336792 40672 336798 40684
rect 338022 40672 338028 40684
rect 338080 40672 338086 40724
rect 121454 39448 121460 39500
rect 121512 39488 121518 39500
rect 271230 39488 271236 39500
rect 121512 39460 271236 39488
rect 121512 39448 121518 39460
rect 271230 39448 271236 39460
rect 271288 39448 271294 39500
rect 256050 39380 256056 39432
rect 256108 39420 256114 39432
rect 445846 39420 445852 39432
rect 256108 39392 445852 39420
rect 256108 39380 256114 39392
rect 445846 39380 445852 39392
rect 445904 39380 445910 39432
rect 37274 39312 37280 39364
rect 37332 39352 37338 39364
rect 307110 39352 307116 39364
rect 37332 39324 307116 39352
rect 37332 39312 37338 39324
rect 307110 39312 307116 39324
rect 307168 39312 307174 39364
rect 209682 38564 209688 38616
rect 209740 38604 209746 38616
rect 324314 38604 324320 38616
rect 209740 38576 324320 38604
rect 209740 38564 209746 38576
rect 324314 38564 324320 38576
rect 324372 38604 324378 38616
rect 324958 38604 324964 38616
rect 324372 38576 324964 38604
rect 324372 38564 324378 38576
rect 324958 38564 324964 38576
rect 325016 38564 325022 38616
rect 364978 38564 364984 38616
rect 365036 38604 365042 38616
rect 365622 38604 365628 38616
rect 365036 38576 365628 38604
rect 365036 38564 365042 38576
rect 365622 38564 365628 38576
rect 365680 38604 365686 38616
rect 451274 38604 451280 38616
rect 365680 38576 451280 38604
rect 365680 38564 365686 38576
rect 451274 38564 451280 38576
rect 451332 38564 451338 38616
rect 128354 37952 128360 38004
rect 128412 37992 128418 38004
rect 216674 37992 216680 38004
rect 128412 37964 216680 37992
rect 128412 37952 128418 37964
rect 216674 37952 216680 37964
rect 216732 37952 216738 38004
rect 251174 37952 251180 38004
rect 251232 37992 251238 38004
rect 365070 37992 365076 38004
rect 251232 37964 365076 37992
rect 251232 37952 251238 37964
rect 365070 37952 365076 37964
rect 365128 37952 365134 38004
rect 27614 37884 27620 37936
rect 27672 37924 27678 37936
rect 279418 37924 279424 37936
rect 27672 37896 279424 37924
rect 27672 37884 27678 37896
rect 279418 37884 279424 37896
rect 279476 37884 279482 37936
rect 329834 37884 329840 37936
rect 329892 37924 329898 37936
rect 365622 37924 365628 37936
rect 329892 37896 365628 37924
rect 329892 37884 329898 37896
rect 365622 37884 365628 37896
rect 365680 37884 365686 37936
rect 240778 36660 240784 36712
rect 240836 36700 240842 36712
rect 407206 36700 407212 36712
rect 240836 36672 407212 36700
rect 240836 36660 240842 36672
rect 407206 36660 407212 36672
rect 407264 36660 407270 36712
rect 11146 36592 11152 36644
rect 11204 36632 11210 36644
rect 255958 36632 255964 36644
rect 11204 36604 255964 36632
rect 11204 36592 11210 36604
rect 255958 36592 255964 36604
rect 256016 36592 256022 36644
rect 35986 36524 35992 36576
rect 36044 36564 36050 36576
rect 305822 36564 305828 36576
rect 36044 36536 305828 36564
rect 36044 36524 36050 36536
rect 305822 36524 305828 36536
rect 305880 36524 305886 36576
rect 179414 35300 179420 35352
rect 179472 35340 179478 35352
rect 254670 35340 254676 35352
rect 179472 35312 254676 35340
rect 179472 35300 179478 35312
rect 254670 35300 254676 35312
rect 254728 35300 254734 35352
rect 207014 35232 207020 35284
rect 207072 35272 207078 35284
rect 345750 35272 345756 35284
rect 207072 35244 345756 35272
rect 207072 35232 207078 35244
rect 345750 35232 345756 35244
rect 345808 35232 345814 35284
rect 48314 35164 48320 35216
rect 48372 35204 48378 35216
rect 272518 35204 272524 35216
rect 48372 35176 272524 35204
rect 48372 35164 48378 35176
rect 272518 35164 272524 35176
rect 272576 35164 272582 35216
rect 292022 35164 292028 35216
rect 292080 35204 292086 35216
rect 398834 35204 398840 35216
rect 292080 35176 398840 35204
rect 292080 35164 292086 35176
rect 398834 35164 398840 35176
rect 398892 35164 398898 35216
rect 427722 35164 427728 35216
rect 427780 35204 427786 35216
rect 464614 35204 464620 35216
rect 427780 35176 464620 35204
rect 427780 35164 427786 35176
rect 464614 35164 464620 35176
rect 464672 35164 464678 35216
rect 254670 34484 254676 34536
rect 254728 34524 254734 34536
rect 256050 34524 256056 34536
rect 254728 34496 256056 34524
rect 254728 34484 254734 34496
rect 256050 34484 256056 34496
rect 256108 34484 256114 34536
rect 143534 33872 143540 33924
rect 143592 33912 143598 33924
rect 331950 33912 331956 33924
rect 143592 33884 331956 33912
rect 143592 33872 143598 33884
rect 331950 33872 331956 33884
rect 332008 33872 332014 33924
rect 30374 33804 30380 33856
rect 30432 33844 30438 33856
rect 265618 33844 265624 33856
rect 30432 33816 265624 33844
rect 30432 33804 30438 33816
rect 265618 33804 265624 33816
rect 265676 33804 265682 33856
rect 52454 33736 52460 33788
rect 52512 33776 52518 33788
rect 304350 33776 304356 33788
rect 52512 33748 304356 33776
rect 52512 33736 52518 33748
rect 304350 33736 304356 33748
rect 304408 33736 304414 33788
rect 349798 33736 349804 33788
rect 349856 33776 349862 33788
rect 438118 33776 438124 33788
rect 349856 33748 438124 33776
rect 349856 33736 349862 33748
rect 438118 33736 438124 33748
rect 438176 33736 438182 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 35158 33096 35164 33108
rect 3568 33068 35164 33096
rect 3568 33056 3574 33068
rect 35158 33056 35164 33068
rect 35216 33056 35222 33108
rect 337470 33056 337476 33108
rect 337528 33096 337534 33108
rect 449986 33096 449992 33108
rect 337528 33068 449992 33096
rect 337528 33056 337534 33068
rect 449986 33056 449992 33068
rect 450044 33056 450050 33108
rect 464614 33056 464620 33108
rect 464672 33096 464678 33108
rect 579890 33096 579896 33108
rect 464672 33068 579896 33096
rect 464672 33056 464678 33068
rect 579890 33056 579896 33068
rect 579948 33056 579954 33108
rect 91094 32376 91100 32428
rect 91152 32416 91158 32428
rect 264330 32416 264336 32428
rect 91152 32388 264336 32416
rect 91152 32376 91158 32388
rect 264330 32376 264336 32388
rect 264388 32376 264394 32428
rect 309870 32376 309876 32428
rect 309928 32416 309934 32428
rect 324958 32416 324964 32428
rect 309928 32388 324964 32416
rect 309928 32376 309934 32388
rect 324958 32376 324964 32388
rect 325016 32376 325022 32428
rect 336734 31764 336740 31816
rect 336792 31804 336798 31816
rect 337470 31804 337476 31816
rect 336792 31776 337476 31804
rect 336792 31764 336798 31776
rect 337470 31764 337476 31776
rect 337528 31764 337534 31816
rect 320818 31696 320824 31748
rect 320876 31736 320882 31748
rect 396902 31736 396908 31748
rect 320876 31708 396908 31736
rect 320876 31696 320882 31708
rect 396902 31696 396908 31708
rect 396960 31696 396966 31748
rect 320174 31220 320180 31272
rect 320232 31260 320238 31272
rect 320818 31260 320824 31272
rect 320232 31232 320824 31260
rect 320232 31220 320238 31232
rect 320818 31220 320824 31232
rect 320876 31220 320882 31272
rect 201494 31152 201500 31204
rect 201552 31192 201558 31204
rect 335998 31192 336004 31204
rect 201552 31164 336004 31192
rect 201552 31152 201558 31164
rect 335998 31152 336004 31164
rect 336056 31152 336062 31204
rect 66254 31084 66260 31136
rect 66312 31124 66318 31136
rect 302970 31124 302976 31136
rect 66312 31096 302976 31124
rect 66312 31084 66318 31096
rect 302970 31084 302976 31096
rect 303028 31084 303034 31136
rect 5534 31016 5540 31068
rect 5592 31056 5598 31068
rect 251910 31056 251916 31068
rect 5592 31028 251916 31056
rect 5592 31016 5598 31028
rect 251910 31016 251916 31028
rect 251968 31016 251974 31068
rect 97994 29588 98000 29640
rect 98052 29628 98058 29640
rect 260098 29628 260104 29640
rect 98052 29600 260104 29628
rect 98052 29588 98058 29600
rect 260098 29588 260104 29600
rect 260156 29588 260162 29640
rect 317506 28908 317512 28960
rect 317564 28948 317570 28960
rect 318702 28948 318708 28960
rect 317564 28920 318708 28948
rect 317564 28908 317570 28920
rect 318702 28908 318708 28920
rect 318760 28948 318766 28960
rect 391290 28948 391296 28960
rect 318760 28920 391296 28948
rect 318760 28908 318766 28920
rect 391290 28908 391296 28920
rect 391348 28908 391354 28960
rect 86954 28296 86960 28348
rect 87012 28336 87018 28348
rect 287790 28336 287796 28348
rect 87012 28308 287796 28336
rect 87012 28296 87018 28308
rect 287790 28296 287796 28308
rect 287848 28296 287854 28348
rect 93854 28228 93860 28280
rect 93912 28268 93918 28280
rect 305638 28268 305644 28280
rect 93912 28240 305644 28268
rect 93912 28228 93918 28240
rect 305638 28228 305644 28240
rect 305696 28228 305702 28280
rect 309134 27616 309140 27668
rect 309192 27656 309198 27668
rect 318702 27656 318708 27668
rect 309192 27628 318708 27656
rect 309192 27616 309198 27628
rect 318702 27616 318708 27628
rect 318760 27616 318766 27668
rect 200114 27548 200120 27600
rect 200172 27588 200178 27600
rect 311894 27588 311900 27600
rect 200172 27560 311900 27588
rect 200172 27548 200178 27560
rect 311894 27548 311900 27560
rect 311952 27588 311958 27600
rect 312538 27588 312544 27600
rect 311952 27560 312544 27588
rect 311952 27548 311958 27560
rect 312538 27548 312544 27560
rect 312596 27548 312602 27600
rect 117314 26936 117320 26988
rect 117372 26976 117378 26988
rect 282270 26976 282276 26988
rect 117372 26948 282276 26976
rect 117372 26936 117378 26948
rect 282270 26936 282276 26948
rect 282328 26936 282334 26988
rect 78674 26868 78680 26920
rect 78732 26908 78738 26920
rect 305730 26908 305736 26920
rect 78732 26880 305736 26908
rect 78732 26868 78738 26880
rect 305730 26868 305736 26880
rect 305788 26868 305794 26920
rect 336826 26188 336832 26240
rect 336884 26228 336890 26240
rect 442994 26228 443000 26240
rect 336884 26200 443000 26228
rect 336884 26188 336890 26200
rect 442994 26188 443000 26200
rect 443052 26188 443058 26240
rect 179322 25644 179328 25696
rect 179380 25684 179386 25696
rect 299474 25684 299480 25696
rect 179380 25656 299480 25684
rect 179380 25644 179386 25656
rect 299474 25644 299480 25656
rect 299532 25684 299538 25696
rect 300762 25684 300768 25696
rect 299532 25656 300768 25684
rect 299532 25644 299538 25656
rect 300762 25644 300768 25656
rect 300820 25644 300826 25696
rect 82814 25576 82820 25628
rect 82872 25616 82878 25628
rect 273898 25616 273904 25628
rect 82872 25588 273904 25616
rect 82872 25576 82878 25588
rect 273898 25576 273904 25588
rect 273956 25576 273962 25628
rect 4154 25508 4160 25560
rect 4212 25548 4218 25560
rect 298922 25548 298928 25560
rect 4212 25520 298928 25548
rect 4212 25508 4218 25520
rect 298922 25508 298928 25520
rect 298980 25508 298986 25560
rect 305638 25508 305644 25560
rect 305696 25548 305702 25560
rect 378870 25548 378876 25560
rect 305696 25520 378876 25548
rect 305696 25508 305702 25520
rect 378870 25508 378876 25520
rect 378928 25508 378934 25560
rect 300762 24760 300768 24812
rect 300820 24800 300826 24812
rect 369118 24800 369124 24812
rect 300820 24772 369124 24800
rect 300820 24760 300826 24772
rect 369118 24760 369124 24772
rect 369176 24760 369182 24812
rect 113174 24080 113180 24132
rect 113232 24120 113238 24132
rect 250438 24120 250444 24132
rect 113232 24092 250444 24120
rect 113232 24080 113238 24092
rect 250438 24080 250444 24092
rect 250496 24080 250502 24132
rect 176562 23400 176568 23452
rect 176620 23440 176626 23452
rect 331214 23440 331220 23452
rect 176620 23412 331220 23440
rect 176620 23400 176626 23412
rect 331214 23400 331220 23412
rect 331272 23400 331278 23452
rect 331214 22924 331220 22976
rect 331272 22964 331278 22976
rect 332042 22964 332048 22976
rect 331272 22936 332048 22964
rect 331272 22924 331278 22936
rect 332042 22924 332048 22936
rect 332100 22924 332106 22976
rect 52546 22788 52552 22840
rect 52604 22828 52610 22840
rect 293218 22828 293224 22840
rect 52604 22800 293224 22828
rect 52604 22788 52610 22800
rect 293218 22788 293224 22800
rect 293276 22788 293282 22840
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 268378 22760 268384 22772
rect 12492 22732 268384 22760
rect 12492 22720 12498 22732
rect 268378 22720 268384 22732
rect 268436 22720 268442 22772
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 249794 22080 249800 22092
rect 1360 22052 249800 22080
rect 1360 22040 1366 22052
rect 249794 22040 249800 22052
rect 249852 22040 249858 22092
rect 314654 22040 314660 22092
rect 314712 22080 314718 22092
rect 392578 22080 392584 22092
rect 314712 22052 392584 22080
rect 314712 22040 314718 22052
rect 392578 22040 392584 22052
rect 392636 22040 392642 22092
rect 14 21564 20 21616
rect 72 21604 78 21616
rect 1302 21604 1308 21616
rect 72 21576 1308 21604
rect 72 21564 78 21576
rect 1302 21564 1308 21576
rect 1360 21564 1366 21616
rect 281534 21428 281540 21480
rect 281592 21468 281598 21480
rect 314654 21468 314660 21480
rect 281592 21440 314660 21468
rect 281592 21428 281598 21440
rect 314654 21428 314660 21440
rect 314712 21428 314718 21480
rect 111794 21360 111800 21412
rect 111852 21400 111858 21412
rect 307018 21400 307024 21412
rect 111852 21372 307024 21400
rect 111852 21360 111858 21372
rect 307018 21360 307024 21372
rect 307076 21360 307082 21412
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 22738 20652 22744 20664
rect 3568 20624 22744 20652
rect 3568 20612 3574 20624
rect 22738 20612 22744 20624
rect 22796 20612 22802 20664
rect 274634 20612 274640 20664
rect 274692 20652 274698 20664
rect 275830 20652 275836 20664
rect 274692 20624 275836 20652
rect 274692 20612 274698 20624
rect 275830 20612 275836 20624
rect 275888 20652 275894 20664
rect 420914 20652 420920 20664
rect 275888 20624 420920 20652
rect 275888 20612 275894 20624
rect 420914 20612 420920 20624
rect 420972 20612 420978 20664
rect 498838 20612 498844 20664
rect 498896 20652 498902 20664
rect 579890 20652 579896 20664
rect 498896 20624 579896 20652
rect 498896 20612 498902 20624
rect 579890 20612 579896 20624
rect 579948 20612 579954 20664
rect 102134 20000 102140 20052
rect 102192 20040 102198 20052
rect 300118 20040 300124 20052
rect 102192 20012 300124 20040
rect 102192 20000 102198 20012
rect 300118 20000 300124 20012
rect 300176 20000 300182 20052
rect 57974 19932 57980 19984
rect 58032 19972 58038 19984
rect 287882 19972 287888 19984
rect 58032 19944 287888 19972
rect 58032 19932 58038 19944
rect 287882 19932 287888 19944
rect 287940 19932 287946 19984
rect 176470 19252 176476 19304
rect 176528 19292 176534 19304
rect 244274 19292 244280 19304
rect 176528 19264 244280 19292
rect 176528 19252 176534 19264
rect 244274 19252 244280 19264
rect 244332 19292 244338 19304
rect 244918 19292 244924 19304
rect 244332 19264 244924 19292
rect 244332 19252 244338 19264
rect 244918 19252 244924 19264
rect 244976 19252 244982 19304
rect 289722 19252 289728 19304
rect 289780 19292 289786 19304
rect 396718 19292 396724 19304
rect 289780 19264 396724 19292
rect 289780 19252 289786 19264
rect 396718 19252 396724 19264
rect 396776 19252 396782 19304
rect 188982 18640 188988 18692
rect 189040 18680 189046 18692
rect 260834 18680 260840 18692
rect 189040 18652 260840 18680
rect 189040 18640 189046 18652
rect 260834 18640 260840 18652
rect 260892 18640 260898 18692
rect 93946 18572 93952 18624
rect 94004 18612 94010 18624
rect 283558 18612 283564 18624
rect 94004 18584 283564 18612
rect 94004 18572 94010 18584
rect 283558 18572 283564 18584
rect 283616 18572 283622 18624
rect 263594 17960 263600 18012
rect 263652 18000 263658 18012
rect 289722 18000 289728 18012
rect 263652 17972 289728 18000
rect 263652 17960 263658 17972
rect 289722 17960 289728 17972
rect 289780 17960 289786 18012
rect 210418 17348 210424 17400
rect 210476 17388 210482 17400
rect 210476 17360 259592 17388
rect 210476 17348 210482 17360
rect 259564 17332 259592 17360
rect 96614 17280 96620 17332
rect 96672 17320 96678 17332
rect 258810 17320 258816 17332
rect 96672 17292 258816 17320
rect 96672 17280 96678 17292
rect 258810 17280 258816 17292
rect 258868 17280 258874 17332
rect 259546 17280 259552 17332
rect 259604 17320 259610 17332
rect 377398 17320 377404 17332
rect 259604 17292 377404 17320
rect 259604 17280 259610 17292
rect 377398 17280 377404 17292
rect 377456 17280 377462 17332
rect 104894 17212 104900 17264
rect 104952 17252 104958 17264
rect 289170 17252 289176 17264
rect 104952 17224 289176 17252
rect 104952 17212 104958 17224
rect 289170 17212 289176 17224
rect 289228 17212 289234 17264
rect 179506 15988 179512 16040
rect 179564 16028 179570 16040
rect 294874 16028 294880 16040
rect 179564 16000 294880 16028
rect 179564 15988 179570 16000
rect 294874 15988 294880 16000
rect 294932 16028 294938 16040
rect 296162 16028 296168 16040
rect 294932 16000 296168 16028
rect 294932 15988 294938 16000
rect 296162 15988 296168 16000
rect 296220 15988 296226 16040
rect 50154 15920 50160 15972
rect 50212 15960 50218 15972
rect 257338 15960 257344 15972
rect 50212 15932 257344 15960
rect 50212 15920 50218 15932
rect 257338 15920 257344 15932
rect 257396 15920 257402 15972
rect 275922 15920 275928 15972
rect 275980 15960 275986 15972
rect 277946 15960 277952 15972
rect 275980 15932 277952 15960
rect 275980 15920 275986 15932
rect 277946 15920 277952 15932
rect 278004 15960 278010 15972
rect 449894 15960 449900 15972
rect 278004 15932 449900 15960
rect 278004 15920 278010 15932
rect 449894 15920 449900 15932
rect 449952 15920 449958 15972
rect 69842 15852 69848 15904
rect 69900 15892 69906 15904
rect 282362 15892 282368 15904
rect 69900 15864 282368 15892
rect 69900 15852 69906 15864
rect 282362 15852 282368 15864
rect 282420 15852 282426 15904
rect 266354 15104 266360 15156
rect 266412 15144 266418 15156
rect 385678 15144 385684 15156
rect 266412 15116 385684 15144
rect 266412 15104 266418 15116
rect 385678 15104 385684 15116
rect 385736 15104 385742 15156
rect 108114 14492 108120 14544
rect 108172 14532 108178 14544
rect 253290 14532 253296 14544
rect 108172 14504 253296 14532
rect 108172 14492 108178 14504
rect 253290 14492 253296 14504
rect 253348 14492 253354 14544
rect 84194 14424 84200 14476
rect 84252 14464 84258 14476
rect 301498 14464 301504 14476
rect 84252 14436 301504 14464
rect 84252 14424 84258 14436
rect 301498 14424 301504 14436
rect 301556 14424 301562 14476
rect 271782 13744 271788 13796
rect 271840 13784 271846 13796
rect 360930 13784 360936 13796
rect 271840 13756 360936 13784
rect 271840 13744 271846 13756
rect 360930 13744 360936 13756
rect 360988 13744 360994 13796
rect 249978 13200 249984 13252
rect 250036 13240 250042 13252
rect 266354 13240 266360 13252
rect 250036 13212 266360 13240
rect 250036 13200 250042 13212
rect 266354 13200 266360 13212
rect 266412 13200 266418 13252
rect 177942 13132 177948 13184
rect 178000 13172 178006 13184
rect 284938 13172 284944 13184
rect 178000 13144 284944 13172
rect 178000 13132 178006 13144
rect 284938 13132 284944 13144
rect 284996 13132 285002 13184
rect 109034 13064 109040 13116
rect 109092 13104 109098 13116
rect 258718 13104 258724 13116
rect 109092 13076 258724 13104
rect 109092 13064 109098 13076
rect 258718 13064 258724 13076
rect 258776 13064 258782 13116
rect 348418 13064 348424 13116
rect 348476 13104 348482 13116
rect 449066 13104 449072 13116
rect 348476 13076 449072 13104
rect 348476 13064 348482 13076
rect 449066 13064 449072 13076
rect 449124 13064 449130 13116
rect 270770 12452 270776 12504
rect 270828 12492 270834 12504
rect 271782 12492 271788 12504
rect 270828 12464 271788 12492
rect 270828 12452 270834 12464
rect 271782 12452 271788 12464
rect 271840 12452 271846 12504
rect 285674 12384 285680 12436
rect 285732 12424 285738 12436
rect 286962 12424 286968 12436
rect 285732 12396 286968 12424
rect 285732 12384 285738 12396
rect 286962 12384 286968 12396
rect 287020 12424 287026 12436
rect 450078 12424 450084 12436
rect 287020 12396 450084 12424
rect 287020 12384 287026 12396
rect 450078 12384 450084 12396
rect 450136 12384 450142 12436
rect 256694 11840 256700 11892
rect 256752 11880 256758 11892
rect 285674 11880 285680 11892
rect 256752 11852 285680 11880
rect 256752 11840 256758 11852
rect 285674 11840 285680 11852
rect 285732 11840 285738 11892
rect 28442 11772 28448 11824
rect 28500 11812 28506 11824
rect 264238 11812 264244 11824
rect 28500 11784 264244 11812
rect 28500 11772 28506 11784
rect 264238 11772 264244 11784
rect 264296 11772 264302 11824
rect 34514 11704 34520 11756
rect 34572 11744 34578 11756
rect 294598 11744 294604 11756
rect 34572 11716 294604 11744
rect 34572 11704 34578 11716
rect 294598 11704 294604 11716
rect 294656 11704 294662 11756
rect 183554 10956 183560 11008
rect 183612 10996 183618 11008
rect 349154 10996 349160 11008
rect 183612 10968 349160 10996
rect 183612 10956 183618 10968
rect 349154 10956 349160 10968
rect 349212 10996 349218 11008
rect 349798 10996 349804 11008
rect 349212 10968 349804 10996
rect 349212 10956 349218 10968
rect 349798 10956 349804 10968
rect 349856 10956 349862 11008
rect 345290 10888 345296 10940
rect 345348 10928 345354 10940
rect 345750 10928 345756 10940
rect 345348 10900 345756 10928
rect 345348 10888 345354 10900
rect 345750 10888 345756 10900
rect 345808 10928 345814 10940
rect 400858 10928 400864 10940
rect 345808 10900 400864 10928
rect 345808 10888 345814 10900
rect 400858 10888 400864 10900
rect 400916 10888 400922 10940
rect 120626 10276 120632 10328
rect 120684 10316 120690 10328
rect 253198 10316 253204 10328
rect 120684 10288 253204 10316
rect 120684 10276 120690 10288
rect 253198 10276 253204 10288
rect 253256 10276 253262 10328
rect 287974 9596 287980 9648
rect 288032 9636 288038 9648
rect 429838 9636 429844 9648
rect 288032 9608 429844 9636
rect 288032 9596 288038 9608
rect 429838 9596 429844 9608
rect 429896 9596 429902 9648
rect 123478 9052 123484 9104
rect 123536 9092 123542 9104
rect 275278 9092 275284 9104
rect 123536 9064 275284 9092
rect 123536 9052 123542 9064
rect 275278 9052 275284 9064
rect 275336 9052 275342 9104
rect 119890 8984 119896 9036
rect 119948 9024 119954 9036
rect 291930 9024 291936 9036
rect 119948 8996 291936 9024
rect 119948 8984 119954 8996
rect 291930 8984 291936 8996
rect 291988 8984 291994 9036
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 295978 8956 295984 8968
rect 23072 8928 295984 8956
rect 23072 8916 23078 8928
rect 295978 8916 295984 8928
rect 296036 8916 296042 8968
rect 349430 8236 349436 8288
rect 349488 8276 349494 8288
rect 349706 8276 349712 8288
rect 349488 8248 349712 8276
rect 349488 8236 349494 8248
rect 349706 8236 349712 8248
rect 349764 8276 349770 8288
rect 412634 8276 412640 8288
rect 349764 8248 412640 8276
rect 349764 8236 349770 8248
rect 412634 8236 412640 8248
rect 412692 8236 412698 8288
rect 309870 8168 309876 8220
rect 309928 8208 309934 8220
rect 356790 8208 356796 8220
rect 309928 8180 356796 8208
rect 309928 8168 309934 8180
rect 356790 8168 356796 8180
rect 356848 8168 356854 8220
rect 115198 7624 115204 7676
rect 115256 7664 115262 7676
rect 304258 7664 304264 7676
rect 115256 7636 304264 7664
rect 115256 7624 115262 7636
rect 304258 7624 304264 7636
rect 304316 7624 304322 7676
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 249058 7596 249064 7608
rect 4120 7568 249064 7596
rect 4120 7556 4126 7568
rect 249058 7556 249064 7568
rect 249116 7556 249122 7608
rect 293678 7556 293684 7608
rect 293736 7596 293742 7608
rect 309226 7596 309232 7608
rect 293736 7568 309232 7596
rect 293736 7556 293742 7568
rect 309226 7556 309232 7568
rect 309284 7596 309290 7608
rect 309870 7596 309876 7608
rect 309284 7568 309876 7596
rect 309284 7556 309290 7568
rect 309870 7556 309876 7568
rect 309928 7556 309934 7608
rect 327074 7556 327080 7608
rect 327132 7596 327138 7608
rect 349706 7596 349712 7608
rect 327132 7568 349712 7596
rect 327132 7556 327138 7568
rect 349706 7556 349712 7568
rect 349764 7556 349770 7608
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 31018 6848 31024 6860
rect 3568 6820 31024 6848
rect 3568 6808 3574 6820
rect 31018 6808 31024 6820
rect 31076 6808 31082 6860
rect 324958 6808 324964 6860
rect 325016 6848 325022 6860
rect 414014 6848 414020 6860
rect 325016 6820 414020 6848
rect 325016 6808 325022 6820
rect 414014 6808 414020 6820
rect 414072 6808 414078 6860
rect 418798 6808 418804 6860
rect 418856 6848 418862 6860
rect 580166 6848 580172 6860
rect 418856 6820 580172 6848
rect 418856 6808 418862 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 347038 6740 347044 6792
rect 347096 6780 347102 6792
rect 348418 6780 348424 6792
rect 347096 6752 348424 6780
rect 347096 6740 347102 6752
rect 348418 6740 348424 6752
rect 348476 6740 348482 6792
rect 175182 6264 175188 6316
rect 175240 6304 175246 6316
rect 302050 6304 302056 6316
rect 175240 6276 302056 6304
rect 175240 6264 175246 6276
rect 302050 6264 302056 6276
rect 302108 6264 302114 6316
rect 116394 6196 116400 6248
rect 116452 6236 116458 6248
rect 302878 6236 302884 6248
rect 116452 6208 302884 6236
rect 116452 6196 116458 6208
rect 302878 6196 302884 6208
rect 302936 6196 302942 6248
rect 60826 6128 60832 6180
rect 60884 6168 60890 6180
rect 287698 6168 287704 6180
rect 60884 6140 287704 6168
rect 60884 6128 60890 6140
rect 287698 6128 287704 6140
rect 287756 6128 287762 6180
rect 324406 5516 324412 5568
rect 324464 5556 324470 5568
rect 324958 5556 324964 5568
rect 324464 5528 324964 5556
rect 324464 5516 324470 5528
rect 324958 5516 324964 5528
rect 325016 5516 325022 5568
rect 77386 4904 77392 4956
rect 77444 4944 77450 4956
rect 77444 4916 84194 4944
rect 77444 4904 77450 4916
rect 84166 4876 84194 4916
rect 261478 4876 261484 4888
rect 84166 4848 261484 4876
rect 261478 4836 261484 4848
rect 261536 4836 261542 4888
rect 56042 4768 56048 4820
rect 56100 4808 56106 4820
rect 254578 4808 254584 4820
rect 56100 4780 254584 4808
rect 56100 4768 56106 4780
rect 254578 4768 254584 4780
rect 254636 4768 254642 4820
rect 289722 4768 289728 4820
rect 289780 4808 289786 4820
rect 395338 4808 395344 4820
rect 289780 4780 395344 4808
rect 289780 4768 289786 4780
rect 395338 4768 395344 4780
rect 395396 4768 395402 4820
rect 215938 4088 215944 4140
rect 215996 4128 216002 4140
rect 247586 4128 247592 4140
rect 215996 4100 247592 4128
rect 215996 4088 216002 4100
rect 247586 4088 247592 4100
rect 247644 4088 247650 4140
rect 291838 4088 291844 4140
rect 291896 4128 291902 4140
rect 298462 4128 298468 4140
rect 291896 4100 298468 4128
rect 291896 4088 291902 4100
rect 298462 4088 298468 4100
rect 298520 4088 298526 4140
rect 302050 4088 302056 4140
rect 302108 4128 302114 4140
rect 329190 4128 329196 4140
rect 302108 4100 329196 4128
rect 302108 4088 302114 4100
rect 329190 4088 329196 4100
rect 329248 4088 329254 4140
rect 351178 4088 351184 4140
rect 351236 4128 351242 4140
rect 351638 4128 351644 4140
rect 351236 4100 351644 4128
rect 351236 4088 351242 4100
rect 351638 4088 351644 4100
rect 351696 4128 351702 4140
rect 403618 4128 403624 4140
rect 351696 4100 403624 4128
rect 351696 4088 351702 4100
rect 403618 4088 403624 4100
rect 403676 4088 403682 4140
rect 282178 4020 282184 4072
rect 282236 4060 282242 4072
rect 291378 4060 291384 4072
rect 282236 4032 291384 4060
rect 282236 4020 282242 4032
rect 291378 4020 291384 4032
rect 291436 4060 291442 4072
rect 292022 4060 292028 4072
rect 291436 4032 292028 4060
rect 291436 4020 291442 4032
rect 292022 4020 292028 4032
rect 292080 4020 292086 4072
rect 305638 4020 305644 4072
rect 305696 4060 305702 4072
rect 306742 4060 306748 4072
rect 305696 4032 306748 4060
rect 305696 4020 305702 4032
rect 306742 4020 306748 4032
rect 306800 4020 306806 4072
rect 278682 3952 278688 4004
rect 278740 3992 278746 4004
rect 288986 3992 288992 4004
rect 278740 3964 288992 3992
rect 278740 3952 278746 3964
rect 288986 3952 288992 3964
rect 289044 3992 289050 4004
rect 289722 3992 289728 4004
rect 289044 3964 289728 3992
rect 289044 3952 289050 3964
rect 289722 3952 289728 3964
rect 289780 3952 289786 4004
rect 286594 3816 286600 3868
rect 286652 3856 286658 3868
rect 289078 3856 289084 3868
rect 286652 3828 289084 3856
rect 286652 3816 286658 3828
rect 289078 3816 289084 3828
rect 289136 3816 289142 3868
rect 132954 3612 132960 3664
rect 133012 3652 133018 3664
rect 203518 3652 203524 3664
rect 133012 3624 203524 3652
rect 133012 3612 133018 3624
rect 203518 3612 203524 3624
rect 203576 3612 203582 3664
rect 331858 3652 331864 3664
rect 327644 3624 331864 3652
rect 52454 3544 52460 3596
rect 52512 3584 52518 3596
rect 53374 3584 53380 3596
rect 52512 3556 53380 3584
rect 52512 3544 52518 3556
rect 53374 3544 53380 3556
rect 53432 3544 53438 3596
rect 85574 3544 85580 3596
rect 85632 3584 85638 3596
rect 86494 3584 86500 3596
rect 85632 3556 86500 3584
rect 85632 3544 85638 3556
rect 86494 3544 86500 3556
rect 86552 3544 86558 3596
rect 103330 3544 103336 3596
rect 103388 3584 103394 3596
rect 214558 3584 214564 3596
rect 103388 3556 214564 3584
rect 103388 3544 103394 3556
rect 214558 3544 214564 3556
rect 214616 3544 214622 3596
rect 242986 3544 242992 3596
rect 243044 3584 243050 3596
rect 278038 3584 278044 3596
rect 243044 3556 248414 3584
rect 243044 3544 243050 3556
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 192478 3516 192484 3528
rect 41932 3488 192484 3516
rect 41932 3476 41938 3488
rect 192478 3476 192484 3488
rect 192536 3476 192542 3528
rect 235810 3476 235816 3528
rect 235868 3516 235874 3528
rect 238018 3516 238024 3528
rect 235868 3488 238024 3516
rect 235868 3476 235874 3488
rect 238018 3476 238024 3488
rect 238076 3476 238082 3528
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 244090 3516 244096 3528
rect 242952 3488 244096 3516
rect 242952 3476 242958 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 248386 3516 248414 3556
rect 277366 3556 278044 3584
rect 276658 3516 276664 3528
rect 248386 3488 276664 3516
rect 276658 3476 276664 3488
rect 276716 3476 276722 3528
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 185578 3448 185584 3460
rect 25372 3420 185584 3448
rect 25372 3408 25378 3420
rect 185578 3408 185584 3420
rect 185636 3408 185642 3460
rect 206278 3408 206284 3460
rect 206336 3448 206342 3460
rect 268838 3448 268844 3460
rect 206336 3420 268844 3448
rect 206336 3408 206342 3420
rect 268838 3408 268844 3420
rect 268896 3408 268902 3460
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 135254 3340 135260 3392
rect 135312 3380 135318 3392
rect 136450 3380 136456 3392
rect 135312 3352 136456 3380
rect 135312 3340 135318 3352
rect 136450 3340 136456 3352
rect 136508 3340 136514 3392
rect 277118 3272 277124 3324
rect 277176 3312 277182 3324
rect 277366 3312 277394 3556
rect 278038 3544 278044 3556
rect 278096 3544 278102 3596
rect 299566 3544 299572 3596
rect 299624 3584 299630 3596
rect 300762 3584 300768 3596
rect 299624 3556 300768 3584
rect 299624 3544 299630 3556
rect 300762 3544 300768 3556
rect 300820 3544 300826 3596
rect 309042 3544 309048 3596
rect 309100 3584 309106 3596
rect 311158 3584 311164 3596
rect 309100 3556 311164 3584
rect 309100 3544 309106 3556
rect 311158 3544 311164 3556
rect 311216 3544 311222 3596
rect 316034 3544 316040 3596
rect 316092 3584 316098 3596
rect 317322 3584 317328 3596
rect 316092 3556 317328 3584
rect 316092 3544 316098 3556
rect 317322 3544 317328 3556
rect 317380 3544 317386 3596
rect 322106 3544 322112 3596
rect 322164 3584 322170 3596
rect 327074 3584 327080 3596
rect 322164 3556 327080 3584
rect 322164 3544 322170 3556
rect 327074 3544 327080 3556
rect 327132 3544 327138 3596
rect 284294 3476 284300 3528
rect 284352 3516 284358 3528
rect 284938 3516 284944 3528
rect 284352 3488 284944 3516
rect 284352 3476 284358 3488
rect 284938 3476 284944 3488
rect 284996 3476 285002 3528
rect 298002 3476 298008 3528
rect 298060 3516 298066 3528
rect 315022 3516 315028 3528
rect 298060 3488 315028 3516
rect 298060 3476 298066 3488
rect 315022 3476 315028 3488
rect 315080 3476 315086 3528
rect 315298 3476 315304 3528
rect 315356 3516 315362 3528
rect 316218 3516 316224 3528
rect 315356 3488 316224 3516
rect 315356 3476 315362 3488
rect 316218 3476 316224 3488
rect 316276 3516 316282 3528
rect 327644 3516 327672 3624
rect 331858 3612 331864 3624
rect 331916 3612 331922 3664
rect 340966 3612 340972 3664
rect 341024 3652 341030 3664
rect 342162 3652 342168 3664
rect 341024 3624 342168 3652
rect 341024 3612 341030 3624
rect 342162 3612 342168 3624
rect 342220 3612 342226 3664
rect 327718 3544 327724 3596
rect 327776 3544 327782 3596
rect 335998 3544 336004 3596
rect 336056 3584 336062 3596
rect 344554 3584 344560 3596
rect 336056 3556 344560 3584
rect 336056 3544 336062 3556
rect 344554 3544 344560 3556
rect 344612 3584 344618 3596
rect 344612 3556 345014 3584
rect 344612 3544 344618 3556
rect 316276 3488 327672 3516
rect 316276 3476 316282 3488
rect 305546 3408 305552 3460
rect 305604 3448 305610 3460
rect 327736 3448 327764 3544
rect 332594 3476 332600 3528
rect 332652 3516 332658 3528
rect 333882 3516 333888 3528
rect 332652 3488 333888 3516
rect 332652 3476 332658 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 340966 3476 340972 3528
rect 341024 3516 341030 3528
rect 341518 3516 341524 3528
rect 341024 3488 341524 3516
rect 341024 3476 341030 3488
rect 341518 3476 341524 3488
rect 341576 3476 341582 3528
rect 305604 3420 327764 3448
rect 344986 3448 345014 3556
rect 349246 3476 349252 3528
rect 349304 3516 349310 3528
rect 350442 3516 350448 3528
rect 349304 3488 350448 3516
rect 349304 3476 349310 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 355318 3448 355324 3460
rect 344986 3420 355324 3448
rect 305604 3408 305610 3420
rect 355318 3408 355324 3420
rect 355376 3408 355382 3460
rect 324314 3340 324320 3392
rect 324372 3380 324378 3392
rect 325602 3380 325608 3392
rect 324372 3352 325608 3380
rect 324372 3340 324378 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 277176 3284 277394 3312
rect 277176 3272 277182 3284
rect 271138 3000 271144 3052
rect 271196 3040 271202 3052
rect 276014 3040 276020 3052
rect 271196 3012 276020 3040
rect 271196 3000 271202 3012
rect 276014 3000 276020 3012
rect 276072 3000 276078 3052
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 3418 2972 3424 2984
rect 1728 2944 3424 2972
rect 1728 2932 1734 2944
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 40678 2048 40684 2100
rect 40736 2088 40742 2100
rect 294690 2088 294696 2100
rect 40736 2060 294696 2088
rect 40736 2048 40742 2060
rect 294690 2048 294696 2060
rect 294748 2048 294754 2100
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 63408 702788 63460 702840
rect 218980 702788 219032 702840
rect 412640 702788 412692 702840
rect 413652 702788 413704 702840
rect 72976 702720 73028 702772
rect 245660 702720 245712 702772
rect 53748 702652 53800 702704
rect 202788 702652 202840 702704
rect 416780 702652 416832 702704
rect 40500 702584 40552 702636
rect 217324 702584 217376 702636
rect 300124 702584 300176 702636
rect 538220 702584 538272 702636
rect 8116 702516 8168 702568
rect 210424 702516 210476 702568
rect 251088 702516 251140 702568
rect 527180 702516 527232 702568
rect 130384 702448 130436 702500
rect 412640 702448 412692 702500
rect 235172 700340 235224 700392
rect 269120 700340 269172 700392
rect 359464 700340 359516 700392
rect 397460 700340 397512 700392
rect 24308 700272 24360 700324
rect 39304 700272 39356 700324
rect 52368 700272 52420 700324
rect 137836 700272 137888 700324
rect 154120 700272 154172 700324
rect 247040 700272 247092 700324
rect 332416 700272 332468 700324
rect 429844 700272 429896 700324
rect 494796 700272 494848 700324
rect 518164 700272 518216 700324
rect 102784 699660 102836 699712
rect 105452 699660 105504 699712
rect 261484 699660 261536 699712
rect 300124 699660 300176 699712
rect 348792 699660 348844 699712
rect 351184 699660 351236 699712
rect 540244 699660 540296 699712
rect 543464 699660 543516 699712
rect 552664 699660 552716 699712
rect 559656 699660 559708 699712
rect 265624 698912 265676 698964
rect 348792 698912 348844 698964
rect 570604 696940 570656 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 7564 683136 7616 683188
rect 549904 683136 549956 683188
rect 580172 683136 580224 683188
rect 543004 670692 543056 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 18604 656888 18656 656940
rect 338764 643084 338816 643136
rect 580172 643084 580224 643136
rect 351184 632680 351236 632732
rect 488540 632680 488592 632732
rect 3424 632068 3476 632120
rect 17224 632068 17276 632120
rect 337936 630640 337988 630692
rect 580172 630640 580224 630692
rect 39304 620236 39356 620288
rect 51080 620236 51132 620288
rect 220728 620236 220780 620288
rect 282920 620236 282972 620288
rect 51080 619624 51132 619676
rect 52276 619624 52328 619676
rect 185584 619624 185636 619676
rect 88340 618876 88392 618928
rect 236644 618876 236696 618928
rect 412640 618876 412692 618928
rect 534356 618876 534408 618928
rect 3148 618264 3200 618316
rect 40684 618264 40736 618316
rect 289728 618264 289780 618316
rect 456800 618264 456852 618316
rect 17224 617516 17276 617568
rect 229100 617516 229152 617568
rect 391020 616836 391072 616888
rect 580172 616836 580224 616888
rect 358084 616700 358136 616752
rect 359464 616700 359516 616752
rect 227628 616088 227680 616140
rect 331220 616088 331272 616140
rect 400864 616088 400916 616140
rect 552664 616088 552716 616140
rect 260104 615476 260156 615528
rect 510620 615476 510672 615528
rect 169760 614728 169812 614780
rect 245844 614728 245896 614780
rect 288348 614184 288400 614236
rect 483848 614184 483900 614236
rect 229468 614116 229520 614168
rect 264244 614116 264296 614168
rect 536932 614116 536984 614168
rect 338028 613368 338080 613420
rect 364340 613368 364392 613420
rect 420184 613368 420236 613420
rect 477500 613368 477552 613420
rect 289084 612824 289136 612876
rect 390560 612824 390612 612876
rect 391020 612824 391072 612876
rect 300216 612756 300268 612808
rect 493508 612756 493560 612808
rect 537024 612688 537076 612740
rect 540244 612688 540296 612740
rect 275284 611464 275336 611516
rect 402980 611464 403032 611516
rect 327908 611396 327960 611448
rect 537024 611396 537076 611448
rect 178684 611328 178736 611380
rect 450360 611328 450412 611380
rect 292396 610104 292448 610156
rect 388536 610104 388588 610156
rect 223028 610036 223080 610088
rect 249800 610036 249852 610088
rect 491300 610036 491352 610088
rect 191104 609968 191156 610020
rect 469680 609968 469732 610020
rect 273904 608744 273956 608796
rect 431960 608744 432012 608796
rect 207572 608676 207624 608728
rect 253940 608676 253992 608728
rect 436192 608676 436244 608728
rect 232688 608608 232740 608660
rect 252560 608608 252612 608660
rect 498660 608608 498712 608660
rect 462320 607860 462372 607912
rect 534264 607860 534316 607912
rect 306288 607384 306340 607436
rect 452936 607384 452988 607436
rect 169024 607316 169076 607368
rect 412640 607316 412692 607368
rect 295984 607248 296036 607300
rect 562324 607248 562376 607300
rect 63132 607180 63184 607232
rect 443276 607180 443328 607232
rect 319444 606092 319496 606144
rect 378876 606092 378928 606144
rect 324228 606024 324280 606076
rect 448520 606024 448572 606076
rect 333336 605956 333388 606008
rect 520280 605956 520332 606008
rect 119344 605888 119396 605940
rect 409880 605888 409932 605940
rect 3240 605820 3292 605872
rect 46204 605820 46256 605872
rect 63500 605820 63552 605872
rect 459560 605820 459612 605872
rect 357440 605140 357492 605192
rect 358084 605140 358136 605192
rect 332508 604732 332560 604784
rect 400220 604732 400272 604784
rect 400864 604732 400916 604784
rect 287704 604664 287756 604716
rect 357440 604664 357492 604716
rect 308404 604596 308456 604648
rect 386420 604596 386472 604648
rect 166264 604528 166316 604580
rect 312544 604528 312596 604580
rect 396080 604528 396132 604580
rect 86224 604460 86276 604512
rect 524420 604460 524472 604512
rect 321468 603304 321520 603356
rect 423956 603304 424008 603356
rect 204352 603168 204404 603220
rect 251180 603236 251232 603288
rect 414388 603236 414440 603288
rect 252468 603168 252520 603220
rect 486884 603168 486936 603220
rect 63316 603100 63368 603152
rect 381452 603100 381504 603152
rect 283564 602012 283616 602064
rect 376760 602012 376812 602064
rect 298008 601944 298060 601996
rect 398196 601944 398248 601996
rect 339040 601876 339092 601928
rect 496084 601876 496136 601928
rect 317236 601808 317288 601860
rect 536840 601808 536892 601860
rect 305644 601740 305696 601792
rect 549260 601740 549312 601792
rect 549904 601740 549956 601792
rect 112444 601672 112496 601724
rect 440700 601672 440752 601724
rect 307024 600652 307076 600704
rect 393320 600652 393372 600704
rect 336648 600584 336700 600636
rect 474188 600584 474240 600636
rect 334808 600516 334860 600568
rect 500960 600516 501012 600568
rect 253204 600448 253256 600500
rect 438860 600448 438912 600500
rect 134524 600380 134576 600432
rect 349896 600380 349948 600432
rect 17224 600312 17276 600364
rect 374000 600312 374052 600364
rect 376760 600312 376812 600364
rect 544476 600312 544528 600364
rect 331864 599292 331916 599344
rect 347964 599292 348016 599344
rect 311808 599224 311860 599276
rect 371792 599224 371844 599276
rect 327816 599156 327868 599208
rect 415400 599156 415452 599208
rect 327724 599088 327776 599140
rect 422300 599088 422352 599140
rect 512828 599088 512880 599140
rect 542452 599088 542504 599140
rect 334716 599020 334768 599072
rect 537024 599020 537076 599072
rect 80704 598952 80756 599004
rect 534080 598952 534132 599004
rect 414388 598204 414440 598256
rect 482008 598204 482060 598256
rect 140228 597864 140280 597916
rect 407304 597864 407356 597916
rect 518164 597864 518216 597916
rect 552020 597864 552072 597916
rect 333428 597796 333480 597848
rect 345480 597796 345532 597848
rect 503628 597796 503680 597848
rect 547880 597796 547932 597848
rect 326436 597728 326488 597780
rect 367100 597728 367152 597780
rect 477408 597728 477460 597780
rect 538312 597728 538364 597780
rect 339684 597660 339736 597712
rect 405740 597660 405792 597712
rect 472992 597660 473044 597712
rect 543740 597660 543792 597712
rect 279424 597592 279476 597644
rect 369308 597592 369360 597644
rect 486884 597592 486936 597644
rect 574744 597592 574796 597644
rect 407028 597524 407080 597576
rect 527180 597524 527232 597576
rect 532608 597524 532660 597576
rect 561680 597524 561732 597576
rect 236000 597456 236052 597508
rect 236644 597456 236696 597508
rect 90364 596776 90416 596828
rect 102784 596776 102836 596828
rect 323584 596504 323636 596556
rect 465264 596504 465316 596556
rect 329196 596436 329248 596488
rect 539692 596436 539744 596488
rect 309048 596368 309100 596420
rect 535552 596368 535604 596420
rect 153844 596300 153896 596352
rect 383660 596300 383712 596352
rect 331036 596232 331088 596284
rect 582380 596232 582432 596284
rect 38568 596164 38620 596216
rect 143540 596164 143592 596216
rect 236000 596164 236052 596216
rect 256608 596164 256660 596216
rect 529940 596164 529992 596216
rect 220728 596096 220780 596148
rect 407028 596096 407080 596148
rect 569960 595620 570012 595672
rect 570604 595620 570656 595672
rect 459560 595484 459612 595536
rect 460434 595484 460486 595536
rect 92940 595416 92992 595468
rect 317420 595416 317472 595468
rect 325056 595076 325108 595128
rect 352564 595076 352616 595128
rect 460572 595076 460624 595128
rect 544384 595076 544436 595128
rect 338856 595008 338908 595060
rect 426624 595008 426676 595060
rect 456248 595008 456300 595060
rect 553492 595008 553544 595060
rect 337844 594940 337896 594992
rect 538864 594940 538916 594992
rect 318064 594872 318116 594924
rect 535828 594872 535880 594924
rect 53564 594804 53616 594856
rect 140596 594804 140648 594856
rect 331956 594804 332008 594856
rect 569960 594804 570012 594856
rect 339500 594736 339552 594788
rect 342904 594736 342956 594788
rect 535644 594532 535696 594584
rect 537116 594532 537168 594584
rect 127624 594056 127676 594108
rect 339500 594056 339552 594108
rect 54944 593376 54996 593428
rect 169024 593376 169076 593428
rect 169576 593376 169628 593428
rect 143816 593308 143868 593360
rect 339684 593308 339736 593360
rect 45468 592084 45520 592136
rect 127624 592084 127676 592136
rect 39948 592016 40000 592068
rect 163228 592016 163280 592068
rect 55036 591268 55088 591320
rect 327908 591268 327960 591320
rect 562324 591268 562376 591320
rect 579804 591268 579856 591320
rect 60004 590860 60056 590912
rect 86224 590860 86276 590912
rect 86500 590860 86552 590912
rect 41328 590792 41380 590844
rect 92940 590792 92992 590844
rect 48136 590724 48188 590776
rect 159916 590724 159968 590776
rect 56324 590656 56376 590708
rect 191104 590656 191156 590708
rect 191472 590656 191524 590708
rect 197268 590656 197320 590708
rect 273996 590656 274048 590708
rect 535644 590656 535696 590708
rect 554044 590656 554096 590708
rect 106188 589908 106240 589960
rect 336556 589908 336608 589960
rect 38476 589500 38528 589552
rect 105820 589500 105872 589552
rect 106188 589500 106240 589552
rect 99380 589432 99432 589484
rect 251824 589432 251876 589484
rect 35808 589364 35860 589416
rect 77484 589364 77536 589416
rect 257344 589364 257396 589416
rect 59084 589296 59136 589348
rect 309784 589296 309836 589348
rect 50344 588276 50396 588328
rect 197268 588276 197320 588328
rect 57704 588208 57756 588260
rect 90364 588208 90416 588260
rect 59268 588140 59320 588192
rect 112444 588140 112496 588192
rect 56232 588072 56284 588124
rect 130384 588072 130436 588124
rect 214104 588072 214156 588124
rect 248512 588072 248564 588124
rect 194784 588004 194836 588056
rect 253296 588004 253348 588056
rect 60556 587936 60608 587988
rect 153844 587936 153896 587988
rect 163228 587936 163280 587988
rect 318156 587936 318208 587988
rect 8944 587868 8996 587920
rect 172888 587868 172940 587920
rect 266360 587868 266412 587920
rect 324964 587868 325016 587920
rect 337660 587868 337712 587920
rect 197268 587528 197320 587580
rect 198004 587528 198056 587580
rect 299388 587120 299440 587172
rect 337108 587120 337160 587172
rect 49608 586848 49660 586900
rect 83372 586848 83424 586900
rect 49516 586780 49568 586832
rect 96252 586780 96304 586832
rect 122012 586780 122064 586832
rect 244924 586780 244976 586832
rect 63224 586712 63276 586764
rect 137468 586712 137520 586764
rect 217324 586712 217376 586764
rect 245108 586712 245160 586764
rect 57244 586644 57296 586696
rect 166264 586644 166316 586696
rect 201224 586644 201276 586696
rect 217232 586644 217284 586696
rect 239220 586644 239272 586696
rect 277400 586644 277452 586696
rect 31024 586576 31076 586628
rect 147128 586576 147180 586628
rect 181904 586576 181956 586628
rect 243084 586576 243136 586628
rect 44088 586508 44140 586560
rect 125232 586508 125284 586560
rect 50988 585488 51040 585540
rect 67916 585488 67968 585540
rect 46848 585420 46900 585472
rect 102692 585420 102744 585472
rect 15108 585352 15160 585404
rect 71136 585352 71188 585404
rect 226340 585352 226392 585404
rect 227628 585352 227680 585404
rect 247776 585352 247828 585404
rect 60740 585284 60792 585336
rect 150348 585284 150400 585336
rect 185124 585284 185176 585336
rect 185584 585284 185636 585336
rect 247684 585284 247736 585336
rect 48228 585216 48280 585268
rect 109132 585216 109184 585268
rect 137468 585216 137520 585268
rect 260196 585216 260248 585268
rect 35164 585148 35216 585200
rect 255320 585148 255372 585200
rect 333244 585148 333296 585200
rect 337660 585148 337712 585200
rect 217232 585080 217284 585132
rect 295340 585080 295392 585132
rect 295340 584604 295392 584656
rect 295984 584604 296036 584656
rect 61476 584536 61528 584588
rect 245936 584536 245988 584588
rect 292488 583720 292540 583772
rect 337660 583720 337712 583772
rect 245752 582360 245804 582412
rect 318800 582360 318852 582412
rect 320088 582360 320140 582412
rect 245752 582224 245804 582276
rect 245936 582224 245988 582276
rect 297364 581000 297416 581052
rect 337660 581000 337712 581052
rect 535736 581000 535788 581052
rect 563704 581000 563756 581052
rect 244188 580932 244240 580984
rect 336096 580932 336148 580984
rect 242992 580524 243044 580576
rect 243544 580524 243596 580576
rect 3332 579640 3384 579692
rect 57612 579640 57664 579692
rect 60740 579640 60792 579692
rect 242992 579640 243044 579692
rect 244188 579640 244240 579692
rect 535736 579164 535788 579216
rect 538220 579164 538272 579216
rect 245108 578892 245160 578944
rect 276020 578892 276072 578944
rect 276020 578212 276072 578264
rect 276664 578212 276716 578264
rect 337660 578212 337712 578264
rect 329748 576852 329800 576904
rect 337660 576852 337712 576904
rect 535736 576852 535788 576904
rect 539600 576852 539652 576904
rect 560944 576852 560996 576904
rect 580172 576852 580224 576904
rect 245660 576512 245712 576564
rect 245936 576512 245988 576564
rect 314936 576104 314988 576156
rect 339040 576104 339092 576156
rect 59176 575492 59228 575544
rect 61568 575492 61620 575544
rect 245660 575492 245712 575544
rect 314752 575492 314804 575544
rect 314936 575492 314988 575544
rect 331036 572636 331088 572688
rect 337660 572636 337712 572688
rect 245660 571956 245712 572008
rect 293960 571956 294012 572008
rect 55128 571344 55180 571396
rect 60740 571344 60792 571396
rect 293960 571276 294012 571328
rect 295248 571276 295300 571328
rect 327724 571276 327776 571328
rect 337844 570528 337896 570580
rect 338764 570528 338816 570580
rect 245660 569168 245712 569220
rect 245936 569168 245988 569220
rect 262220 569168 262272 569220
rect 535460 569168 535512 569220
rect 538404 569168 538456 569220
rect 304264 568624 304316 568676
rect 337660 568624 337712 568676
rect 53656 568556 53708 568608
rect 60740 568556 60792 568608
rect 262220 568556 262272 568608
rect 325148 568556 325200 568608
rect 243544 568488 243596 568540
rect 305644 568488 305696 568540
rect 315304 566448 315356 566500
rect 333336 566448 333388 566500
rect 3424 565836 3476 565888
rect 22744 565836 22796 565888
rect 245936 565836 245988 565888
rect 314660 565836 314712 565888
rect 315304 565836 315356 565888
rect 27528 564408 27580 564460
rect 60740 564408 60792 564460
rect 535460 563864 535512 563916
rect 538220 563864 538272 563916
rect 538864 563660 538916 563712
rect 575480 563660 575532 563712
rect 575480 563048 575532 563100
rect 579804 563048 579856 563100
rect 244924 562300 244976 562352
rect 317328 562300 317380 562352
rect 317328 561688 317380 561740
rect 337384 561688 337436 561740
rect 244924 561620 244976 561672
rect 245568 561620 245620 561672
rect 329196 561620 329248 561672
rect 250444 560260 250496 560312
rect 337660 560260 337712 560312
rect 318156 560192 318208 560244
rect 336924 560192 336976 560244
rect 269028 559512 269080 559564
rect 334808 559512 334860 559564
rect 245936 558900 245988 558952
rect 267740 558900 267792 558952
rect 269028 558900 269080 558952
rect 249708 556792 249760 556844
rect 337936 556792 337988 556844
rect 59084 556112 59136 556164
rect 60740 556112 60792 556164
rect 35716 555432 35768 555484
rect 59084 555432 59136 555484
rect 3148 554684 3200 554736
rect 35164 554684 35216 554736
rect 535460 554684 535512 554736
rect 562324 554684 562376 554736
rect 257252 552644 257304 552696
rect 338948 552644 339000 552696
rect 39856 552032 39908 552084
rect 60740 552032 60792 552084
rect 245936 552032 245988 552084
rect 256700 552032 256752 552084
rect 257252 552032 257304 552084
rect 245660 551284 245712 551336
rect 269764 551284 269816 551336
rect 245936 549244 245988 549296
rect 255228 549244 255280 549296
rect 331956 549176 332008 549228
rect 37188 547884 37240 547936
rect 60740 547884 60792 547936
rect 307208 547884 307260 547936
rect 337660 547884 337712 547936
rect 245936 546456 245988 546508
rect 264336 546456 264388 546508
rect 56508 545776 56560 545828
rect 60740 545776 60792 545828
rect 245292 543668 245344 543720
rect 329104 543668 329156 543720
rect 40684 542376 40736 542428
rect 42800 542376 42852 542428
rect 60740 542376 60792 542428
rect 311164 542376 311216 542428
rect 337660 542376 337712 542428
rect 290464 540948 290516 541000
rect 337476 540948 337528 541000
rect 322204 539520 322256 539572
rect 337660 539520 337712 539572
rect 41236 538228 41288 538280
rect 60740 538228 60792 538280
rect 574744 538160 574796 538212
rect 580172 538160 580224 538212
rect 309784 536732 309836 536784
rect 337292 536732 337344 536784
rect 245844 536052 245896 536104
rect 311716 536052 311768 536104
rect 338856 536052 338908 536104
rect 59084 535440 59136 535492
rect 61568 535440 61620 535492
rect 244188 534012 244240 534064
rect 334716 534012 334768 534064
rect 535552 533400 535604 533452
rect 539692 533400 539744 533452
rect 242992 532720 243044 532772
rect 244188 532720 244240 532772
rect 326344 532720 326396 532772
rect 337660 532720 337712 532772
rect 54484 531972 54536 532024
rect 58992 531972 59044 532024
rect 60740 531972 60792 532024
rect 264336 531972 264388 532024
rect 336832 531972 336884 532024
rect 7564 529184 7616 529236
rect 43904 529184 43956 529236
rect 246948 529184 247000 529236
rect 321560 529184 321612 529236
rect 329104 528912 329156 528964
rect 336832 528912 336884 528964
rect 43904 528572 43956 528624
rect 60740 528572 60792 528624
rect 535552 528572 535604 528624
rect 537116 528572 537168 528624
rect 246856 528504 246908 528556
rect 336004 528504 336056 528556
rect 249064 527824 249116 527876
rect 309048 527824 309100 527876
rect 3424 527144 3476 527196
rect 48964 527144 49016 527196
rect 246304 527144 246356 527196
rect 246856 527144 246908 527196
rect 309048 527144 309100 527196
rect 309784 527144 309836 527196
rect 21364 527076 21416 527128
rect 269764 527076 269816 527128
rect 317236 527076 317288 527128
rect 21364 526396 21416 526448
rect 314844 526396 314896 526448
rect 337844 526396 337896 526448
rect 264336 525784 264388 525836
rect 314844 525784 314896 525836
rect 315304 525784 315356 525836
rect 317236 525784 317288 525836
rect 317420 525784 317472 525836
rect 53840 525716 53892 525768
rect 55036 525716 55088 525768
rect 60740 525716 60792 525768
rect 544476 525716 544528 525768
rect 579804 525716 579856 525768
rect 33048 525036 33100 525088
rect 53840 525036 53892 525088
rect 300124 525036 300176 525088
rect 337384 525036 337436 525088
rect 55036 524288 55088 524340
rect 57244 524288 57296 524340
rect 535828 523676 535880 523728
rect 536840 523676 536892 523728
rect 558184 523676 558236 523728
rect 307116 522996 307168 523048
rect 337476 522996 337528 523048
rect 245844 521636 245896 521688
rect 303528 521636 303580 521688
rect 314016 520276 314068 520328
rect 337476 520276 337528 520328
rect 535552 520276 535604 520328
rect 549352 520276 549404 520328
rect 245844 518916 245896 518968
rect 270500 518916 270552 518968
rect 336004 518916 336056 518968
rect 535552 518848 535604 518900
rect 549260 518848 549312 518900
rect 3424 516060 3476 516112
rect 61476 516060 61528 516112
rect 535552 515040 535604 515092
rect 538404 515040 538456 515092
rect 250536 514768 250588 514820
rect 337660 514768 337712 514820
rect 305736 513340 305788 513392
rect 337660 513340 337712 513392
rect 535552 513340 535604 513392
rect 548524 513340 548576 513392
rect 245660 513272 245712 513324
rect 264336 513272 264388 513324
rect 563704 511232 563756 511284
rect 579620 511232 579672 511284
rect 330576 510620 330628 510672
rect 337660 510620 337712 510672
rect 245844 509872 245896 509924
rect 251088 509872 251140 509924
rect 259460 509872 259512 509924
rect 535552 507832 535604 507884
rect 550640 507832 550692 507884
rect 255228 507356 255280 507408
rect 258080 507356 258132 507408
rect 535552 506404 535604 506456
rect 569960 506404 570012 506456
rect 245844 505724 245896 505776
rect 255320 505724 255372 505776
rect 260196 505724 260248 505776
rect 310428 505724 310480 505776
rect 310428 505112 310480 505164
rect 337108 505112 337160 505164
rect 57796 504500 57848 504552
rect 62304 504500 62356 504552
rect 255320 504364 255372 504416
rect 311900 504364 311952 504416
rect 311900 503684 311952 503736
rect 312636 503684 312688 503736
rect 337752 503684 337804 503736
rect 251824 502936 251876 502988
rect 303620 502936 303672 502988
rect 303620 502324 303672 502376
rect 304356 502324 304408 502376
rect 337660 502324 337712 502376
rect 535552 502324 535604 502376
rect 546500 502324 546552 502376
rect 246948 501576 247000 501628
rect 322940 501576 322992 501628
rect 3056 500964 3108 501016
rect 50436 500964 50488 501016
rect 245844 500488 245896 500540
rect 249064 500488 249116 500540
rect 535552 499536 535604 499588
rect 547972 499536 548024 499588
rect 278044 496816 278096 496868
rect 337660 496816 337712 496868
rect 245844 495456 245896 495508
rect 265716 495456 265768 495508
rect 333336 495456 333388 495508
rect 337476 495456 337528 495508
rect 535552 495456 535604 495508
rect 546592 495456 546644 495508
rect 535552 492668 535604 492720
rect 550732 492668 550784 492720
rect 57888 491308 57940 491360
rect 60740 491308 60792 491360
rect 269764 491308 269816 491360
rect 328276 491308 328328 491360
rect 337476 491308 337528 491360
rect 249064 489880 249116 489932
rect 337660 489880 337712 489932
rect 56416 488520 56468 488572
rect 60740 488520 60792 488572
rect 247776 487772 247828 487824
rect 256792 487772 256844 487824
rect 256792 487160 256844 487212
rect 339316 487160 339368 487212
rect 245844 485800 245896 485852
rect 289176 485800 289228 485852
rect 327724 485800 327776 485852
rect 328276 485800 328328 485852
rect 253296 485052 253348 485104
rect 337752 485052 337804 485104
rect 48044 484372 48096 484424
rect 60740 484372 60792 484424
rect 535552 484372 535604 484424
rect 549444 484372 549496 484424
rect 247684 484304 247736 484356
rect 337936 484304 337988 484356
rect 535552 483012 535604 483064
rect 553400 483012 553452 483064
rect 535552 482876 535604 482928
rect 535736 482876 535788 482928
rect 245752 482264 245804 482316
rect 247684 482264 247736 482316
rect 331864 482264 331916 482316
rect 45376 481652 45428 481704
rect 60740 481652 60792 481704
rect 327908 479476 327960 479528
rect 336740 479476 336792 479528
rect 8208 477504 8260 477556
rect 60740 477504 60792 477556
rect 535736 477504 535788 477556
rect 549260 477504 549312 477556
rect 3884 475328 3936 475380
rect 4804 475328 4856 475380
rect 17224 475328 17276 475380
rect 245752 474716 245804 474768
rect 280804 474716 280856 474768
rect 310428 474716 310480 474768
rect 337660 474716 337712 474768
rect 535736 474716 535788 474768
rect 543832 474716 543884 474768
rect 329288 474104 329340 474156
rect 337752 474104 337804 474156
rect 535736 472200 535788 472252
rect 538496 472200 538548 472252
rect 245844 471996 245896 472048
rect 269212 471996 269264 472048
rect 58992 471656 59044 471708
rect 63408 471656 63460 471708
rect 535736 470568 535788 470620
rect 545212 470568 545264 470620
rect 297916 469820 297968 469872
rect 336740 469820 336792 469872
rect 245844 469140 245896 469192
rect 269764 469140 269816 469192
rect 269212 468460 269264 468512
rect 318708 468460 318760 468512
rect 338028 468460 338080 468512
rect 535736 467984 535788 468036
rect 539692 467984 539744 468036
rect 31668 467848 31720 467900
rect 60740 467848 60792 467900
rect 331956 467440 332008 467492
rect 336832 467440 336884 467492
rect 41144 466420 41196 466472
rect 42800 466420 42852 466472
rect 245844 465060 245896 465112
rect 255320 465060 255372 465112
rect 535736 465060 535788 465112
rect 545304 465060 545356 465112
rect 37096 464312 37148 464364
rect 58992 464312 59044 464364
rect 49424 463700 49476 463752
rect 60740 463700 60792 463752
rect 3424 462612 3476 462664
rect 8944 462612 8996 462664
rect 293960 462340 294012 462392
rect 297364 462340 297416 462392
rect 535736 462340 535788 462392
rect 540980 462340 541032 462392
rect 245844 461592 245896 461644
rect 293960 461592 294012 461644
rect 301504 461592 301556 461644
rect 337660 461592 337712 461644
rect 8944 460912 8996 460964
rect 63132 460912 63184 460964
rect 335268 459552 335320 459604
rect 337660 459552 337712 459604
rect 535736 459552 535788 459604
rect 552112 459552 552164 459604
rect 280068 458804 280120 458856
rect 305736 458804 305788 458856
rect 245844 458192 245896 458244
rect 279516 458192 279568 458244
rect 280068 458192 280120 458244
rect 43812 456764 43864 456816
rect 60740 456764 60792 456816
rect 331864 456764 331916 456816
rect 337660 456764 337712 456816
rect 535736 456764 535788 456816
rect 543924 456764 543976 456816
rect 556804 456764 556856 456816
rect 580908 456764 580960 456816
rect 265532 456016 265584 456068
rect 327816 456016 327868 456068
rect 245844 455404 245896 455456
rect 264980 455404 265032 455456
rect 265532 455404 265584 455456
rect 245844 454044 245896 454096
rect 308496 454044 308548 454096
rect 330484 454044 330536 454096
rect 337660 454044 337712 454096
rect 535736 452616 535788 452668
rect 541072 452616 541124 452668
rect 327816 451868 327868 451920
rect 337568 451868 337620 451920
rect 34428 451256 34480 451308
rect 60740 451256 60792 451308
rect 52184 450508 52236 450560
rect 60004 450508 60056 450560
rect 254584 449896 254636 449948
rect 337292 449896 337344 449948
rect 3424 449556 3476 449608
rect 8944 449556 8996 449608
rect 60372 448536 60424 448588
rect 61476 448536 61528 448588
rect 535736 447108 535788 447160
rect 542544 447108 542596 447160
rect 305736 446360 305788 446412
rect 337108 446360 337160 446412
rect 245844 445748 245896 445800
rect 261576 445748 261628 445800
rect 265624 445748 265676 445800
rect 42616 444388 42668 444440
rect 60740 444388 60792 444440
rect 535736 444388 535788 444440
rect 550824 444388 550876 444440
rect 336096 443096 336148 443148
rect 338028 443096 338080 443148
rect 46572 441600 46624 441652
rect 60740 441600 60792 441652
rect 535736 441600 535788 441652
rect 548156 441600 548208 441652
rect 245844 438880 245896 438932
rect 283656 438880 283708 438932
rect 329196 438880 329248 438932
rect 337292 438880 337344 438932
rect 247776 436092 247828 436144
rect 337292 436092 337344 436144
rect 245752 434732 245804 434784
rect 322204 434732 322256 434784
rect 535736 434732 535788 434784
rect 546684 434732 546736 434784
rect 288624 433236 288676 433288
rect 289084 433236 289136 433288
rect 245844 432556 245896 432608
rect 288624 432556 288676 432608
rect 253296 431944 253348 431996
rect 317512 431944 317564 431996
rect 337660 431944 337712 431996
rect 288624 431332 288676 431384
rect 293040 431332 293092 431384
rect 326528 431196 326580 431248
rect 337384 431196 337436 431248
rect 548524 431196 548576 431248
rect 571248 431196 571300 431248
rect 53472 430584 53524 430636
rect 60740 430584 60792 430636
rect 570604 429836 570656 429888
rect 571248 429836 571300 429888
rect 580172 429836 580224 429888
rect 282828 429156 282880 429208
rect 336924 429156 336976 429208
rect 4804 428408 4856 428460
rect 51080 428408 51132 428460
rect 51080 427796 51132 427848
rect 52092 427796 52144 427848
rect 60740 427796 60792 427848
rect 245752 427796 245804 427848
rect 323676 427796 323728 427848
rect 256516 426436 256568 426488
rect 336924 426436 336976 426488
rect 535828 426436 535880 426488
rect 548064 426436 548116 426488
rect 245844 425076 245896 425128
rect 251916 425076 251968 425128
rect 264888 425076 264940 425128
rect 337660 425076 337712 425128
rect 32956 423648 33008 423700
rect 60740 423648 60792 423700
rect 251824 422288 251876 422340
rect 337660 422288 337712 422340
rect 535828 422288 535880 422340
rect 539784 422288 539836 422340
rect 50712 420928 50764 420980
rect 60740 420928 60792 420980
rect 245752 420928 245804 420980
rect 322296 420928 322348 420980
rect 251088 420180 251140 420232
rect 307208 420180 307260 420232
rect 535828 419500 535880 419552
rect 545396 419500 545448 419552
rect 558184 419432 558236 419484
rect 580172 419432 580224 419484
rect 535828 417324 535880 417376
rect 539876 417324 539928 417376
rect 4804 416780 4856 416832
rect 61016 416780 61068 416832
rect 245844 415352 245896 415404
rect 253296 415352 253348 415404
rect 257344 415352 257396 415404
rect 336832 415352 336884 415404
rect 46756 413992 46808 414044
rect 60832 413992 60884 414044
rect 535828 413992 535880 414044
rect 563060 413992 563112 414044
rect 307668 411884 307720 411936
rect 318064 411884 318116 411936
rect 58992 411272 59044 411324
rect 61384 411272 61436 411324
rect 245844 411272 245896 411324
rect 307208 411340 307260 411392
rect 307668 411340 307720 411392
rect 306564 411272 306616 411324
rect 320824 411272 320876 411324
rect 535828 411272 535880 411324
rect 541164 411272 541216 411324
rect 25688 410524 25740 410576
rect 50344 410524 50396 410576
rect 3148 409844 3200 409896
rect 25688 409844 25740 409896
rect 26148 409844 26200 409896
rect 271144 409844 271196 409896
rect 337476 409844 337528 409896
rect 245844 409096 245896 409148
rect 269120 409096 269172 409148
rect 269764 409096 269816 409148
rect 335360 408484 335412 408536
rect 336924 408484 336976 408536
rect 53748 407736 53800 407788
rect 60740 407736 60792 407788
rect 300308 407124 300360 407176
rect 335176 407124 335228 407176
rect 337660 407124 337712 407176
rect 245844 406376 245896 406428
rect 306564 406376 306616 406428
rect 554044 406376 554096 406428
rect 576860 406376 576912 406428
rect 328460 405628 328512 405680
rect 329288 405628 329340 405680
rect 333980 405628 334032 405680
rect 335360 405628 335412 405680
rect 57704 405016 57756 405068
rect 68284 405016 68336 405068
rect 159364 405016 159416 405068
rect 271144 405016 271196 405068
rect 61936 404948 61988 405000
rect 328460 404948 328512 405000
rect 574744 404948 574796 405000
rect 576860 404948 576912 405000
rect 579712 404948 579764 405000
rect 4068 404472 4120 404524
rect 9588 404472 9640 404524
rect 75920 404472 75972 404524
rect 50436 404404 50488 404456
rect 178040 404404 178092 404456
rect 201408 404404 201460 404456
rect 249064 404404 249116 404456
rect 46204 404336 46256 404388
rect 117964 404336 118016 404388
rect 120724 404336 120776 404388
rect 171600 404336 171652 404388
rect 333980 404336 334032 404388
rect 334808 404336 334860 404388
rect 337752 404336 337804 404388
rect 535460 404336 535512 404388
rect 542360 404336 542412 404388
rect 22744 404268 22796 404320
rect 241796 404268 241848 404320
rect 48964 404200 49016 404252
rect 200580 404200 200632 404252
rect 201408 404200 201460 404252
rect 241796 404064 241848 404116
rect 242808 404064 242860 404116
rect 232504 403792 232556 403844
rect 249800 403792 249852 403844
rect 168288 403724 168340 403776
rect 253940 403724 253992 403776
rect 56232 403656 56284 403708
rect 66904 403656 66956 403708
rect 232136 403656 232188 403708
rect 339132 403656 339184 403708
rect 56324 403588 56376 403640
rect 104164 403588 104216 403640
rect 169024 403588 169076 403640
rect 194140 403588 194192 403640
rect 338580 403588 338632 403640
rect 252468 402976 252520 403028
rect 298100 402976 298152 403028
rect 75920 402908 75972 402960
rect 181444 402908 181496 402960
rect 219348 402908 219400 402960
rect 247040 402908 247092 402960
rect 323584 402908 323636 402960
rect 18604 402840 18656 402892
rect 79324 402840 79376 402892
rect 222476 402840 222528 402892
rect 252468 402840 252520 402892
rect 238668 402772 238720 402824
rect 253204 402772 253256 402824
rect 52276 402432 52328 402484
rect 73804 402432 73856 402484
rect 60556 402364 60608 402416
rect 82820 402364 82872 402416
rect 48136 402296 48188 402348
rect 83464 402296 83516 402348
rect 117504 402296 117556 402348
rect 144920 402296 144972 402348
rect 172428 402296 172480 402348
rect 187700 402296 187752 402348
rect 57612 402228 57664 402280
rect 121460 402228 121512 402280
rect 130384 402228 130436 402280
rect 135904 402228 135956 402280
rect 155868 402228 155920 402280
rect 190920 402228 190972 402280
rect 191748 402228 191800 402280
rect 248512 402228 248564 402280
rect 146484 402024 146536 402076
rect 147680 402024 147732 402076
rect 102784 401616 102836 401668
rect 105268 401616 105320 401668
rect 129648 401616 129700 401668
rect 130384 401616 130436 401668
rect 157984 401616 158036 401668
rect 158720 401616 158772 401668
rect 535828 401616 535880 401668
rect 541256 401616 541308 401668
rect 63132 401004 63184 401056
rect 71136 401004 71188 401056
rect 53564 400936 53616 400988
rect 86224 400936 86276 400988
rect 119344 400936 119396 400988
rect 251180 400936 251232 400988
rect 50896 400868 50948 400920
rect 76288 400868 76340 400920
rect 339868 400868 339920 400920
rect 533988 400596 534040 400648
rect 538312 400596 538364 400648
rect 339500 399780 339552 399832
rect 340006 399780 340058 399832
rect 347872 399780 347924 399832
rect 349022 399780 349074 399832
rect 357440 399780 357492 399832
rect 358682 399780 358734 399832
rect 367100 399780 367152 399832
rect 368342 399780 368394 399832
rect 386420 399780 386472 399832
rect 387662 399780 387714 399832
rect 396080 399780 396132 399832
rect 397322 399780 397374 399832
rect 405740 399780 405792 399832
rect 406982 399780 407034 399832
rect 474740 399780 474792 399832
rect 475890 399780 475942 399832
rect 494060 399780 494112 399832
rect 495210 399780 495262 399832
rect 503720 399780 503772 399832
rect 504870 399780 504922 399832
rect 513380 399780 513432 399832
rect 514530 399780 514582 399832
rect 523040 399780 523092 399832
rect 524190 399780 524242 399832
rect 339132 399576 339184 399628
rect 359280 399576 359332 399628
rect 45468 399508 45520 399560
rect 75920 399508 75972 399560
rect 132408 399508 132460 399560
rect 246304 399508 246356 399560
rect 325148 399508 325200 399560
rect 368388 399508 368440 399560
rect 38476 399440 38528 399492
rect 71044 399440 71096 399492
rect 111064 399440 111116 399492
rect 126980 399440 127032 399492
rect 151084 399440 151136 399492
rect 174820 399440 174872 399492
rect 380624 399440 380676 399492
rect 526444 399440 526496 399492
rect 543924 399440 543976 399492
rect 368388 398964 368440 399016
rect 428188 398964 428240 399016
rect 168380 398896 168432 398948
rect 169760 398896 169812 398948
rect 242808 398896 242860 398948
rect 440332 398896 440384 398948
rect 64696 398828 64748 398880
rect 339500 398828 339552 398880
rect 358820 398828 358872 398880
rect 359280 398828 359332 398880
rect 533436 398828 533488 398880
rect 127532 398760 127584 398812
rect 411444 398760 411496 398812
rect 457260 398760 457312 398812
rect 543004 398760 543056 398812
rect 169760 398692 169812 398744
rect 454592 398692 454644 398744
rect 512000 398692 512052 398744
rect 560944 398692 560996 398744
rect 100024 398624 100076 398676
rect 102048 398624 102100 398676
rect 380532 398624 380584 398676
rect 380624 398624 380676 398676
rect 464252 398624 464304 398676
rect 338580 398556 338632 398608
rect 485504 398556 485556 398608
rect 336004 398488 336056 398540
rect 385132 398488 385184 398540
rect 440332 398488 440384 398540
rect 497740 398488 497792 398540
rect 339868 398420 339920 398472
rect 353392 398420 353444 398472
rect 354128 398420 354180 398472
rect 530584 398216 530636 398268
rect 539876 398216 539928 398268
rect 41328 398148 41380 398200
rect 75184 398148 75236 398200
rect 120724 398148 120776 398200
rect 127532 398148 127584 398200
rect 530676 398148 530728 398200
rect 541072 398148 541124 398200
rect 3976 398080 4028 398132
rect 31024 398080 31076 398132
rect 62120 398080 62172 398132
rect 63316 398080 63368 398132
rect 331220 398080 331272 398132
rect 331956 398080 332008 398132
rect 356796 398080 356848 398132
rect 452016 398080 452068 398132
rect 502984 398080 503036 398132
rect 539692 398080 539744 398132
rect 355232 397468 355284 397520
rect 356704 397468 356756 397520
rect 385132 397468 385184 397520
rect 385684 397468 385736 397520
rect 464344 397468 464396 397520
rect 466184 397468 466236 397520
rect 500224 397468 500276 397520
rect 502340 397468 502392 397520
rect 512000 397468 512052 397520
rect 512644 397468 512696 397520
rect 525064 397468 525116 397520
rect 526076 397468 526128 397520
rect 41144 397400 41196 397452
rect 41328 397400 41380 397452
rect 545304 397400 545356 397452
rect 140596 397332 140648 397384
rect 545212 397332 545264 397384
rect 161940 397264 161992 397316
rect 162768 397264 162820 397316
rect 283564 397264 283616 397316
rect 322296 397264 322348 397316
rect 322756 397264 322808 397316
rect 552112 397264 552164 397316
rect 265716 397196 265768 397248
rect 331312 397196 331364 397248
rect 54944 396856 54996 396908
rect 89720 396856 89772 396908
rect 335268 396856 335320 396908
rect 347780 396856 347832 396908
rect 45468 396788 45520 396840
rect 85948 396788 86000 396840
rect 163504 396788 163556 396840
rect 206376 396788 206428 396840
rect 227628 396788 227680 396840
rect 250536 396788 250588 396840
rect 331312 396788 331364 396840
rect 332416 396788 332468 396840
rect 48136 396720 48188 396772
rect 95608 396720 95660 396772
rect 195244 396720 195296 396772
rect 256792 396720 256844 396772
rect 273996 396720 274048 396772
rect 341524 396720 341576 396772
rect 355232 396720 355284 396772
rect 365076 396720 365128 396772
rect 408868 396720 408920 396772
rect 414112 396720 414164 396772
rect 425612 396720 425664 396772
rect 489184 396720 489236 396772
rect 546592 396720 546644 396772
rect 37096 395972 37148 396024
rect 540980 395972 541032 396024
rect 308496 395904 308548 395956
rect 309048 395904 309100 395956
rect 538496 395904 538548 395956
rect 322204 395836 322256 395888
rect 322848 395836 322900 395888
rect 549444 395836 549496 395888
rect 260748 395768 260800 395820
rect 363604 395768 363656 395820
rect 357348 395428 357400 395480
rect 375380 395428 375432 395480
rect 173164 395360 173216 395412
rect 259460 395360 259512 395412
rect 260748 395360 260800 395412
rect 371976 395360 372028 395412
rect 382464 395360 382516 395412
rect 391204 395360 391256 395412
rect 414020 395360 414072 395412
rect 520924 395360 520976 395412
rect 542452 395360 542504 395412
rect 168196 395292 168248 395344
rect 197360 395292 197412 395344
rect 214564 395292 214616 395344
rect 244372 395292 244424 395344
rect 357348 395292 357400 395344
rect 369676 395292 369728 395344
rect 401784 395292 401836 395344
rect 416044 395292 416096 395344
rect 452844 395292 452896 395344
rect 522304 395292 522356 395344
rect 545120 395292 545172 395344
rect 61844 394612 61896 394664
rect 62028 394612 62080 394664
rect 246396 394612 246448 394664
rect 246948 394612 247000 394664
rect 542544 394612 542596 394664
rect 251916 394544 251968 394596
rect 252468 394544 252520 394596
rect 335176 394544 335228 394596
rect 582472 394544 582524 394596
rect 337936 394476 337988 394528
rect 434812 394476 434864 394528
rect 580264 394476 580316 394528
rect 323676 394408 323728 394460
rect 550824 394408 550876 394460
rect 178040 394340 178092 394392
rect 178684 394340 178736 394392
rect 46664 394068 46716 394120
rect 88340 394068 88392 394120
rect 189724 394068 189776 394120
rect 262220 394068 262272 394120
rect 43996 394000 44048 394052
rect 133880 394000 133932 394052
rect 179328 394000 179380 394052
rect 337384 394000 337436 394052
rect 62028 393932 62080 393984
rect 335360 393932 335412 393984
rect 336096 393932 336148 393984
rect 355508 393932 355560 393984
rect 421104 393932 421156 393984
rect 472624 393932 472676 393984
rect 492680 393932 492732 393984
rect 496084 393932 496136 393984
rect 531320 393932 531372 393984
rect 160744 393320 160796 393372
rect 178684 393320 178736 393372
rect 252468 393320 252520 393372
rect 373908 393252 373960 393304
rect 457444 393252 457496 393304
rect 329748 392776 329800 392828
rect 346492 392776 346544 392828
rect 321468 392708 321520 392760
rect 343824 392708 343876 392760
rect 374644 392708 374696 392760
rect 405740 392708 405792 392760
rect 171048 392640 171100 392692
rect 252468 392640 252520 392692
rect 324228 392640 324280 392692
rect 351920 392640 351972 392692
rect 377404 392640 377456 392692
rect 418160 392640 418212 392692
rect 95884 392572 95936 392624
rect 242900 392572 242952 392624
rect 292028 392572 292080 392624
rect 300216 392572 300268 392624
rect 337844 392572 337896 392624
rect 368480 392572 368532 392624
rect 379428 392572 379480 392624
rect 579620 392572 579672 392624
rect 238760 392028 238812 392080
rect 292028 392028 292080 392080
rect 142804 391960 142856 392012
rect 245660 391960 245712 392012
rect 292304 391960 292356 392012
rect 350540 391960 350592 392012
rect 541256 391892 541308 391944
rect 135904 391348 135956 391400
rect 205640 391348 205692 391400
rect 197360 391280 197412 391332
rect 292304 391280 292356 391332
rect 158628 391212 158680 391264
rect 258080 391212 258132 391264
rect 166816 389784 166868 389836
rect 267740 389784 267792 389836
rect 286968 389784 287020 389836
rect 343732 389784 343784 389836
rect 409788 389784 409840 389836
rect 539784 389784 539836 389836
rect 245016 389172 245068 389224
rect 531964 389172 532016 389224
rect 52092 388492 52144 388544
rect 153200 388492 153252 388544
rect 154120 388492 154172 388544
rect 152556 388424 152608 388476
rect 270500 388424 270552 388476
rect 317236 388424 317288 388476
rect 333428 388424 333480 388476
rect 339316 388424 339368 388476
rect 406384 388424 406436 388476
rect 482284 388424 482336 388476
rect 518900 388424 518952 388476
rect 154120 387880 154172 387932
rect 202972 387880 203024 387932
rect 218704 387880 218756 387932
rect 219348 387880 219400 387932
rect 270500 387880 270552 387932
rect 182180 387812 182232 387864
rect 316040 387812 316092 387864
rect 317236 387812 317288 387864
rect 367008 387812 367060 387864
rect 440516 387812 440568 387864
rect 60372 387744 60424 387796
rect 60556 387744 60608 387796
rect 288348 387200 288400 387252
rect 306472 387200 306524 387252
rect 181444 387132 181496 387184
rect 241520 387132 241572 387184
rect 365720 387132 365772 387184
rect 367008 387132 367060 387184
rect 60556 387064 60608 387116
rect 327172 387064 327224 387116
rect 327908 387064 327960 387116
rect 381544 387064 381596 387116
rect 534356 387064 534408 387116
rect 125600 386384 125652 386436
rect 273996 386384 274048 386436
rect 227720 386316 227772 386368
rect 228364 386316 228416 386368
rect 545396 386316 545448 386368
rect 155960 386248 156012 386300
rect 156420 386248 156472 386300
rect 440240 386248 440292 386300
rect 255320 386180 255372 386232
rect 347872 386180 347924 386232
rect 79324 385636 79376 385688
rect 118608 385636 118660 385688
rect 140688 385636 140740 385688
rect 156420 385636 156472 385688
rect 202144 385636 202196 385688
rect 255320 385636 255372 385688
rect 118608 385024 118660 385076
rect 234712 385024 234764 385076
rect 52368 384956 52420 385008
rect 113180 384956 113232 385008
rect 114468 384956 114520 385008
rect 320824 384956 320876 385008
rect 321468 384956 321520 385008
rect 541164 384956 541216 385008
rect 179880 384412 179932 384464
rect 260104 384412 260156 384464
rect 122748 384344 122800 384396
rect 244280 384344 244332 384396
rect 63500 384276 63552 384328
rect 98644 384276 98696 384328
rect 114468 384276 114520 384328
rect 293316 384276 293368 384328
rect 531964 384276 532016 384328
rect 563060 384276 563112 384328
rect 66260 383460 66312 383512
rect 67272 383460 67324 383512
rect 135904 383052 135956 383104
rect 183560 383052 183612 383104
rect 231124 383052 231176 383104
rect 234620 383052 234672 383104
rect 323124 383052 323176 383104
rect 178684 382984 178736 383036
rect 292580 382984 292632 383036
rect 293316 382984 293368 383036
rect 302976 382984 303028 383036
rect 307024 382984 307076 383036
rect 546684 382984 546736 383036
rect 67272 382916 67324 382968
rect 340972 382916 341024 382968
rect 292580 382168 292632 382220
rect 293132 382168 293184 382220
rect 549352 382168 549404 382220
rect 219440 381624 219492 381676
rect 244924 381624 244976 381676
rect 176568 381556 176620 381608
rect 275284 381556 275336 381608
rect 166908 381488 166960 381540
rect 290464 381488 290516 381540
rect 399484 381488 399536 381540
rect 543832 381488 543884 381540
rect 177948 380196 178000 380248
rect 247776 380196 247828 380248
rect 69112 380128 69164 380180
rect 218704 380128 218756 380180
rect 269764 380128 269816 380180
rect 311900 380128 311952 380180
rect 456800 380128 456852 380180
rect 534264 380128 534316 380180
rect 222200 379584 222252 379636
rect 273904 379584 273956 379636
rect 311900 379584 311952 379636
rect 312728 379584 312780 379636
rect 389180 379584 389232 379636
rect 389824 379584 389876 379636
rect 209780 379516 209832 379568
rect 456800 379516 456852 379568
rect 152924 379448 152976 379500
rect 287704 379448 287756 379500
rect 563060 379448 563112 379500
rect 580172 379448 580224 379500
rect 50804 378836 50856 378888
rect 151820 378836 151872 378888
rect 152924 378836 152976 378888
rect 191104 378836 191156 378888
rect 191748 378836 191800 378888
rect 380900 378836 380952 378888
rect 381544 378836 381596 378888
rect 111708 378768 111760 378820
rect 252560 378768 252612 378820
rect 342996 378768 343048 378820
rect 535644 378768 535696 378820
rect 200764 377612 200816 377664
rect 265624 377612 265676 377664
rect 148324 377544 148376 377596
rect 238024 377544 238076 377596
rect 234712 377476 234764 377528
rect 404360 377476 404412 377528
rect 405004 377476 405056 377528
rect 139308 377408 139360 377460
rect 256700 377408 256752 377460
rect 291108 377408 291160 377460
rect 499580 377408 499632 377460
rect 37004 376728 37056 376780
rect 62672 376728 62724 376780
rect 259460 376728 259512 376780
rect 291108 376728 291160 376780
rect 164240 376660 164292 376712
rect 164884 376660 164936 376712
rect 62672 376116 62724 376168
rect 237380 376116 237432 376168
rect 164884 376048 164936 376100
rect 356060 376048 356112 376100
rect 356704 376048 356756 376100
rect 186964 375980 187016 376032
rect 548156 375980 548208 376032
rect 92388 375300 92440 375352
rect 93768 375300 93820 375352
rect 215300 375300 215352 375352
rect 279424 375300 279476 375352
rect 60464 374620 60516 374672
rect 90364 374620 90416 374672
rect 160836 374620 160888 374672
rect 264980 374620 265032 374672
rect 364984 374620 365036 374672
rect 521660 374620 521712 374672
rect 157984 374076 158036 374128
rect 160928 374076 160980 374128
rect 267740 374076 267792 374128
rect 364984 374076 365036 374128
rect 93768 374008 93820 374060
rect 295432 374008 295484 374060
rect 243084 373940 243136 373992
rect 386420 373940 386472 373992
rect 172336 373328 172388 373380
rect 243084 373328 243136 373380
rect 2964 373260 3016 373312
rect 15108 373260 15160 373312
rect 130568 373260 130620 373312
rect 251824 373260 251876 373312
rect 384304 373260 384356 373312
rect 473360 373260 473412 373312
rect 160928 371900 160980 371952
rect 245660 371900 245712 371952
rect 237380 371832 237432 371884
rect 444472 371832 444524 371884
rect 310244 371152 310296 371204
rect 508504 371152 508556 371204
rect 208492 370676 208544 370728
rect 245016 370676 245068 370728
rect 171784 370608 171836 370660
rect 242808 370608 242860 370660
rect 262864 370608 262916 370660
rect 177764 370540 177816 370592
rect 250444 370540 250496 370592
rect 281448 370540 281500 370592
rect 320180 370540 320232 370592
rect 52368 370472 52420 370524
rect 100024 370472 100076 370524
rect 110328 370472 110380 370524
rect 232504 370472 232556 370524
rect 310336 370472 310388 370524
rect 352564 370472 352616 370524
rect 274640 369928 274692 369980
rect 309232 369928 309284 369980
rect 310244 369928 310296 369980
rect 255320 369860 255372 369912
rect 256516 369860 256568 369912
rect 302240 369860 302292 369912
rect 276848 369792 276900 369844
rect 278044 369792 278096 369844
rect 52184 369180 52236 369232
rect 112444 369180 112496 369232
rect 224960 369180 225012 369232
rect 255320 369180 255372 369232
rect 53748 369112 53800 369164
rect 116676 369112 116728 369164
rect 125508 369112 125560 369164
rect 246580 369112 246632 369164
rect 369124 369112 369176 369164
rect 376760 369112 376812 369164
rect 379336 369112 379388 369164
rect 523040 369112 523092 369164
rect 245660 368500 245712 368552
rect 276848 368500 276900 368552
rect 277308 368500 277360 368552
rect 313280 368432 313332 368484
rect 314016 368432 314068 368484
rect 208400 367820 208452 367872
rect 260748 367820 260800 367872
rect 261484 367820 261536 367872
rect 50988 367752 51040 367804
rect 120080 367752 120132 367804
rect 122104 367752 122156 367804
rect 244188 367752 244240 367804
rect 319536 367752 319588 367804
rect 366364 367752 366416 367804
rect 535736 367752 535788 367804
rect 263600 367276 263652 367328
rect 264888 367276 264940 367328
rect 309968 367276 310020 367328
rect 218060 367208 218112 367260
rect 313280 367208 313332 367260
rect 145564 367140 145616 367192
rect 208492 367140 208544 367192
rect 255964 367140 256016 367192
rect 256608 367140 256660 367192
rect 403624 367140 403676 367192
rect 300860 367072 300912 367124
rect 66904 367004 66956 367056
rect 128360 367004 128412 367056
rect 301044 367004 301096 367056
rect 301504 367004 301556 367056
rect 53472 366324 53524 366376
rect 138020 366324 138072 366376
rect 216680 366324 216732 366376
rect 263600 366324 263652 366376
rect 417424 366324 417476 366376
rect 477500 366324 477552 366376
rect 283656 365916 283708 365968
rect 423680 365916 423732 365968
rect 424324 365916 424376 365968
rect 189080 365848 189132 365900
rect 338764 365848 338816 365900
rect 138020 365780 138072 365832
rect 296812 365780 296864 365832
rect 101404 365712 101456 365764
rect 301044 365712 301096 365764
rect 273996 365644 274048 365696
rect 274548 365644 274600 365696
rect 300308 365644 300360 365696
rect 544384 365644 544436 365696
rect 580172 365644 580224 365696
rect 179236 365100 179288 365152
rect 264244 365100 264296 365152
rect 314016 365168 314068 365220
rect 300768 365100 300820 365152
rect 372620 365100 372672 365152
rect 173716 365032 173768 365084
rect 42616 364964 42668 365016
rect 96620 364964 96672 365016
rect 126244 364964 126296 365016
rect 245752 364964 245804 365016
rect 363604 365032 363656 365084
rect 440332 365032 440384 365084
rect 279516 364964 279568 365016
rect 418804 364964 418856 365016
rect 96620 364420 96672 364472
rect 300952 364420 301004 364472
rect 83464 364352 83516 364404
rect 307852 364352 307904 364404
rect 273904 363808 273956 363860
rect 298192 363808 298244 363860
rect 277308 363740 277360 363792
rect 347044 363740 347096 363792
rect 228824 363672 228876 363724
rect 336648 363672 336700 363724
rect 41236 363604 41288 363656
rect 305000 363604 305052 363656
rect 389824 363604 389876 363656
rect 431960 363604 432012 363656
rect 432052 363604 432104 363656
rect 452660 363604 452712 363656
rect 305000 363400 305052 363452
rect 305736 363400 305788 363452
rect 144184 362992 144236 363044
rect 212540 362992 212592 363044
rect 245752 362992 245804 363044
rect 246948 362992 247000 363044
rect 315396 362992 315448 363044
rect 162308 362924 162360 362976
rect 162768 362924 162820 362976
rect 294052 362924 294104 362976
rect 336648 362924 336700 362976
rect 340880 362924 340932 362976
rect 212540 362312 212592 362364
rect 256700 362312 256752 362364
rect 140044 362244 140096 362296
rect 245752 362244 245804 362296
rect 95148 362176 95200 362228
rect 117964 362176 118016 362228
rect 122656 362176 122708 362228
rect 242992 362176 243044 362228
rect 258908 362176 258960 362228
rect 289728 362176 289780 362228
rect 336740 362176 336792 362228
rect 340144 361700 340196 361752
rect 413284 361700 413336 361752
rect 153108 361632 153160 361684
rect 201592 361632 201644 361684
rect 202144 361632 202196 361684
rect 227352 361632 227404 361684
rect 227628 361632 227680 361684
rect 342260 361632 342312 361684
rect 175096 361564 175148 361616
rect 359464 361564 359516 361616
rect 287704 360816 287756 360868
rect 316132 360816 316184 360868
rect 250536 360340 250588 360392
rect 251088 360340 251140 360392
rect 349436 360340 349488 360392
rect 113180 360272 113232 360324
rect 317512 360272 317564 360324
rect 70400 360204 70452 360256
rect 71136 360204 71188 360256
rect 291200 360204 291252 360256
rect 243912 359660 243964 359712
rect 277400 359660 277452 359712
rect 177856 359592 177908 359644
rect 254584 359592 254636 359644
rect 166632 359524 166684 359576
rect 248420 359524 248472 359576
rect 170956 359456 171008 359508
rect 255964 359456 256016 359508
rect 375104 359456 375156 359508
rect 391940 359456 391992 359508
rect 393964 359456 394016 359508
rect 489920 359456 489972 359508
rect 68284 358912 68336 358964
rect 193404 358912 193456 358964
rect 146944 358844 146996 358896
rect 276664 358844 276716 358896
rect 277124 358844 277176 358896
rect 349804 358912 349856 358964
rect 279424 358844 279476 358896
rect 454040 358844 454092 358896
rect 166264 358776 166316 358828
rect 166816 358776 166868 358828
rect 445024 358776 445076 358828
rect 2780 358436 2832 358488
rect 4804 358436 4856 358488
rect 290464 358096 290516 358148
rect 298008 358096 298060 358148
rect 175924 357756 175976 357808
rect 195244 357756 195296 357808
rect 212356 357756 212408 357808
rect 214564 357756 214616 357808
rect 285956 357756 286008 357808
rect 286968 357756 287020 357808
rect 306380 357756 306432 357808
rect 162124 357688 162176 357740
rect 247684 357688 247736 357740
rect 248144 357688 248196 357740
rect 262864 357688 262916 357740
rect 265348 357688 265400 357740
rect 265624 357688 265676 357740
rect 300308 357688 300360 357740
rect 170496 357620 170548 357672
rect 283656 357620 283708 357672
rect 287336 357620 287388 357672
rect 91744 357552 91796 357604
rect 212448 357552 212500 357604
rect 231124 357552 231176 357604
rect 293224 357552 293276 357604
rect 169116 357484 169168 357536
rect 202880 357484 202932 357536
rect 307760 357484 307812 357536
rect 43996 357416 44048 357468
rect 243912 357416 243964 357468
rect 251088 357416 251140 357468
rect 253940 357416 253992 357468
rect 256700 357416 256752 357468
rect 304540 357416 304592 357468
rect 212448 357348 212500 357400
rect 261576 357348 261628 357400
rect 262128 357348 262180 357400
rect 273720 357348 273772 357400
rect 274548 357348 274600 357400
rect 117964 356736 118016 356788
rect 212356 356736 212408 356788
rect 262128 356736 262180 356788
rect 297456 356736 297508 356788
rect 109684 356668 109736 356720
rect 251088 356668 251140 356720
rect 262864 356668 262916 356720
rect 429844 356668 429896 356720
rect 171140 356260 171192 356312
rect 199660 356260 199712 356312
rect 262772 356260 262824 356312
rect 351184 356260 351236 356312
rect 154488 356192 154540 356244
rect 186780 356192 186832 356244
rect 193404 356192 193456 356244
rect 297640 356192 297692 356244
rect 134616 356124 134668 356176
rect 266360 356124 266412 356176
rect 266820 356124 266872 356176
rect 270408 356124 270460 356176
rect 273720 356124 273772 356176
rect 298744 356124 298796 356176
rect 170588 356056 170640 356108
rect 326436 356056 326488 356108
rect 270408 355988 270460 356040
rect 417424 355988 417476 356040
rect 164148 355444 164200 355496
rect 191104 355444 191156 355496
rect 49424 355376 49476 355428
rect 167000 355376 167052 355428
rect 173808 355376 173860 355428
rect 189724 355376 189776 355428
rect 254400 355376 254452 355428
rect 425704 355376 425756 355428
rect 112536 355308 112588 355360
rect 289176 355308 289228 355360
rect 295524 355308 295576 355360
rect 424324 355308 424376 355360
rect 450544 355308 450596 355360
rect 292304 354900 292356 354952
rect 292580 354900 292632 354952
rect 179420 354832 179472 354884
rect 219440 354832 219492 354884
rect 220452 354832 220504 354884
rect 301504 354832 301556 354884
rect 174544 354764 174596 354816
rect 279056 354764 279108 354816
rect 284024 354764 284076 354816
rect 302884 354764 302936 354816
rect 167000 354696 167052 354748
rect 209872 354696 209924 354748
rect 271144 354696 271196 354748
rect 385040 354696 385092 354748
rect 292488 354492 292540 354544
rect 293316 354492 293368 354544
rect 295432 354424 295484 354476
rect 295616 354424 295668 354476
rect 53748 353948 53800 354000
rect 179420 353948 179472 354000
rect 295432 353268 295484 353320
rect 346308 353268 346360 353320
rect 43904 353200 43956 353252
rect 171140 353200 171192 353252
rect 54944 352520 54996 352572
rect 68284 352520 68336 352572
rect 295432 352520 295484 352572
rect 297916 352520 297968 352572
rect 346308 352520 346360 352572
rect 442172 352520 442224 352572
rect 345664 352452 345716 352504
rect 437388 351908 437440 351960
rect 580172 351908 580224 351960
rect 442172 351840 442224 351892
rect 442908 351840 442960 351892
rect 548064 351840 548116 351892
rect 293224 351160 293276 351212
rect 438860 351160 438912 351212
rect 295432 350480 295484 350532
rect 302332 350480 302384 350532
rect 302976 350480 303028 350532
rect 438860 350480 438912 350532
rect 440148 350480 440200 350532
rect 547880 350480 547932 350532
rect 45284 349800 45336 349852
rect 171784 349800 171836 349852
rect 302332 349800 302384 349852
rect 325148 349800 325200 349852
rect 63224 348372 63276 348424
rect 133144 348372 133196 348424
rect 429108 348372 429160 348424
rect 574744 348372 574796 348424
rect 132592 347760 132644 347812
rect 133144 347760 133196 347812
rect 176660 347760 176712 347812
rect 49424 347012 49476 347064
rect 179236 347012 179288 347064
rect 295432 347012 295484 347064
rect 295800 347012 295852 347064
rect 300768 347012 300820 347064
rect 311256 347012 311308 347064
rect 355324 347012 355376 347064
rect 437480 347012 437532 347064
rect 3332 345652 3384 345704
rect 44824 345652 44876 345704
rect 118516 345652 118568 345704
rect 130476 345652 130528 345704
rect 173716 345652 173768 345704
rect 176660 345652 176712 345704
rect 295616 345652 295668 345704
rect 318616 345652 318668 345704
rect 534172 345652 534224 345704
rect 118516 344972 118568 345024
rect 178684 344972 178736 345024
rect 295432 342864 295484 342916
rect 296812 342864 296864 342916
rect 299940 342864 299992 342916
rect 359464 342184 359516 342236
rect 502984 342184 503036 342236
rect 359464 341572 359516 341624
rect 360016 341572 360068 341624
rect 78588 341504 78640 341556
rect 132500 341504 132552 341556
rect 175004 340824 175056 340876
rect 176660 340824 176712 340876
rect 295432 340824 295484 340876
rect 311808 340824 311860 340876
rect 68652 340144 68704 340196
rect 175924 340144 175976 340196
rect 311808 340144 311860 340196
rect 344284 340144 344336 340196
rect 362224 340144 362276 340196
rect 528560 340144 528612 340196
rect 295432 339396 295484 339448
rect 301044 339396 301096 339448
rect 301320 339396 301372 339448
rect 301320 338784 301372 338836
rect 325240 338784 325292 338836
rect 295984 338716 296036 338768
rect 538404 338716 538456 338768
rect 175096 338104 175148 338156
rect 176660 338104 176712 338156
rect 49516 337356 49568 337408
rect 122932 337356 122984 337408
rect 175004 337356 175056 337408
rect 299940 335996 299992 336048
rect 401600 335996 401652 336048
rect 371884 334636 371936 334688
rect 396080 334636 396132 334688
rect 477960 334636 478012 334688
rect 552020 334636 552072 334688
rect 175188 334568 175240 334620
rect 176660 334568 176712 334620
rect 295708 334568 295760 334620
rect 365260 334568 365312 334620
rect 379244 334568 379296 334620
rect 512644 334568 512696 334620
rect 401600 333956 401652 334008
rect 477500 333956 477552 334008
rect 477960 333956 478012 334008
rect 169760 333888 169812 333940
rect 170956 333888 171008 333940
rect 176660 333888 176712 333940
rect 130660 333276 130712 333328
rect 169760 333276 169812 333328
rect 295432 333276 295484 333328
rect 353944 333276 353996 333328
rect 66904 333208 66956 333260
rect 149060 333208 149112 333260
rect 304448 333208 304500 333260
rect 513380 333208 513432 333260
rect 106924 331848 106976 331900
rect 175188 331848 175240 331900
rect 355416 331848 355468 331900
rect 441620 331848 441672 331900
rect 293868 331236 293920 331288
rect 337384 331236 337436 331288
rect 295432 330488 295484 330540
rect 300952 330488 301004 330540
rect 301320 330488 301372 330540
rect 58992 329060 59044 329112
rect 74632 329060 74684 329112
rect 75276 329060 75328 329112
rect 301320 329060 301372 329112
rect 440240 329060 440292 329112
rect 75276 328448 75328 328500
rect 134524 328448 134576 328500
rect 440240 328380 440292 328432
rect 440884 328380 440936 328432
rect 543740 328380 543792 328432
rect 295524 327700 295576 327752
rect 310428 327700 310480 327752
rect 293132 327020 293184 327072
rect 310336 327020 310388 327072
rect 310336 326408 310388 326460
rect 348424 326408 348476 326460
rect 296628 326340 296680 326392
rect 537116 326340 537168 326392
rect 173256 325660 173308 325712
rect 176660 325660 176712 325712
rect 310336 324912 310388 324964
rect 391204 324912 391256 324964
rect 337936 323552 337988 323604
rect 458180 323552 458232 323604
rect 294328 322940 294380 322992
rect 337936 322940 337988 322992
rect 81532 322872 81584 322924
rect 82820 322872 82872 322924
rect 146300 322872 146352 322924
rect 300216 322192 300268 322244
rect 369860 322192 369912 322244
rect 370504 322192 370556 322244
rect 434720 322192 434772 322244
rect 438768 322192 438820 322244
rect 509240 322192 509292 322244
rect 413284 321648 413336 321700
rect 420184 321648 420236 321700
rect 175188 321580 175240 321632
rect 177580 321580 177632 321632
rect 177764 321580 177816 321632
rect 295340 321512 295392 321564
rect 305736 321512 305788 321564
rect 306288 321512 306340 321564
rect 310428 321512 310480 321564
rect 393964 321512 394016 321564
rect 305736 320832 305788 320884
rect 319628 320832 319680 320884
rect 359464 320832 359516 320884
rect 448520 320832 448572 320884
rect 3148 320084 3200 320136
rect 59268 320084 59320 320136
rect 367744 319472 367796 319524
rect 394700 319472 394752 319524
rect 59268 319404 59320 319456
rect 87604 319404 87656 319456
rect 313372 319404 313424 319456
rect 314568 319404 314620 319456
rect 325056 319404 325108 319456
rect 379520 319404 379572 319456
rect 483020 319404 483072 319456
rect 295340 318792 295392 318844
rect 313372 318792 313424 318844
rect 447140 318792 447192 318844
rect 466460 318792 466512 318844
rect 81440 318724 81492 318776
rect 106280 318724 106332 318776
rect 106924 318724 106976 318776
rect 33048 318044 33100 318096
rect 136732 318044 136784 318096
rect 147588 318044 147640 318096
rect 173256 318044 173308 318096
rect 379152 318044 379204 318096
rect 447140 318044 447192 318096
rect 136732 317432 136784 317484
rect 147588 317432 147640 317484
rect 177948 317364 178000 317416
rect 179144 317364 179196 317416
rect 345848 316820 345900 316872
rect 377404 316820 377456 316872
rect 304540 316752 304592 316804
rect 362960 316752 363012 316804
rect 59176 316684 59228 316736
rect 105544 316684 105596 316736
rect 295340 316684 295392 316736
rect 299296 316684 299348 316736
rect 338028 316684 338080 316736
rect 443092 316684 443144 316736
rect 362960 316004 363012 316056
rect 364248 316004 364300 316056
rect 415584 316004 415636 316056
rect 299296 315936 299348 315988
rect 305000 315936 305052 315988
rect 49608 315256 49660 315308
rect 59268 315256 59320 315308
rect 87604 315256 87656 315308
rect 116768 315256 116820 315308
rect 305000 315256 305052 315308
rect 373264 315256 373316 315308
rect 452568 315256 452620 315308
rect 556804 315256 556856 315308
rect 59268 314644 59320 314696
rect 157248 314644 157300 314696
rect 179328 314644 179380 314696
rect 295340 314576 295392 314628
rect 317604 314576 317656 314628
rect 318524 314576 318576 314628
rect 320824 314576 320876 314628
rect 386512 314576 386564 314628
rect 451280 314644 451332 314696
rect 452568 314644 452620 314696
rect 34428 313896 34480 313948
rect 124220 313896 124272 313948
rect 296076 313896 296128 313948
rect 306472 313896 306524 313948
rect 318524 313896 318576 313948
rect 386328 313896 386380 313948
rect 385684 313420 385736 313472
rect 389180 313420 389232 313472
rect 57796 313216 57848 313268
rect 109040 313216 109092 313268
rect 109040 312604 109092 312656
rect 109684 312604 109736 312656
rect 420184 312604 420236 312656
rect 440976 312604 441028 312656
rect 170680 312536 170732 312588
rect 171048 312536 171100 312588
rect 176660 312536 176712 312588
rect 295340 312536 295392 312588
rect 305000 312536 305052 312588
rect 360844 312536 360896 312588
rect 430580 312536 430632 312588
rect 450544 312536 450596 312588
rect 458180 312536 458232 312588
rect 305000 311856 305052 311908
rect 372620 311856 372672 311908
rect 458180 311856 458232 311908
rect 579988 311856 580040 311908
rect 457444 311788 457496 311840
rect 460940 311788 460992 311840
rect 79324 311176 79376 311228
rect 157984 311176 158036 311228
rect 43812 311108 43864 311160
rect 132500 311108 132552 311160
rect 85580 310972 85632 311024
rect 86224 310972 86276 311024
rect 86224 310496 86276 310548
rect 170404 310496 170456 310548
rect 295340 310428 295392 310480
rect 307852 310428 307904 310480
rect 308956 310428 309008 310480
rect 173348 310224 173400 310276
rect 173808 310224 173860 310276
rect 176660 310224 176712 310276
rect 386328 309884 386380 309936
rect 395344 309884 395396 309936
rect 308956 309816 309008 309868
rect 360292 309816 360344 309868
rect 372620 309816 372672 309868
rect 391204 309816 391256 309868
rect 41236 309748 41288 309800
rect 68284 309748 68336 309800
rect 326436 309748 326488 309800
rect 419540 309748 419592 309800
rect 360292 309136 360344 309188
rect 361488 309136 361540 309188
rect 384304 309136 384356 309188
rect 419540 309068 419592 309120
rect 420184 309068 420236 309120
rect 436928 309068 436980 309120
rect 437388 309068 437440 309120
rect 39764 308456 39816 308508
rect 69020 308456 69072 308508
rect 93768 308456 93820 308508
rect 114560 308456 114612 308508
rect 436928 308456 436980 308508
rect 465080 308456 465132 308508
rect 48044 308388 48096 308440
rect 131856 308388 131908 308440
rect 458364 308388 458416 308440
rect 575480 308388 575532 308440
rect 73068 307776 73120 307828
rect 75920 307776 75972 307828
rect 295340 307776 295392 307828
rect 303620 307776 303672 307828
rect 399484 307776 399536 307828
rect 434168 307776 434220 307828
rect 458364 307776 458416 307828
rect 88432 307300 88484 307352
rect 89720 307300 89772 307352
rect 379612 307164 379664 307216
rect 386420 307164 386472 307216
rect 377496 307096 377548 307148
rect 398840 307096 398892 307148
rect 300308 307028 300360 307080
rect 441712 307028 441764 307080
rect 89720 306960 89772 307012
rect 90364 306960 90416 307012
rect 80060 306688 80112 306740
rect 83464 306688 83516 306740
rect 113272 306484 113324 306536
rect 113824 306484 113876 306536
rect 159456 306484 159508 306536
rect 102140 306416 102192 306468
rect 160928 306416 160980 306468
rect 90364 306348 90416 306400
rect 152464 306348 152516 306400
rect 391204 306348 391256 306400
rect 469220 306348 469272 306400
rect 172336 306076 172388 306128
rect 176660 306076 176712 306128
rect 76656 305668 76708 305720
rect 112536 305668 112588 305720
rect 121368 305668 121420 305720
rect 172336 305668 172388 305720
rect 45376 305600 45428 305652
rect 127072 305600 127124 305652
rect 410524 305600 410576 305652
rect 448612 305600 448664 305652
rect 294052 305328 294104 305380
rect 295340 305328 295392 305380
rect 88340 305056 88392 305108
rect 88984 305056 89036 305108
rect 136088 305056 136140 305108
rect 405004 305056 405056 305108
rect 455420 305056 455472 305108
rect 3240 304988 3292 305040
rect 120264 304988 120316 305040
rect 121368 304988 121420 305040
rect 409604 304988 409656 305040
rect 463700 304988 463752 305040
rect 134524 304376 134576 304428
rect 173256 304376 173308 304428
rect 114744 304308 114796 304360
rect 173348 304308 173400 304360
rect 104992 304240 105044 304292
rect 167736 304240 167788 304292
rect 295340 304240 295392 304292
rect 441620 304240 441672 304292
rect 103520 303900 103572 303952
rect 104992 303900 105044 303952
rect 429844 303900 429896 303952
rect 430304 303900 430356 303952
rect 447140 303900 447192 303952
rect 98552 303832 98604 303884
rect 98736 303832 98788 303884
rect 129004 303832 129056 303884
rect 406384 303832 406436 303884
rect 443000 303832 443052 303884
rect 81440 303764 81492 303816
rect 138664 303764 138716 303816
rect 417608 303764 417660 303816
rect 458180 303764 458232 303816
rect 70492 303696 70544 303748
rect 71044 303696 71096 303748
rect 153844 303696 153896 303748
rect 373724 303696 373776 303748
rect 380900 303696 380952 303748
rect 399484 303696 399536 303748
rect 444380 303696 444432 303748
rect 22744 303628 22796 303680
rect 117872 303628 117924 303680
rect 362868 303628 362920 303680
rect 389180 303628 389232 303680
rect 395344 303628 395396 303680
rect 471980 303628 472032 303680
rect 295340 303560 295392 303612
rect 300860 303560 300912 303612
rect 398104 303560 398156 303612
rect 405004 303560 405056 303612
rect 111800 303016 111852 303068
rect 128360 303016 128412 303068
rect 46848 302948 46900 303000
rect 68744 302948 68796 303000
rect 102140 302948 102192 303000
rect 106188 302948 106240 303000
rect 122840 302948 122892 303000
rect 300860 302948 300912 303000
rect 356796 302948 356848 303000
rect 35716 302880 35768 302932
rect 126428 302880 126480 302932
rect 297548 302880 297600 302932
rect 304356 302880 304408 302932
rect 374736 302880 374788 302932
rect 403624 302540 403676 302592
rect 459652 302540 459704 302592
rect 425888 302472 425940 302524
rect 446404 302472 446456 302524
rect 428372 302404 428424 302456
rect 429108 302404 429160 302456
rect 451372 302404 451424 302456
rect 360108 302336 360160 302388
rect 385040 302336 385092 302388
rect 385776 302336 385828 302388
rect 440148 302336 440200 302388
rect 470692 302336 470744 302388
rect 88432 302268 88484 302320
rect 157984 302268 158036 302320
rect 376208 302268 376260 302320
rect 423864 302268 423916 302320
rect 456800 302268 456852 302320
rect 90272 302200 90324 302252
rect 162216 302200 162268 302252
rect 374736 302200 374788 302252
rect 375288 302200 375340 302252
rect 407672 302200 407724 302252
rect 103612 301588 103664 301640
rect 130660 301588 130712 301640
rect 107660 301520 107712 301572
rect 139308 301520 139360 301572
rect 144276 301520 144328 301572
rect 129188 301452 129240 301504
rect 162308 301452 162360 301504
rect 418804 301452 418856 301504
rect 448520 301452 448572 301504
rect 74540 300976 74592 301028
rect 149796 300976 149848 301028
rect 393596 300976 393648 301028
rect 393964 300976 394016 301028
rect 446496 300976 446548 301028
rect 79232 300908 79284 300960
rect 164976 300908 165028 300960
rect 376116 300908 376168 300960
rect 409604 300908 409656 300960
rect 412364 300908 412416 300960
rect 484400 300908 484452 300960
rect 59084 300840 59136 300892
rect 295340 300840 295392 300892
rect 300308 300840 300360 300892
rect 301596 300840 301648 300892
rect 436008 300840 436060 300892
rect 438492 300840 438544 300892
rect 449900 300840 449952 300892
rect 155776 300772 155828 300824
rect 159364 300772 159416 300824
rect 421012 300772 421064 300824
rect 421840 300772 421892 300824
rect 116584 300228 116636 300280
rect 129740 300228 129792 300280
rect 91100 300160 91152 300212
rect 170680 300160 170732 300212
rect 39856 300092 39908 300144
rect 127164 300092 127216 300144
rect 101496 299616 101548 299668
rect 137284 299616 137336 299668
rect 416504 299616 416556 299668
rect 438860 299616 438912 299668
rect 86960 299548 87012 299600
rect 142804 299548 142856 299600
rect 358084 299548 358136 299600
rect 414020 299548 414072 299600
rect 422024 299548 422076 299600
rect 454132 299548 454184 299600
rect 67456 299480 67508 299532
rect 152556 299480 152608 299532
rect 293224 299480 293276 299532
rect 411812 299480 411864 299532
rect 414480 299480 414532 299532
rect 476212 299480 476264 299532
rect 105544 299412 105596 299464
rect 106096 299412 106148 299464
rect 167092 299412 167144 299464
rect 168196 299412 168248 299464
rect 176660 299412 176712 299464
rect 438860 299412 438912 299464
rect 553492 299412 553544 299464
rect 579620 299412 579672 299464
rect 108672 299344 108724 299396
rect 111800 299344 111852 299396
rect 53564 298732 53616 298784
rect 167092 298732 167144 298784
rect 112904 298392 112956 298444
rect 149704 298392 149756 298444
rect 106096 298324 106148 298376
rect 145656 298324 145708 298376
rect 84200 298256 84252 298308
rect 141516 298256 141568 298308
rect 68468 298188 68520 298240
rect 160836 298188 160888 298240
rect 72976 298120 73028 298172
rect 170588 298120 170640 298172
rect 52460 298052 52512 298104
rect 53656 298052 53708 298104
rect 101404 298052 101456 298104
rect 44824 297372 44876 297424
rect 52460 297372 52512 297424
rect 314016 297372 314068 297424
rect 369768 297372 369820 297424
rect 102876 297032 102928 297084
rect 134524 297032 134576 297084
rect 93216 296964 93268 297016
rect 124864 296964 124916 297016
rect 83556 296896 83608 296948
rect 144368 296896 144420 296948
rect 172336 296896 172388 296948
rect 176660 296896 176712 296948
rect 442816 296896 442868 296948
rect 444564 296896 444616 296948
rect 93860 296828 93912 296880
rect 159364 296828 159416 296880
rect 95148 296760 95200 296812
rect 102784 296760 102836 296812
rect 172336 296760 172388 296812
rect 50712 296692 50764 296744
rect 158168 296692 158220 296744
rect 369768 296692 369820 296744
rect 376944 296692 376996 296744
rect 60464 296012 60516 296064
rect 84844 296012 84896 296064
rect 67364 295944 67416 295996
rect 169116 295944 169168 295996
rect 113824 295604 113876 295656
rect 123576 295604 123628 295656
rect 118516 295536 118568 295588
rect 119620 295536 119672 295588
rect 82912 295468 82964 295520
rect 134708 295468 134760 295520
rect 100944 295400 100996 295452
rect 155224 295400 155276 295452
rect 69020 295332 69072 295384
rect 71780 295332 71832 295384
rect 94504 295332 94556 295384
rect 95056 295332 95108 295384
rect 148508 295332 148560 295384
rect 295340 295332 295392 295384
rect 309876 295332 309928 295384
rect 310336 295332 310388 295384
rect 46572 295264 46624 295316
rect 72976 295264 73028 295316
rect 73896 295264 73948 295316
rect 297640 295264 297692 295316
rect 379152 295264 379204 295316
rect 310336 295196 310388 295248
rect 319444 295196 319496 295248
rect 73252 294924 73304 294976
rect 74632 294924 74684 294976
rect 73804 294788 73856 294840
rect 84844 294788 84896 294840
rect 70032 294652 70084 294704
rect 101496 294652 101548 294704
rect 9588 294584 9640 294636
rect 72608 294584 72660 294636
rect 95792 294584 95844 294636
rect 168288 294584 168340 294636
rect 442816 294584 442868 294636
rect 452752 294584 452804 294636
rect 75184 294244 75236 294296
rect 141424 294244 141476 294296
rect 85488 294176 85540 294228
rect 91744 294176 91796 294228
rect 91928 294176 91980 294228
rect 133144 294176 133196 294228
rect 62764 294108 62816 294160
rect 96620 294108 96672 294160
rect 102232 294108 102284 294160
rect 151176 294108 151228 294160
rect 78404 294040 78456 294092
rect 129096 294040 129148 294092
rect 70400 293972 70452 294024
rect 71044 293972 71096 294024
rect 76472 293972 76524 294024
rect 77944 293972 77996 294024
rect 81440 293972 81492 294024
rect 81900 293972 81952 294024
rect 88340 293972 88392 294024
rect 89076 293972 89128 294024
rect 103612 293972 103664 294024
rect 104532 293972 104584 294024
rect 109040 293972 109092 294024
rect 109684 293972 109736 294024
rect 111892 293972 111944 294024
rect 114560 293972 114612 294024
rect 115388 293972 115440 294024
rect 120356 293972 120408 294024
rect 173348 293972 173400 294024
rect 176660 293972 176712 294024
rect 79048 293496 79100 293548
rect 79324 293496 79376 293548
rect 98368 293496 98420 293548
rect 98644 293496 98696 293548
rect 296720 293224 296772 293276
rect 307024 293224 307076 293276
rect 116400 292884 116452 292936
rect 116768 292884 116820 292936
rect 123668 292884 123720 292936
rect 99656 292816 99708 292868
rect 131764 292816 131816 292868
rect 58716 292748 58768 292800
rect 92572 292748 92624 292800
rect 105452 292748 105504 292800
rect 106188 292748 106240 292800
rect 152648 292748 152700 292800
rect 88064 292680 88116 292732
rect 136180 292680 136232 292732
rect 57244 292612 57296 292664
rect 79048 292612 79100 292664
rect 80980 292612 81032 292664
rect 138756 292612 138808 292664
rect 4068 292544 4120 292596
rect 95976 292544 96028 292596
rect 98368 292544 98420 292596
rect 178684 292544 178736 292596
rect 295340 292476 295392 292528
rect 305092 292476 305144 292528
rect 305552 292476 305604 292528
rect 86408 291864 86460 291916
rect 3240 291796 3292 291848
rect 17224 291796 17276 291848
rect 68468 291796 68520 291848
rect 68652 291796 68704 291848
rect 110788 291864 110840 291916
rect 122564 291864 122616 291916
rect 122748 291864 122800 291916
rect 120356 291796 120408 291848
rect 141608 291796 141660 291848
rect 151360 291252 151412 291304
rect 147036 291184 147088 291236
rect 163688 291116 163740 291168
rect 164148 291116 164200 291168
rect 294052 291116 294104 291168
rect 343732 291116 343784 291168
rect 13084 290436 13136 290488
rect 39948 290436 40000 290488
rect 49608 290436 49660 290488
rect 126336 290436 126388 290488
rect 148324 290436 148376 290488
rect 163688 290436 163740 290488
rect 176660 290436 176712 290488
rect 343732 290436 343784 290488
rect 365168 290436 365220 290488
rect 373264 290436 373316 290488
rect 373816 290436 373868 290488
rect 376944 290436 376996 290488
rect 49608 289892 49660 289944
rect 67732 289892 67784 289944
rect 121552 289892 121604 289944
rect 140136 289892 140188 289944
rect 43812 289824 43864 289876
rect 67640 289824 67692 289876
rect 121644 289824 121696 289876
rect 167644 289824 167696 289876
rect 295340 289824 295392 289876
rect 440332 289824 440384 289876
rect 449992 289824 450044 289876
rect 121552 289756 121604 289808
rect 145564 289756 145616 289808
rect 306288 289756 306340 289808
rect 307760 289756 307812 289808
rect 377956 289756 378008 289808
rect 378784 289756 378836 289808
rect 121644 289688 121696 289740
rect 133880 289688 133932 289740
rect 135168 289688 135220 289740
rect 300308 289688 300360 289740
rect 311900 289688 311952 289740
rect 43904 289076 43956 289128
rect 64880 289076 64932 289128
rect 67732 289076 67784 289128
rect 311900 289076 311952 289128
rect 312544 289076 312596 289128
rect 367008 289076 367060 289128
rect 64604 288396 64656 288448
rect 67640 288396 67692 288448
rect 367008 288396 367060 288448
rect 376944 288396 376996 288448
rect 121552 288328 121604 288380
rect 174544 288328 174596 288380
rect 170588 288260 170640 288312
rect 176660 288260 176712 288312
rect 48044 287036 48096 287088
rect 67640 287036 67692 287088
rect 296168 287036 296220 287088
rect 342904 287036 342956 287088
rect 441528 287036 441580 287088
rect 447784 287036 447836 287088
rect 138848 286356 138900 286408
rect 142160 286356 142212 286408
rect 157156 286356 157208 286408
rect 173348 286356 173400 286408
rect 121736 286288 121788 286340
rect 124312 286288 124364 286340
rect 163596 286288 163648 286340
rect 325240 286288 325292 286340
rect 369860 286288 369912 286340
rect 50988 285676 51040 285728
rect 67732 285676 67784 285728
rect 369860 285676 369912 285728
rect 371148 285676 371200 285728
rect 376944 285676 376996 285728
rect 445024 285676 445076 285728
rect 480352 285676 480404 285728
rect 121460 285608 121512 285660
rect 125600 285608 125652 285660
rect 442172 285608 442224 285660
rect 122472 284928 122524 284980
rect 169116 284928 169168 284980
rect 41236 284316 41288 284368
rect 67640 284316 67692 284368
rect 160836 284316 160888 284368
rect 162768 284316 162820 284368
rect 174636 284316 174688 284368
rect 50712 284248 50764 284300
rect 67732 284248 67784 284300
rect 122748 284248 122800 284300
rect 124220 284248 124272 284300
rect 158628 284248 158680 284300
rect 176660 284248 176712 284300
rect 121460 283568 121512 283620
rect 173164 283568 173216 283620
rect 173348 283568 173400 283620
rect 298744 283568 298796 283620
rect 377312 283568 377364 283620
rect 377864 283568 377916 283620
rect 294788 282888 294840 282940
rect 310520 282888 310572 282940
rect 376024 282888 376076 282940
rect 166264 282820 166316 282872
rect 176660 282820 176712 282872
rect 442724 281800 442776 281852
rect 450084 281800 450136 281852
rect 121552 281596 121604 281648
rect 148324 281596 148376 281648
rect 311716 281596 311768 281648
rect 313372 281596 313424 281648
rect 354588 281596 354640 281648
rect 121460 281528 121512 281580
rect 158076 281528 158128 281580
rect 295340 281528 295392 281580
rect 298284 281528 298336 281580
rect 349896 281528 349948 281580
rect 376944 281528 376996 281580
rect 360016 280848 360068 280900
rect 371240 280848 371292 280900
rect 56324 280780 56376 280832
rect 67640 280780 67692 280832
rect 125140 280780 125192 280832
rect 163688 280780 163740 280832
rect 300308 280780 300360 280832
rect 376208 280780 376260 280832
rect 476120 280780 476172 280832
rect 496084 280780 496136 280832
rect 52184 280168 52236 280220
rect 67640 280168 67692 280220
rect 121460 280168 121512 280220
rect 134800 280168 134852 280220
rect 371240 280168 371292 280220
rect 372528 280168 372580 280220
rect 376944 280168 376996 280220
rect 442816 280168 442868 280220
rect 476120 280168 476172 280220
rect 174636 280100 174688 280152
rect 176660 280100 176712 280152
rect 31024 279420 31076 279472
rect 67456 279420 67508 279472
rect 67640 279420 67692 279472
rect 122656 279420 122708 279472
rect 160836 279420 160888 279472
rect 296536 279420 296588 279472
rect 351276 279420 351328 279472
rect 39948 278740 40000 278792
rect 58624 278740 58676 278792
rect 121460 278740 121512 278792
rect 145564 278740 145616 278792
rect 67640 278672 67692 278724
rect 121552 278672 121604 278724
rect 132408 278672 132460 278724
rect 152648 278128 152700 278180
rect 166724 278128 166776 278180
rect 132408 278060 132460 278112
rect 164884 278060 164936 278112
rect 122748 277992 122800 278044
rect 169208 277992 169260 278044
rect 305736 277992 305788 278044
rect 371976 277992 372028 278044
rect 375196 277584 375248 277636
rect 376760 277584 376812 277636
rect 53656 277380 53708 277432
rect 67640 277380 67692 277432
rect 121460 277312 121512 277364
rect 126428 277380 126480 277432
rect 142896 277380 142948 277432
rect 166724 277380 166776 277432
rect 176660 277380 176712 277432
rect 373908 277380 373960 277432
rect 375196 277380 375248 277432
rect 442632 277380 442684 277432
rect 467932 277380 467984 277432
rect 56416 276632 56468 276684
rect 67640 276632 67692 276684
rect 293040 276632 293092 276684
rect 299572 276700 299624 276752
rect 300308 276700 300360 276752
rect 308496 276632 308548 276684
rect 355508 276632 355560 276684
rect 46848 276020 46900 276072
rect 67732 276020 67784 276072
rect 121460 276020 121512 276072
rect 166264 276020 166316 276072
rect 371976 276020 372028 276072
rect 377772 276020 377824 276072
rect 54852 275952 54904 276004
rect 55128 275952 55180 276004
rect 67640 275952 67692 276004
rect 123668 275272 123720 275324
rect 160100 275272 160152 275324
rect 301320 275272 301372 275324
rect 376116 275272 376168 275324
rect 121460 274728 121512 274780
rect 144460 274728 144512 274780
rect 160100 274728 160152 274780
rect 161296 274728 161348 274780
rect 176660 274728 176712 274780
rect 121552 274660 121604 274712
rect 170588 274660 170640 274712
rect 295340 274660 295392 274712
rect 300860 274660 300912 274712
rect 301320 274660 301372 274712
rect 121460 274592 121512 274644
rect 170496 274592 170548 274644
rect 41328 273912 41380 273964
rect 56508 273912 56560 273964
rect 306288 273912 306340 273964
rect 359648 273912 359700 273964
rect 463608 273912 463660 273964
rect 531964 273912 532016 273964
rect 121460 273368 121512 273420
rect 123484 273368 123536 273420
rect 66168 273300 66220 273352
rect 67824 273300 67876 273352
rect 56232 273232 56284 273284
rect 56508 273232 56560 273284
rect 67640 273232 67692 273284
rect 359648 273232 359700 273284
rect 360016 273232 360068 273284
rect 377772 273232 377824 273284
rect 442724 273232 442776 273284
rect 462320 273232 462372 273284
rect 463608 273232 463660 273284
rect 121460 272552 121512 272604
rect 121644 272552 121696 272604
rect 143080 272552 143132 272604
rect 120816 272484 120868 272536
rect 130568 272484 130620 272536
rect 158720 272484 158772 272536
rect 442816 272076 442868 272128
rect 448612 272076 448664 272128
rect 66076 271872 66128 271924
rect 67640 271872 67692 271924
rect 158720 271872 158772 271924
rect 160008 271872 160060 271924
rect 176660 271872 176712 271924
rect 295340 271872 295392 271924
rect 301688 271872 301740 271924
rect 176292 271804 176344 271856
rect 179696 271804 179748 271856
rect 296536 271804 296588 271856
rect 298100 271804 298152 271856
rect 64788 270580 64840 270632
rect 67732 270580 67784 270632
rect 41328 270512 41380 270564
rect 54484 270512 54536 270564
rect 59176 270512 59228 270564
rect 67640 270512 67692 270564
rect 121460 270512 121512 270564
rect 152740 270512 152792 270564
rect 67732 270444 67784 270496
rect 165528 269764 165580 269816
rect 177304 269764 177356 269816
rect 121460 269152 121512 269204
rect 130568 269152 130620 269204
rect 61844 269084 61896 269136
rect 67640 269084 67692 269136
rect 121552 269084 121604 269136
rect 151268 269084 151320 269136
rect 442264 269084 442316 269136
rect 448796 269084 448848 269136
rect 121460 269016 121512 269068
rect 160744 269016 160796 269068
rect 126888 268948 126940 269000
rect 130384 268948 130436 269000
rect 121368 268336 121420 268388
rect 163688 268336 163740 268388
rect 294236 268336 294288 268388
rect 299388 268336 299440 268388
rect 356704 268336 356756 268388
rect 35716 267792 35768 267844
rect 67640 267792 67692 267844
rect 3516 267656 3568 267708
rect 8208 267724 8260 267776
rect 48964 267724 49016 267776
rect 53472 267724 53524 267776
rect 67732 267724 67784 267776
rect 121460 267724 121512 267776
rect 126888 267724 126940 267776
rect 161388 267724 161440 267776
rect 176660 267724 176712 267776
rect 45284 267656 45336 267708
rect 67640 267656 67692 267708
rect 301504 267656 301556 267708
rect 379244 267656 379296 267708
rect 59084 267588 59136 267640
rect 67732 267588 67784 267640
rect 125048 267044 125100 267096
rect 169024 267044 169076 267096
rect 122472 266976 122524 267028
rect 169300 266976 169352 267028
rect 442816 266364 442868 266416
rect 460204 266364 460256 266416
rect 49424 266296 49476 266348
rect 67640 266296 67692 266348
rect 152556 266296 152608 266348
rect 176660 266296 176712 266348
rect 542360 266296 542412 266348
rect 133328 265684 133380 265736
rect 163504 265684 163556 265736
rect 121460 265616 121512 265668
rect 125508 265616 125560 265668
rect 174544 265616 174596 265668
rect 442356 265072 442408 265124
rect 444656 265072 444708 265124
rect 364156 264936 364208 264988
rect 376944 264936 376996 264988
rect 49516 263644 49568 263696
rect 67640 263644 67692 263696
rect 8944 263576 8996 263628
rect 54852 263576 54904 263628
rect 67732 263576 67784 263628
rect 121460 263576 121512 263628
rect 171876 263576 171928 263628
rect 376576 263576 376628 263628
rect 377496 263576 377548 263628
rect 121552 263508 121604 263560
rect 132500 263508 132552 263560
rect 133788 263508 133840 263560
rect 296352 263508 296404 263560
rect 345756 263508 345808 263560
rect 353944 263508 353996 263560
rect 377312 263508 377364 263560
rect 121460 262828 121512 262880
rect 153200 262828 153252 262880
rect 153936 262828 153988 262880
rect 60372 262284 60424 262336
rect 67732 262284 67784 262336
rect 55128 262216 55180 262268
rect 67640 262216 67692 262268
rect 442724 262216 442776 262268
rect 467104 262216 467156 262268
rect 60556 262148 60608 262200
rect 67732 262148 67784 262200
rect 121460 262148 121512 262200
rect 171140 262148 171192 262200
rect 302884 262148 302936 262200
rect 303712 262148 303764 262200
rect 61936 262080 61988 262132
rect 67640 262080 67692 262132
rect 158168 261468 158220 261520
rect 158628 261468 158680 261520
rect 176660 261468 176712 261520
rect 442816 261468 442868 261520
rect 570604 261468 570656 261520
rect 295340 261128 295392 261180
rect 299388 261128 299440 261180
rect 304448 261128 304500 261180
rect 303712 260856 303764 260908
rect 379336 260856 379388 260908
rect 21364 260788 21416 260840
rect 67640 260788 67692 260840
rect 121460 260788 121512 260840
rect 127164 260788 127216 260840
rect 127440 260788 127492 260840
rect 63316 260720 63368 260772
rect 67732 260720 67784 260772
rect 127440 260176 127492 260228
rect 149980 260176 150032 260228
rect 121644 260108 121696 260160
rect 167828 260108 167880 260160
rect 121460 259428 121512 259480
rect 131948 259428 132000 259480
rect 293868 259360 293920 259412
rect 308404 259360 308456 259412
rect 365260 259360 365312 259412
rect 371056 259360 371108 259412
rect 440240 259360 440292 259412
rect 454040 259360 454092 259412
rect 446496 259292 446548 259344
rect 448612 259292 448664 259344
rect 3976 258680 4028 258732
rect 62856 258680 62908 258732
rect 57796 258068 57848 258120
rect 67732 258068 67784 258120
rect 121460 258068 121512 258120
rect 156696 258068 156748 258120
rect 371056 258068 371108 258120
rect 376944 258068 376996 258120
rect 448612 258068 448664 258120
rect 580172 258068 580224 258120
rect 53748 258000 53800 258052
rect 67640 258000 67692 258052
rect 18604 257320 18656 257372
rect 53748 257320 53800 257372
rect 121460 256776 121512 256828
rect 150072 256776 150124 256828
rect 121552 256708 121604 256760
rect 162308 256708 162360 256760
rect 140596 256640 140648 256692
rect 176660 256708 176712 256760
rect 295340 256708 295392 256760
rect 302332 256708 302384 256760
rect 379888 256708 379940 256760
rect 440516 256708 440568 256760
rect 446496 256708 446548 256760
rect 121460 256096 121512 256148
rect 127072 256096 127124 256148
rect 122196 256028 122248 256080
rect 130384 256028 130436 256080
rect 63408 255960 63460 256012
rect 67640 255960 67692 256012
rect 122472 255960 122524 256012
rect 155316 255960 155368 256012
rect 318616 255960 318668 256012
rect 377312 255960 377364 256012
rect 127072 255348 127124 255400
rect 127624 255348 127676 255400
rect 60556 255280 60608 255332
rect 67732 255280 67784 255332
rect 121460 255280 121512 255332
rect 152648 255280 152700 255332
rect 166632 255212 166684 255264
rect 176660 255212 176712 255264
rect 295340 254532 295392 254584
rect 300124 254532 300176 254584
rect 300768 254532 300820 254584
rect 61660 253988 61712 254040
rect 67640 253988 67692 254040
rect 123668 253988 123720 254040
rect 164148 253988 164200 254040
rect 166632 253988 166684 254040
rect 61936 253920 61988 253972
rect 67732 253920 67784 253972
rect 121460 253920 121512 253972
rect 173164 253920 173216 253972
rect 36820 253852 36872 253904
rect 37004 253852 37056 253904
rect 67640 253852 67692 253904
rect 121552 253852 121604 253904
rect 140044 253852 140096 253904
rect 4804 253172 4856 253224
rect 36820 253172 36872 253224
rect 300768 253172 300820 253224
rect 373264 253172 373316 253224
rect 64512 252560 64564 252612
rect 66904 252560 66956 252612
rect 67548 252560 67600 252612
rect 121460 252560 121512 252612
rect 158168 252560 158220 252612
rect 62028 252492 62080 252544
rect 67640 252492 67692 252544
rect 296628 251880 296680 251932
rect 311164 251880 311216 251932
rect 56416 251812 56468 251864
rect 68284 251812 68336 251864
rect 297456 251812 297508 251864
rect 368296 251812 368348 251864
rect 442908 251812 442960 251864
rect 448520 251812 448572 251864
rect 462412 251812 462464 251864
rect 295340 251744 295392 251796
rect 297364 251744 297416 251796
rect 121552 251268 121604 251320
rect 159548 251268 159600 251320
rect 121460 251200 121512 251252
rect 170680 251200 170732 251252
rect 368296 251200 368348 251252
rect 376944 251200 376996 251252
rect 442724 251200 442776 251252
rect 460940 251200 460992 251252
rect 120632 251132 120684 251184
rect 132592 251132 132644 251184
rect 295340 250452 295392 250504
rect 296628 250452 296680 250504
rect 300124 250452 300176 250504
rect 57704 249840 57756 249892
rect 67640 249840 67692 249892
rect 121460 249772 121512 249824
rect 133236 249772 133288 249824
rect 52276 249704 52328 249756
rect 67640 249704 67692 249756
rect 121552 249704 121604 249756
rect 129740 249704 129792 249756
rect 121460 249636 121512 249688
rect 129188 249636 129240 249688
rect 119804 249092 119856 249144
rect 130660 249092 130712 249144
rect 129740 249024 129792 249076
rect 175924 249024 175976 249076
rect 65800 248616 65852 248668
rect 68008 248616 68060 248668
rect 121460 248344 121512 248396
rect 162124 248344 162176 248396
rect 295340 248344 295392 248396
rect 316132 248344 316184 248396
rect 317236 248344 317288 248396
rect 317236 247664 317288 247716
rect 373356 247664 373408 247716
rect 63224 247120 63276 247172
rect 67640 247120 67692 247172
rect 59084 247052 59136 247104
rect 67732 247052 67784 247104
rect 121552 247052 121604 247104
rect 129188 247052 129240 247104
rect 362960 247052 363012 247104
rect 376944 247052 376996 247104
rect 50804 246984 50856 247036
rect 67640 246984 67692 247036
rect 65984 246916 66036 246968
rect 68100 246916 68152 246968
rect 301044 246508 301096 246560
rect 301596 246508 301648 246560
rect 294328 246304 294380 246356
rect 301044 246304 301096 246356
rect 318708 246304 318760 246356
rect 362960 246304 363012 246356
rect 363696 246304 363748 246356
rect 442908 246304 442960 246356
rect 534080 246304 534132 246356
rect 121552 245760 121604 245812
rect 124956 245760 125008 245812
rect 121460 245692 121512 245744
rect 148416 245692 148468 245744
rect 131856 245624 131908 245676
rect 164056 245624 164108 245676
rect 176660 245624 176712 245676
rect 318064 245624 318116 245676
rect 318708 245624 318760 245676
rect 364708 245624 364760 245676
rect 365628 245624 365680 245676
rect 376944 245624 376996 245676
rect 26148 245556 26200 245608
rect 67640 245556 67692 245608
rect 121460 245556 121512 245608
rect 167000 245556 167052 245608
rect 467104 245556 467156 245608
rect 533988 245556 534040 245608
rect 580172 245556 580224 245608
rect 121552 244264 121604 244316
rect 147496 244264 147548 244316
rect 35808 244196 35860 244248
rect 67640 244196 67692 244248
rect 121644 244196 121696 244248
rect 135996 244196 136048 244248
rect 17224 244128 17276 244180
rect 43996 244128 44048 244180
rect 67732 244128 67784 244180
rect 121460 244128 121512 244180
rect 126244 244128 126296 244180
rect 159456 243516 159508 243568
rect 171784 243516 171836 243568
rect 128360 242904 128412 242956
rect 129648 242904 129700 242956
rect 162124 242904 162176 242956
rect 296260 242904 296312 242956
rect 300952 242904 301004 242956
rect 318156 242904 318208 242956
rect 357532 242904 357584 242956
rect 358820 242904 358872 242956
rect 442172 242904 442224 242956
rect 443276 242904 443328 242956
rect 121460 242836 121512 242888
rect 138848 242836 138900 242888
rect 121552 242768 121604 242820
rect 128360 242768 128412 242820
rect 142988 242292 143040 242344
rect 175004 242292 175056 242344
rect 145656 242224 145708 242276
rect 179880 242224 179932 242276
rect 63408 242156 63460 242208
rect 69664 242156 69716 242208
rect 119988 242156 120040 242208
rect 170496 242156 170548 242208
rect 442908 242156 442960 242208
rect 444472 242156 444524 242208
rect 63316 241544 63368 241596
rect 67640 241544 67692 241596
rect 61752 241476 61804 241528
rect 67732 241476 67784 241528
rect 175004 241476 175056 241528
rect 176660 241476 176712 241528
rect 53564 241408 53616 241460
rect 67640 241408 67692 241460
rect 296444 241408 296496 241460
rect 296628 241408 296680 241460
rect 300216 241408 300268 241460
rect 150072 240864 150124 240916
rect 155776 240796 155828 240848
rect 42708 240728 42760 240780
rect 67640 240728 67692 240780
rect 127624 240728 127676 240780
rect 179512 240728 179564 240780
rect 184204 240592 184256 240644
rect 284208 240592 284260 240644
rect 306380 240796 306432 240848
rect 372528 240796 372580 240848
rect 301136 240728 301188 240780
rect 301688 240728 301740 240780
rect 381544 240660 381596 240712
rect 476120 240728 476172 240780
rect 191932 240456 191984 240508
rect 121460 240116 121512 240168
rect 149888 240116 149940 240168
rect 3424 240048 3476 240100
rect 48228 240048 48280 240100
rect 148508 240048 148560 240100
rect 301136 240048 301188 240100
rect 310428 240048 310480 240100
rect 310612 240048 310664 240100
rect 439504 239640 439556 239692
rect 444564 239640 444616 239692
rect 395988 239504 396040 239556
rect 440424 239504 440476 239556
rect 117136 239436 117188 239488
rect 134616 239436 134668 239488
rect 158628 239436 158680 239488
rect 220176 239436 220228 239488
rect 382188 239436 382240 239488
rect 441712 239436 441764 239488
rect 48228 239368 48280 239420
rect 71688 239368 71740 239420
rect 116768 239368 116820 239420
rect 136732 239368 136784 239420
rect 161296 239368 161348 239420
rect 323400 239368 323452 239420
rect 382096 239368 382148 239420
rect 441620 239368 441672 239420
rect 443736 239368 443788 239420
rect 580264 239368 580316 239420
rect 189080 239096 189132 239148
rect 190184 239096 190236 239148
rect 382188 239096 382240 239148
rect 64696 239028 64748 239080
rect 70032 239028 70084 239080
rect 316132 239028 316184 239080
rect 317328 239028 317380 239080
rect 390468 239028 390520 239080
rect 60464 238960 60516 239012
rect 80336 238960 80388 239012
rect 119988 238960 120040 239012
rect 125048 238960 125100 239012
rect 263048 238960 263100 239012
rect 297548 238960 297600 239012
rect 376024 238960 376076 239012
rect 435364 238960 435416 239012
rect 438584 238960 438636 239012
rect 59268 238892 59320 238944
rect 91284 238892 91336 238944
rect 117228 238892 117280 238944
rect 210516 238892 210568 238944
rect 219440 238892 219492 238944
rect 382096 238892 382148 238944
rect 390468 238892 390520 238944
rect 438860 238892 438912 238944
rect 48964 238824 49016 238876
rect 85580 238824 85632 238876
rect 99012 238824 99064 238876
rect 120816 238824 120868 238876
rect 173348 238824 173400 238876
rect 215300 238824 215352 238876
rect 269212 238824 269264 238876
rect 395988 238824 396040 238876
rect 37096 238756 37148 238808
rect 81624 238756 81676 238808
rect 91928 238756 91980 238808
rect 144184 238756 144236 238808
rect 179512 238756 179564 238808
rect 189080 238756 189132 238808
rect 223764 238756 223816 238808
rect 269120 238756 269172 238808
rect 379612 238756 379664 238808
rect 398932 238756 398984 238808
rect 399944 238756 399996 238808
rect 436744 238756 436796 238808
rect 443092 238756 443144 238808
rect 3332 238688 3384 238740
rect 55036 238688 55088 238740
rect 103520 238688 103572 238740
rect 114468 238688 114520 238740
rect 117136 238688 117188 238740
rect 118976 238688 119028 238740
rect 131856 238688 131908 238740
rect 178684 238688 178736 238740
rect 196440 238688 196492 238740
rect 204812 238688 204864 238740
rect 376576 238688 376628 238740
rect 424324 238688 424376 238740
rect 438584 238688 438636 238740
rect 443736 238688 443788 238740
rect 71688 238620 71740 238672
rect 112536 238620 112588 238672
rect 117228 238620 117280 238672
rect 117688 238620 117740 238672
rect 250536 238620 250588 238672
rect 264980 238620 265032 238672
rect 279424 238620 279476 238672
rect 296536 238620 296588 238672
rect 387248 238620 387300 238672
rect 420184 238620 420236 238672
rect 458272 238620 458324 238672
rect 57888 238552 57940 238604
rect 74540 238552 74592 238604
rect 85580 238552 85632 238604
rect 86776 238552 86828 238604
rect 117044 238552 117096 238604
rect 123668 238552 123720 238604
rect 219348 238552 219400 238604
rect 341524 238552 341576 238604
rect 407764 238552 407816 238604
rect 50896 238484 50948 238536
rect 73252 238484 73304 238536
rect 118332 238484 118384 238536
rect 240140 238484 240192 238536
rect 75828 238416 75880 238468
rect 80888 238416 80940 238468
rect 115112 238416 115164 238468
rect 236368 238416 236420 238468
rect 296536 238416 296588 238468
rect 108028 238348 108080 238400
rect 119988 238348 120040 238400
rect 196440 238348 196492 238400
rect 219440 238348 219492 238400
rect 253204 238348 253256 238400
rect 307208 238484 307260 238536
rect 393596 238484 393648 238536
rect 312636 238416 312688 238468
rect 384304 238416 384356 238468
rect 240140 238280 240192 238332
rect 315304 238280 315356 238332
rect 46664 238008 46716 238060
rect 77208 238008 77260 238060
rect 86776 238008 86828 238060
rect 208492 238008 208544 238060
rect 257620 238008 257672 238060
rect 262128 238008 262180 238060
rect 291200 238008 291252 238060
rect 312636 238008 312688 238060
rect 315304 238008 315356 238060
rect 405648 238008 405700 238060
rect 432236 238008 432288 238060
rect 454040 238008 454092 238060
rect 456892 238008 456944 238060
rect 77208 237804 77260 237856
rect 77760 237804 77812 237856
rect 422300 237668 422352 237720
rect 426348 237668 426400 237720
rect 74540 237396 74592 237448
rect 75184 237396 75236 237448
rect 79048 237396 79100 237448
rect 80796 237396 80848 237448
rect 82084 237396 82136 237448
rect 82912 237396 82964 237448
rect 208492 237396 208544 237448
rect 209688 237396 209740 237448
rect 210608 237396 210660 237448
rect 432696 237396 432748 237448
rect 434076 237396 434128 237448
rect 46756 237328 46808 237380
rect 107384 237328 107436 237380
rect 116768 237328 116820 237380
rect 172336 237328 172388 237380
rect 458364 237328 458416 237380
rect 54760 237260 54812 237312
rect 325700 237260 325752 237312
rect 326344 237260 326396 237312
rect 357348 237260 357400 237312
rect 411904 237260 411956 237312
rect 54944 237192 54996 237244
rect 89352 237192 89404 237244
rect 106740 237192 106792 237244
rect 140596 237192 140648 237244
rect 156696 237192 156748 237244
rect 276020 237192 276072 237244
rect 288256 237192 288308 237244
rect 313372 237192 313424 237244
rect 325148 237192 325200 237244
rect 422300 237192 422352 237244
rect 45468 237124 45520 237176
rect 77116 237124 77168 237176
rect 88708 237124 88760 237176
rect 120724 237124 120776 237176
rect 179880 237124 179932 237176
rect 204812 237124 204864 237176
rect 284668 237124 284720 237176
rect 285588 237124 285640 237176
rect 308496 237124 308548 237176
rect 375104 237124 375156 237176
rect 402980 237124 403032 237176
rect 403808 237124 403860 237176
rect 115848 237056 115900 237108
rect 133328 237056 133380 237108
rect 86132 236988 86184 237040
rect 130476 236988 130528 237040
rect 429108 236920 429160 236972
rect 440240 236920 440292 236972
rect 443184 236920 443236 236972
rect 459744 236920 459796 236972
rect 426440 236852 426492 236904
rect 451280 236852 451332 236904
rect 414020 236784 414072 236836
rect 449992 236784 450044 236836
rect 163688 236716 163740 236768
rect 193956 236716 194008 236768
rect 261484 236716 261536 236768
rect 291844 236716 291896 236768
rect 394608 236716 394660 236768
rect 452844 236716 452896 236768
rect 140596 236648 140648 236700
rect 288532 236648 288584 236700
rect 378048 236648 378100 236700
rect 392584 236648 392636 236700
rect 432604 236648 432656 236700
rect 561680 236648 561732 236700
rect 76564 235968 76616 236020
rect 77116 235968 77168 236020
rect 393596 235968 393648 236020
rect 395344 235968 395396 236020
rect 250536 235900 250588 235952
rect 316132 235900 316184 235952
rect 373356 235900 373408 235952
rect 467932 235900 467984 235952
rect 37188 235832 37240 235884
rect 94412 235832 94464 235884
rect 95148 235832 95200 235884
rect 113824 235832 113876 235884
rect 138020 235832 138072 235884
rect 166724 235832 166776 235884
rect 358084 235832 358136 235884
rect 368388 235832 368440 235884
rect 398104 235832 398156 235884
rect 48136 235764 48188 235816
rect 79324 235764 79376 235816
rect 109684 235764 109736 235816
rect 125140 235764 125192 235816
rect 155316 235764 155368 235816
rect 269212 235764 269264 235816
rect 269304 235764 269356 235816
rect 317420 235764 317472 235816
rect 377404 235764 377456 235816
rect 159548 235696 159600 235748
rect 273996 235696 274048 235748
rect 286600 235696 286652 235748
rect 286876 235696 286928 235748
rect 307116 235696 307168 235748
rect 347044 235696 347096 235748
rect 402244 235696 402296 235748
rect 234068 235628 234120 235680
rect 318064 235628 318116 235680
rect 352564 235628 352616 235680
rect 391296 235628 391348 235680
rect 61936 235560 61988 235612
rect 263048 235560 263100 235612
rect 67640 235220 67692 235272
rect 242164 235220 242216 235272
rect 323400 235220 323452 235272
rect 397368 235220 397420 235272
rect 448796 235220 448848 235272
rect 289820 234608 289872 234660
rect 294144 234608 294196 234660
rect 349896 234608 349948 234660
rect 353392 234608 353444 234660
rect 35164 234540 35216 234592
rect 35716 234540 35768 234592
rect 303620 234540 303672 234592
rect 321376 234540 321428 234592
rect 326528 234540 326580 234592
rect 331312 234540 331364 234592
rect 332508 234540 332560 234592
rect 376116 234540 376168 234592
rect 95792 234472 95844 234524
rect 146944 234472 146996 234524
rect 277952 234472 278004 234524
rect 449900 234472 449952 234524
rect 162124 234404 162176 234456
rect 331312 234404 331364 234456
rect 276020 234336 276072 234388
rect 311900 234336 311952 234388
rect 100300 233996 100352 234048
rect 117964 233996 118016 234048
rect 151360 233996 151412 234048
rect 215944 233996 215996 234048
rect 84200 233928 84252 233980
rect 84844 233928 84896 233980
rect 95240 233928 95292 233980
rect 96436 233928 96488 233980
rect 104808 233928 104860 233980
rect 210424 233928 210476 233980
rect 221556 233928 221608 233980
rect 271236 233928 271288 233980
rect 311900 233928 311952 233980
rect 312728 233928 312780 233980
rect 353944 233928 353996 233980
rect 377404 233928 377456 233980
rect 387064 233928 387116 233980
rect 27528 233860 27580 233912
rect 113088 233860 113140 233912
rect 169300 233860 169352 233912
rect 321376 233860 321428 233912
rect 349804 233860 349856 233912
rect 408500 233860 408552 233912
rect 444656 233860 444708 233912
rect 485780 233860 485832 233912
rect 582380 233860 582432 233912
rect 385868 233248 385920 233300
rect 39764 233112 39816 233164
rect 71964 233180 72016 233232
rect 72424 233180 72476 233232
rect 102232 233180 102284 233232
rect 103428 233180 103480 233232
rect 151084 233180 151136 233232
rect 158260 233180 158312 233232
rect 321560 233180 321612 233232
rect 579988 233180 580040 233232
rect 76472 233112 76524 233164
rect 135904 233112 135956 233164
rect 152648 233112 152700 233164
rect 299572 233112 299624 233164
rect 337384 233112 337436 233164
rect 431960 233112 432012 233164
rect 432696 233112 432748 233164
rect 52368 233044 52420 233096
rect 80704 233044 80756 233096
rect 98368 233044 98420 233096
rect 234068 233044 234120 233096
rect 271236 233044 271288 233096
rect 304264 233044 304316 233096
rect 382280 233044 382332 233096
rect 450084 233044 450136 233096
rect 83556 232976 83608 233028
rect 126336 232976 126388 233028
rect 129096 232976 129148 233028
rect 223764 232976 223816 233028
rect 356796 232976 356848 233028
rect 410524 232976 410576 233028
rect 32956 232908 33008 232960
rect 104164 232908 104216 232960
rect 382004 232568 382056 232620
rect 388444 232568 388496 232620
rect 369676 232500 369728 232552
rect 387156 232500 387208 232552
rect 450084 232296 450136 232348
rect 450544 232296 450596 232348
rect 110420 232160 110472 232212
rect 111248 232160 111300 232212
rect 61752 231752 61804 231804
rect 264060 231752 264112 231804
rect 314476 231752 314528 231804
rect 314752 231752 314804 231804
rect 31668 231684 31720 231736
rect 106188 231684 106240 231736
rect 166908 231684 166960 231736
rect 198740 231684 198792 231736
rect 199384 231684 199436 231736
rect 214564 231684 214616 231736
rect 362960 231684 363012 231736
rect 93952 231548 94004 231600
rect 94504 231548 94556 231600
rect 278780 231344 278832 231396
rect 294236 231344 294288 231396
rect 167736 231276 167788 231328
rect 279424 231276 279476 231328
rect 106188 231208 106240 231260
rect 243544 231208 243596 231260
rect 248420 231208 248472 231260
rect 282184 231208 282236 231260
rect 296812 231208 296864 231260
rect 301044 231208 301096 231260
rect 391204 231208 391256 231260
rect 141608 231140 141660 231192
rect 314476 231140 314528 231192
rect 78404 231072 78456 231124
rect 126244 231072 126296 231124
rect 158168 231072 158220 231124
rect 220084 231072 220136 231124
rect 220176 231072 220228 231124
rect 426624 231072 426676 231124
rect 451372 231072 451424 231124
rect 289084 231004 289136 231056
rect 295616 231004 295668 231056
rect 59176 230392 59228 230444
rect 288256 230392 288308 230444
rect 297364 230392 297416 230444
rect 365076 230392 365128 230444
rect 396080 230392 396132 230444
rect 143080 230324 143132 230376
rect 300860 230324 300912 230376
rect 184204 230256 184256 230308
rect 310520 230256 310572 230308
rect 396080 229984 396132 230036
rect 396724 229984 396776 230036
rect 171876 229848 171928 229900
rect 189724 229848 189776 229900
rect 371148 229848 371200 229900
rect 458272 229848 458324 229900
rect 64512 229780 64564 229832
rect 98644 229780 98696 229832
rect 131948 229780 132000 229832
rect 203524 229780 203576 229832
rect 244280 229780 244332 229832
rect 266268 229780 266320 229832
rect 305736 229780 305788 229832
rect 3424 229712 3476 229764
rect 120172 229712 120224 229764
rect 165068 229712 165120 229764
rect 261484 229712 261536 229764
rect 281540 229712 281592 229764
rect 386328 229780 386380 229832
rect 489184 229780 489236 229832
rect 418804 229712 418856 229764
rect 533344 229712 533396 229764
rect 61660 229032 61712 229084
rect 297364 229032 297416 229084
rect 56324 228488 56376 228540
rect 158168 228488 158220 228540
rect 314568 228488 314620 228540
rect 351184 228488 351236 228540
rect 122288 228420 122340 228472
rect 320088 228420 320140 228472
rect 379244 228420 379296 228472
rect 409880 228420 409932 228472
rect 157156 228352 157208 228404
rect 377956 228352 378008 228404
rect 467104 228352 467156 228404
rect 231860 227740 231912 227792
rect 233148 227740 233200 227792
rect 149980 227672 150032 227724
rect 448704 227672 448756 227724
rect 56232 227604 56284 227656
rect 242256 227604 242308 227656
rect 105452 227536 105504 227588
rect 172428 227536 172480 227588
rect 185584 227536 185636 227588
rect 323584 227536 323636 227588
rect 284116 227060 284168 227112
rect 347780 227060 347832 227112
rect 172428 226992 172480 227044
rect 345572 226992 345624 227044
rect 399116 226992 399168 227044
rect 441620 226992 441672 227044
rect 448704 226380 448756 226432
rect 449164 226380 449216 226432
rect 245660 226312 245712 226364
rect 246948 226312 247000 226364
rect 323032 226312 323084 226364
rect 323584 226312 323636 226364
rect 160008 226244 160060 226296
rect 415400 226244 415452 226296
rect 455512 226312 455564 226364
rect 167828 226176 167880 226228
rect 327264 226176 327316 226228
rect 327724 226176 327776 226228
rect 345572 226176 345624 226228
rect 345756 226176 345808 226228
rect 474740 226176 474792 226228
rect 210516 226108 210568 226160
rect 303712 226108 303764 226160
rect 123576 225632 123628 225684
rect 270316 225632 270368 225684
rect 59084 225564 59136 225616
rect 214564 225564 214616 225616
rect 319628 225564 319680 225616
rect 341524 225564 341576 225616
rect 49608 224884 49660 224936
rect 302332 224884 302384 224936
rect 54852 224816 54904 224868
rect 253204 224816 253256 224868
rect 169208 224748 169260 224800
rect 342996 224748 343048 224800
rect 88064 224272 88116 224324
rect 249800 224272 249852 224324
rect 281448 224272 281500 224324
rect 299480 224272 299532 224324
rect 175096 224204 175148 224256
rect 579620 224204 579672 224256
rect 80888 223524 80940 223576
rect 305000 223524 305052 223576
rect 93952 223456 94004 223508
rect 136640 223456 136692 223508
rect 137100 223456 137152 223508
rect 193220 223456 193272 223508
rect 194508 223456 194560 223508
rect 209688 223456 209740 223508
rect 371976 223456 372028 223508
rect 144460 223388 144512 223440
rect 296812 223388 296864 223440
rect 194508 223320 194560 223372
rect 345848 223320 345900 223372
rect 170588 222980 170640 223032
rect 196624 222980 196676 223032
rect 137100 222912 137152 222964
rect 170680 222912 170732 222964
rect 300124 222912 300176 222964
rect 334716 222912 334768 222964
rect 104164 222844 104216 222896
rect 264244 222844 264296 222896
rect 270316 222844 270368 222896
rect 315948 222844 316000 222896
rect 318800 222844 318852 222896
rect 153936 222096 153988 222148
rect 434720 222096 434772 222148
rect 436008 222096 436060 222148
rect 57704 222028 57756 222080
rect 328552 222028 328604 222080
rect 329196 222028 329248 222080
rect 82084 221960 82136 222012
rect 298284 221960 298336 222012
rect 101588 221484 101640 221536
rect 253940 221484 253992 221536
rect 63316 221416 63368 221468
rect 240784 221416 240836 221468
rect 436008 221416 436060 221468
rect 461032 221416 461084 221468
rect 99656 220736 99708 220788
rect 168932 220736 168984 220788
rect 173256 220260 173308 220312
rect 236644 220260 236696 220312
rect 67364 220192 67416 220244
rect 156696 220192 156748 220244
rect 168932 220192 168984 220244
rect 169576 220192 169628 220244
rect 318064 220192 318116 220244
rect 64604 220124 64656 220176
rect 251180 220124 251232 220176
rect 154396 220056 154448 220108
rect 393228 220056 393280 220108
rect 414204 220056 414256 220108
rect 69664 219376 69716 219428
rect 331864 219376 331916 219428
rect 162768 219308 162820 219360
rect 420920 219308 420972 219360
rect 148324 218832 148376 218884
rect 210516 218832 210568 218884
rect 130568 218764 130620 218816
rect 221464 218764 221516 218816
rect 229100 218764 229152 218816
rect 275928 218764 275980 218816
rect 324964 218764 325016 218816
rect 331312 218764 331364 218816
rect 331864 218764 331916 218816
rect 361488 218764 361540 218816
rect 388628 218764 388680 218816
rect 153844 218696 153896 218748
rect 300124 218696 300176 218748
rect 364248 218696 364300 218748
rect 380164 218696 380216 218748
rect 380808 218696 380860 218748
rect 433984 218696 434036 218748
rect 420920 218084 420972 218136
rect 421656 218084 421708 218136
rect 388628 218016 388680 218068
rect 389088 218016 389140 218068
rect 580172 218016 580224 218068
rect 142896 217948 142948 218000
rect 300952 217948 301004 218000
rect 385684 217948 385736 218000
rect 111892 217268 111944 217320
rect 270500 217268 270552 217320
rect 419448 217268 419500 217320
rect 526444 217268 526496 217320
rect 164056 216588 164108 216640
rect 378968 216588 379020 216640
rect 160928 216520 160980 216572
rect 334808 216520 334860 216572
rect 3516 216112 3568 216164
rect 8944 216112 8996 216164
rect 151176 215976 151228 216028
rect 276020 215976 276072 216028
rect 337384 215976 337436 216028
rect 439504 215976 439556 216028
rect 74724 215908 74776 215960
rect 252560 215908 252612 215960
rect 423588 215908 423640 215960
rect 530584 215908 530636 215960
rect 333980 215500 334032 215552
rect 334808 215500 334860 215552
rect 42800 215228 42852 215280
rect 44088 215228 44140 215280
rect 120080 215228 120132 215280
rect 147680 215228 147732 215280
rect 358820 215228 358872 215280
rect 359464 215228 359516 215280
rect 60372 215160 60424 215212
rect 291200 215160 291252 215212
rect 96712 215092 96764 215144
rect 147680 215092 147732 215144
rect 1308 214548 1360 214600
rect 42800 214548 42852 214600
rect 86960 213868 87012 213920
rect 144920 213868 144972 213920
rect 146208 213868 146260 213920
rect 146208 213460 146260 213512
rect 202144 213460 202196 213512
rect 141516 213392 141568 213444
rect 229744 213392 229796 213444
rect 133236 213324 133288 213376
rect 247684 213324 247736 213376
rect 271880 213324 271932 213376
rect 293132 213324 293184 213376
rect 126888 213256 126940 213308
rect 273904 213256 273956 213308
rect 311256 213256 311308 213308
rect 404360 213256 404412 213308
rect 14464 213188 14516 213240
rect 83464 213188 83516 213240
rect 147588 213188 147640 213240
rect 391848 213188 391900 213240
rect 429200 213188 429252 213240
rect 77208 212440 77260 212492
rect 367100 212440 367152 212492
rect 164148 212372 164200 212424
rect 376668 212372 376720 212424
rect 382924 212372 382976 212424
rect 162216 211896 162268 211948
rect 274640 211896 274692 211948
rect 48044 211828 48096 211880
rect 211896 211828 211948 211880
rect 170680 211760 170732 211812
rect 346584 211760 346636 211812
rect 210424 211080 210476 211132
rect 335452 211080 335504 211132
rect 84384 210468 84436 210520
rect 264980 210468 265032 210520
rect 129004 210400 129056 210452
rect 345020 210400 345072 210452
rect 351920 210400 351972 210452
rect 377864 210400 377916 210452
rect 451648 210400 451700 210452
rect 41236 209720 41288 209772
rect 322848 209720 322900 209772
rect 95240 209652 95292 209704
rect 140688 209652 140740 209704
rect 147036 209244 147088 209296
rect 239496 209244 239548 209296
rect 171784 209176 171836 209228
rect 304264 209176 304316 209228
rect 140688 209108 140740 209160
rect 319444 209108 319496 209160
rect 398932 209108 398984 209160
rect 449992 209108 450044 209160
rect 43812 209040 43864 209092
rect 233884 209040 233936 209092
rect 371056 209040 371108 209092
rect 431224 209040 431276 209092
rect 311164 208360 311216 208412
rect 316040 208360 316092 208412
rect 49516 208292 49568 208344
rect 322940 208292 322992 208344
rect 124864 207816 124916 207868
rect 265072 207816 265124 207868
rect 131764 207748 131816 207800
rect 281540 207748 281592 207800
rect 102140 207680 102192 207732
rect 252744 207680 252796 207732
rect 61844 207612 61896 207664
rect 277492 207612 277544 207664
rect 110512 206932 110564 206984
rect 111064 206932 111116 206984
rect 153108 206932 153160 206984
rect 443092 206932 443144 206984
rect 476212 206932 476264 206984
rect 579988 206932 580040 206984
rect 107660 206864 107712 206916
rect 155868 206864 155920 206916
rect 227720 206864 227772 206916
rect 346492 206864 346544 206916
rect 347688 206864 347740 206916
rect 155868 206388 155920 206440
rect 257344 206388 257396 206440
rect 89812 206320 89864 206372
rect 252652 206320 252704 206372
rect 67548 206252 67600 206304
rect 280160 206252 280212 206304
rect 347688 206252 347740 206304
rect 452844 206252 452896 206304
rect 467104 206252 467156 206304
rect 476212 206252 476264 206304
rect 84292 205572 84344 205624
rect 125784 205572 125836 205624
rect 126888 205572 126940 205624
rect 158076 205164 158128 205216
rect 247776 205164 247828 205216
rect 151268 205096 151320 205148
rect 263600 205096 263652 205148
rect 126244 205028 126296 205080
rect 259552 205028 259604 205080
rect 66076 204960 66128 205012
rect 251272 204960 251324 205012
rect 373816 204960 373868 205012
rect 435456 204960 435508 205012
rect 179144 204892 179196 204944
rect 405740 204892 405792 204944
rect 421564 204892 421616 204944
rect 464344 204892 464396 204944
rect 126888 204280 126940 204332
rect 193864 204280 193916 204332
rect 84200 204212 84252 204264
rect 126980 204212 127032 204264
rect 127440 204212 127492 204264
rect 144368 203872 144420 203924
rect 242256 203872 242308 203924
rect 242164 203804 242216 203856
rect 351920 203804 351972 203856
rect 142804 203736 142856 203788
rect 277400 203736 277452 203788
rect 115940 203668 115992 203720
rect 254124 203668 254176 203720
rect 53656 203600 53708 203652
rect 267832 203600 267884 203652
rect 127440 203532 127492 203584
rect 352012 203532 352064 203584
rect 381544 203532 381596 203584
rect 458824 203532 458876 203584
rect 130660 202376 130712 202428
rect 246304 202376 246356 202428
rect 144276 202308 144328 202360
rect 192484 202308 192536 202360
rect 193956 202308 194008 202360
rect 335452 202308 335504 202360
rect 170404 202240 170456 202292
rect 316684 202240 316736 202292
rect 89720 202172 89772 202224
rect 252836 202172 252888 202224
rect 39948 202104 40000 202156
rect 287704 202104 287756 202156
rect 395896 202104 395948 202156
rect 444472 202104 444524 202156
rect 421656 201492 421708 201544
rect 422208 201492 422260 201544
rect 427084 201492 427136 201544
rect 246948 201424 247000 201476
rect 298008 201424 298060 201476
rect 196624 200948 196676 201000
rect 271972 200948 272024 201000
rect 110420 200880 110472 200932
rect 255596 200880 255648 200932
rect 57796 200812 57848 200864
rect 222844 200812 222896 200864
rect 79324 200744 79376 200796
rect 322940 200744 322992 200796
rect 298008 200132 298060 200184
rect 451372 200132 451424 200184
rect 233148 200064 233200 200116
rect 284116 200064 284168 200116
rect 117964 199452 118016 199504
rect 273260 199452 273312 199504
rect 94044 199384 94096 199436
rect 255412 199384 255464 199436
rect 282920 198704 282972 198756
rect 284116 198704 284168 198756
rect 451464 198704 451516 198756
rect 76564 198636 76616 198688
rect 330576 198636 330628 198688
rect 145564 198160 145616 198212
rect 232504 198160 232556 198212
rect 149704 198092 149756 198144
rect 269212 198092 269264 198144
rect 92480 198024 92532 198076
rect 261024 198024 261076 198076
rect 292672 198024 292724 198076
rect 441620 198024 441672 198076
rect 93768 197956 93820 198008
rect 356244 197956 356296 198008
rect 439504 197956 439556 198008
rect 538220 197956 538272 198008
rect 329840 197684 329892 197736
rect 330576 197684 330628 197736
rect 94504 197276 94556 197328
rect 354772 197276 354824 197328
rect 355324 197276 355376 197328
rect 335452 197208 335504 197260
rect 535460 197208 535512 197260
rect 141424 196732 141476 196784
rect 269120 196732 269172 196784
rect 133144 196664 133196 196716
rect 263692 196664 263744 196716
rect 70400 196596 70452 196648
rect 254032 196596 254084 196648
rect 98644 195916 98696 195968
rect 354864 195916 354916 195968
rect 355416 195916 355468 195968
rect 162308 195372 162360 195424
rect 267740 195372 267792 195424
rect 138664 195304 138716 195356
rect 281632 195304 281684 195356
rect 52184 195236 52236 195288
rect 236736 195236 236788 195288
rect 264244 195236 264296 195288
rect 356152 195236 356204 195288
rect 134708 194080 134760 194132
rect 262312 194080 262364 194132
rect 100760 194012 100812 194064
rect 278872 194012 278924 194064
rect 55128 193944 55180 193996
rect 239588 193944 239640 193996
rect 177672 193876 177724 193928
rect 376024 193876 376076 193928
rect 391296 193876 391348 193928
rect 454132 193876 454184 193928
rect 136088 193808 136140 193860
rect 338120 193808 338172 193860
rect 390376 193808 390428 193860
rect 520924 193808 520976 193860
rect 427084 193128 427136 193180
rect 580172 193128 580224 193180
rect 243544 192720 243596 192772
rect 327080 192720 327132 192772
rect 137284 192652 137336 192704
rect 247868 192652 247920 192704
rect 96620 192584 96672 192636
rect 258172 192584 258224 192636
rect 67456 192516 67508 192568
rect 251364 192516 251416 192568
rect 402244 192516 402296 192568
rect 435548 192516 435600 192568
rect 80796 192448 80848 192500
rect 270592 192448 270644 192500
rect 275836 192448 275888 192500
rect 293040 192448 293092 192500
rect 350632 192448 350684 192500
rect 416964 192448 417016 192500
rect 212540 191768 212592 191820
rect 368480 191768 368532 191820
rect 368940 191768 368992 191820
rect 398104 191768 398156 191820
rect 399484 191768 399536 191820
rect 161388 191224 161440 191276
rect 198004 191224 198056 191276
rect 149888 191156 149940 191208
rect 242164 191156 242216 191208
rect 63224 191088 63276 191140
rect 260840 191088 260892 191140
rect 368940 191088 368992 191140
rect 396080 191088 396132 191140
rect 407764 191088 407816 191140
rect 452936 191088 452988 191140
rect 148416 190000 148468 190052
rect 260932 190000 260984 190052
rect 46848 189932 46900 189984
rect 162124 189932 162176 189984
rect 203524 189932 203576 189984
rect 267924 189932 267976 189984
rect 129188 189864 129240 189916
rect 246396 189864 246448 189916
rect 134800 189796 134852 189848
rect 259460 189796 259512 189848
rect 261484 189796 261536 189848
rect 318156 189796 318208 189848
rect 420276 189796 420328 189848
rect 536932 189796 536984 189848
rect 136180 189728 136232 189780
rect 263784 189728 263836 189780
rect 307024 189728 307076 189780
rect 460204 189728 460256 189780
rect 107568 189048 107620 189100
rect 189908 189048 189960 189100
rect 307024 189048 307076 189100
rect 307668 189048 307720 189100
rect 459560 189048 459612 189100
rect 460204 189048 460256 189100
rect 3424 188980 3476 189032
rect 58716 188980 58768 189032
rect 214564 188640 214616 188692
rect 256976 188640 257028 188692
rect 239404 188572 239456 188624
rect 343824 188572 343876 188624
rect 123484 188504 123536 188556
rect 247960 188504 248012 188556
rect 124956 188436 125008 188488
rect 258080 188436 258132 188488
rect 160836 188368 160888 188420
rect 324596 188368 324648 188420
rect 72424 188300 72476 188352
rect 323124 188300 323176 188352
rect 363788 188300 363840 188352
rect 470600 188300 470652 188352
rect 106188 187688 106240 187740
rect 189816 187688 189868 187740
rect 236644 187144 236696 187196
rect 332692 187144 332744 187196
rect 41328 187076 41380 187128
rect 171508 187076 171560 187128
rect 203524 187076 203576 187128
rect 310612 187076 310664 187128
rect 164884 187008 164936 187060
rect 324688 187008 324740 187060
rect 339408 187008 339460 187060
rect 416872 187008 416924 187060
rect 147496 186940 147548 186992
rect 346492 186940 346544 186992
rect 417424 186940 417476 186992
rect 440240 186940 440292 186992
rect 134616 186396 134668 186448
rect 214564 186396 214616 186448
rect 114468 186328 114520 186380
rect 196624 186328 196676 186380
rect 321468 186260 321520 186312
rect 325884 186260 325936 186312
rect 189724 185784 189776 185836
rect 266544 185784 266596 185836
rect 152740 185716 152792 185768
rect 242348 185716 242400 185768
rect 120724 185648 120776 185700
rect 338304 185648 338356 185700
rect 80704 185580 80756 185632
rect 323216 185580 323268 185632
rect 365076 185580 365128 185632
rect 506480 185580 506532 185632
rect 100668 184900 100720 184952
rect 170404 184900 170456 184952
rect 221464 184356 221516 184408
rect 261116 184356 261168 184408
rect 140136 184288 140188 184340
rect 259644 184288 259696 184340
rect 48964 184220 49016 184272
rect 109684 184220 109736 184272
rect 125048 184220 125100 184272
rect 341064 184220 341116 184272
rect 103428 184152 103480 184204
rect 321284 184152 321336 184204
rect 327080 184152 327132 184204
rect 334164 184152 334216 184204
rect 480260 184152 480312 184204
rect 124128 183540 124180 183592
rect 169208 183540 169260 183592
rect 211896 183132 211948 183184
rect 265164 183132 265216 183184
rect 173164 183064 173216 183116
rect 249892 183064 249944 183116
rect 319536 183064 319588 183116
rect 330024 183064 330076 183116
rect 154488 182996 154540 183048
rect 338212 182996 338264 183048
rect 157984 182928 158036 182980
rect 345112 182928 345164 182980
rect 60556 182860 60608 182912
rect 272064 182860 272116 182912
rect 315396 182860 315448 182912
rect 339684 182860 339736 182912
rect 75184 182792 75236 182844
rect 321652 182792 321704 182844
rect 389824 182792 389876 182844
rect 436284 182792 436336 182844
rect 127808 182180 127860 182232
rect 167920 182180 167972 182232
rect 309048 182180 309100 182232
rect 339592 182180 339644 182232
rect 122104 182112 122156 182164
rect 269764 181840 269816 181892
rect 270408 181840 270460 181892
rect 222844 181500 222896 181552
rect 266452 181500 266504 181552
rect 156696 181432 156748 181484
rect 276112 181432 276164 181484
rect 392676 181432 392728 181484
rect 487160 181432 487212 181484
rect 121184 180888 121236 180940
rect 169300 180888 169352 180940
rect 112628 180820 112680 180872
rect 167736 180820 167788 180872
rect 269764 180820 269816 180872
rect 431316 180820 431368 180872
rect 242164 180412 242216 180464
rect 259736 180412 259788 180464
rect 236736 180344 236788 180396
rect 262404 180344 262456 180396
rect 313188 180344 313240 180396
rect 346676 180344 346728 180396
rect 237380 180276 237432 180328
rect 276664 180276 276716 180328
rect 300124 180276 300176 180328
rect 335452 180276 335504 180328
rect 215944 180208 215996 180260
rect 258356 180208 258408 180260
rect 304264 180208 304316 180260
rect 351368 180208 351420 180260
rect 210516 180140 210568 180192
rect 245660 180140 245712 180192
rect 257344 180140 257396 180192
rect 349344 180140 349396 180192
rect 169116 180072 169168 180124
rect 324504 180072 324556 180124
rect 403624 180072 403676 180124
rect 427820 180072 427872 180124
rect 124956 179664 125008 179716
rect 166448 179664 166500 179716
rect 115848 179596 115900 179648
rect 167828 179596 167880 179648
rect 116952 179528 117004 179580
rect 173164 179528 173216 179580
rect 148232 179460 148284 179512
rect 214656 179460 214708 179512
rect 110052 179392 110104 179444
rect 211896 179392 211948 179444
rect 285588 179392 285640 179444
rect 393964 179392 394016 179444
rect 185584 179324 185636 179376
rect 336832 179324 336884 179376
rect 246396 178848 246448 178900
rect 249340 178848 249392 178900
rect 229744 178780 229796 178832
rect 246948 178780 247000 178832
rect 247960 178780 248012 178832
rect 249064 178780 249116 178832
rect 216588 178712 216640 178764
rect 224960 178712 225012 178764
rect 240784 178712 240836 178764
rect 262220 178712 262272 178764
rect 220084 178644 220136 178696
rect 256884 178644 256936 178696
rect 279424 178644 279476 178696
rect 334072 178644 334124 178696
rect 348424 178644 348476 178696
rect 445852 178644 445904 178696
rect 132040 178372 132092 178424
rect 165252 178372 165304 178424
rect 159272 178304 159324 178356
rect 206376 178304 206428 178356
rect 118424 178236 118476 178288
rect 166356 178236 166408 178288
rect 99196 178168 99248 178220
rect 171784 178168 171836 178220
rect 130752 178100 130804 178152
rect 214104 178100 214156 178152
rect 308404 178100 308456 178152
rect 316040 178100 316092 178152
rect 125784 178032 125836 178084
rect 214932 178032 214984 178084
rect 309692 178032 309744 178084
rect 331496 178032 331548 178084
rect 464344 178032 464396 178084
rect 580172 178032 580224 178084
rect 97816 177964 97868 178016
rect 134616 177964 134668 178016
rect 166264 177964 166316 178016
rect 247684 177896 247736 177948
rect 249248 177896 249300 177948
rect 316684 177556 316736 177608
rect 325792 177556 325844 177608
rect 239496 177488 239548 177540
rect 250076 177488 250128 177540
rect 320088 177488 320140 177540
rect 329932 177488 329984 177540
rect 242256 177420 242308 177472
rect 258264 177420 258316 177472
rect 318064 177420 318116 177472
rect 332876 177420 332928 177472
rect 239588 177352 239640 177404
rect 256792 177352 256844 177404
rect 309968 177352 310020 177404
rect 329196 177352 329248 177404
rect 167644 177284 167696 177336
rect 251456 177284 251508 177336
rect 299296 177284 299348 177336
rect 311164 177284 311216 177336
rect 318708 177284 318760 177336
rect 342352 177284 342404 177336
rect 134432 176876 134484 176928
rect 164516 176876 164568 176928
rect 128176 176808 128228 176860
rect 167000 176808 167052 176860
rect 108120 176740 108172 176792
rect 169024 176740 169076 176792
rect 309784 176740 309836 176792
rect 313280 176740 313332 176792
rect 344284 176740 344336 176792
rect 429200 176740 429252 176792
rect 100760 176672 100812 176724
rect 171876 176672 171928 176724
rect 295340 176672 295392 176724
rect 296628 176672 296680 176724
rect 444564 176672 444616 176724
rect 135720 176604 135772 176656
rect 213920 176604 213972 176656
rect 233884 176604 233936 176656
rect 261208 176604 261260 176656
rect 287704 176604 287756 176656
rect 321468 176604 321520 176656
rect 242348 176536 242400 176588
rect 249156 176536 249208 176588
rect 319444 176468 319496 176520
rect 327080 176468 327132 176520
rect 133144 176196 133196 176248
rect 165528 176196 165580 176248
rect 129464 176128 129516 176180
rect 166172 176128 166224 176180
rect 121920 176060 121972 176112
rect 166264 176060 166316 176112
rect 321376 176060 321428 176112
rect 321744 176060 321796 176112
rect 396724 176060 396776 176112
rect 409972 176060 410024 176112
rect 104624 175992 104676 176044
rect 170496 175992 170548 176044
rect 266268 175992 266320 176044
rect 428464 175992 428516 176044
rect 8944 175924 8996 175976
rect 111064 175924 111116 175976
rect 119436 175924 119488 175976
rect 170588 175924 170640 175976
rect 247776 175924 247828 175976
rect 255504 175924 255556 175976
rect 278044 175924 278096 175976
rect 295340 175924 295392 175976
rect 297364 175924 297416 175976
rect 307668 175924 307720 175976
rect 313924 175924 313976 175976
rect 347964 175924 348016 175976
rect 553400 175924 553452 175976
rect 165528 175176 165580 175228
rect 214012 175176 214064 175228
rect 164516 175108 164568 175160
rect 213920 175108 213972 175160
rect 3240 164160 3292 164212
rect 57244 164160 57296 164212
rect 3424 150356 3476 150408
rect 13084 150356 13136 150408
rect 3240 137912 3292 137964
rect 18604 137912 18656 137964
rect 63408 126964 63460 127016
rect 65524 126964 65576 127016
rect 62028 121456 62080 121508
rect 66076 121456 66128 121508
rect 3424 111528 3476 111580
rect 8944 111528 8996 111580
rect 3424 97928 3476 97980
rect 14464 97928 14516 97980
rect 287704 174020 287756 174072
rect 307484 174020 307536 174072
rect 279424 173952 279476 174004
rect 307576 173952 307628 174004
rect 264244 173884 264296 173936
rect 307668 173884 307720 173936
rect 165252 173816 165304 173868
rect 213920 173816 213972 173868
rect 340144 173136 340196 173188
rect 516140 173136 516192 173188
rect 290648 172660 290700 172712
rect 307300 172660 307352 172712
rect 287796 172592 287848 172644
rect 307668 172592 307720 172644
rect 271236 172524 271288 172576
rect 306932 172524 306984 172576
rect 166172 172456 166224 172508
rect 213920 172456 213972 172508
rect 167000 172388 167052 172440
rect 214012 172388 214064 172440
rect 324320 172388 324372 172440
rect 327080 172388 327132 172440
rect 384304 171776 384356 171828
rect 450084 171776 450136 171828
rect 321744 171368 321796 171420
rect 325792 171368 325844 171420
rect 300124 171232 300176 171284
rect 307484 171232 307536 171284
rect 282368 171164 282420 171216
rect 307576 171164 307628 171216
rect 168012 171096 168064 171148
rect 211804 171096 211856 171148
rect 269948 171096 270000 171148
rect 307668 171096 307720 171148
rect 167920 171028 167972 171080
rect 213920 171028 213972 171080
rect 324320 171028 324372 171080
rect 349896 171028 349948 171080
rect 351368 171028 351420 171080
rect 498844 171028 498896 171080
rect 252468 170620 252520 170672
rect 256976 170620 257028 170672
rect 389088 170348 389140 170400
rect 422760 170348 422812 170400
rect 274088 169872 274140 169924
rect 307668 169872 307720 169924
rect 268476 169804 268528 169856
rect 306564 169804 306616 169856
rect 257528 169736 257580 169788
rect 307668 169736 307720 169788
rect 166448 169668 166500 169720
rect 213920 169668 213972 169720
rect 324320 169668 324372 169720
rect 369124 169668 369176 169720
rect 169208 169600 169260 169652
rect 214012 169600 214064 169652
rect 324412 169600 324464 169652
rect 328460 169600 328512 169652
rect 252376 169532 252428 169584
rect 263784 169532 263836 169584
rect 252468 169464 252520 169516
rect 258172 169464 258224 169516
rect 401600 169056 401652 169108
rect 422300 169056 422352 169108
rect 265624 168988 265676 169040
rect 307300 168988 307352 169040
rect 407764 168988 407816 169040
rect 539600 168988 539652 169040
rect 304264 168444 304316 168496
rect 306564 168444 306616 168496
rect 284944 168376 284996 168428
rect 307668 168376 307720 168428
rect 327816 168376 327868 168428
rect 334164 168376 334216 168428
rect 166264 168308 166316 168360
rect 213920 168308 213972 168360
rect 252376 168308 252428 168360
rect 263692 168308 263744 168360
rect 169300 168240 169352 168292
rect 214012 168240 214064 168292
rect 252468 168240 252520 168292
rect 262312 168240 262364 168292
rect 337292 168172 337344 168224
rect 339500 168172 339552 168224
rect 252008 167696 252060 167748
rect 256884 167696 256936 167748
rect 415400 167628 415452 167680
rect 440332 167628 440384 167680
rect 295984 167152 296036 167204
rect 307668 167152 307720 167204
rect 267096 167084 267148 167136
rect 307484 167084 307536 167136
rect 264336 167016 264388 167068
rect 307576 167016 307628 167068
rect 166356 166948 166408 167000
rect 214104 166948 214156 167000
rect 252376 166948 252428 167000
rect 261024 166948 261076 167000
rect 170588 166880 170640 166932
rect 213920 166880 213972 166932
rect 173164 166812 173216 166864
rect 214012 166812 214064 166864
rect 251916 166268 251968 166320
rect 256792 166268 256844 166320
rect 412640 166268 412692 166320
rect 435364 166268 435416 166320
rect 449164 166268 449216 166320
rect 476212 166268 476264 166320
rect 252468 165860 252520 165912
rect 259736 165860 259788 165912
rect 293224 165724 293276 165776
rect 306380 165724 306432 165776
rect 273996 165656 274048 165708
rect 306564 165656 306616 165708
rect 257620 165588 257672 165640
rect 306472 165588 306524 165640
rect 476212 165588 476264 165640
rect 580172 165588 580224 165640
rect 167828 165520 167880 165572
rect 213920 165520 213972 165572
rect 251916 165520 251968 165572
rect 267832 165520 267884 165572
rect 324320 165520 324372 165572
rect 337292 165520 337344 165572
rect 251456 165180 251508 165232
rect 252836 165180 252888 165232
rect 252468 164908 252520 164960
rect 258356 164908 258408 164960
rect 268384 164840 268436 164892
rect 307300 164840 307352 164892
rect 337936 164840 337988 164892
rect 426532 164840 426584 164892
rect 275376 164296 275428 164348
rect 306472 164432 306524 164484
rect 258908 164228 258960 164280
rect 306380 164364 306432 164416
rect 300308 164228 300360 164280
rect 306380 164228 306432 164280
rect 167736 164160 167788 164212
rect 214012 164160 214064 164212
rect 252192 164160 252244 164212
rect 266544 164160 266596 164212
rect 324412 164160 324464 164212
rect 331220 164160 331272 164212
rect 196624 164092 196676 164144
rect 213920 164092 213972 164144
rect 251916 164092 251968 164144
rect 265164 164092 265216 164144
rect 324320 164024 324372 164076
rect 327172 164024 327224 164076
rect 332416 163480 332468 163532
rect 340972 163480 341024 163532
rect 410524 163480 410576 163532
rect 443644 163480 443696 163532
rect 283564 163004 283616 163056
rect 306380 163004 306432 163056
rect 263048 162936 263100 162988
rect 306564 162936 306616 162988
rect 253296 162868 253348 162920
rect 306472 162868 306524 162920
rect 211896 162800 211948 162852
rect 213920 162800 213972 162852
rect 252468 162800 252520 162852
rect 262404 162800 262456 162852
rect 252100 162732 252152 162784
rect 261116 162732 261168 162784
rect 439596 162120 439648 162172
rect 447140 162120 447192 162172
rect 287888 161576 287940 161628
rect 306472 161576 306524 161628
rect 252468 161508 252520 161560
rect 259552 161508 259604 161560
rect 264612 161508 264664 161560
rect 306380 161508 306432 161560
rect 254584 161440 254636 161492
rect 306564 161440 306616 161492
rect 169024 161372 169076 161424
rect 213920 161372 213972 161424
rect 324320 161372 324372 161424
rect 335636 161372 335688 161424
rect 189908 161304 189960 161356
rect 214012 161304 214064 161356
rect 251364 160828 251416 160880
rect 254124 160828 254176 160880
rect 252468 160692 252520 160744
rect 258264 160692 258316 160744
rect 326436 160692 326488 160744
rect 338304 160692 338356 160744
rect 398656 160692 398708 160744
rect 536840 160692 536892 160744
rect 251916 160352 251968 160404
rect 255504 160352 255556 160404
rect 302976 160216 303028 160268
rect 306564 160216 306616 160268
rect 280896 160148 280948 160200
rect 306472 160148 306524 160200
rect 261576 160080 261628 160132
rect 306380 160080 306432 160132
rect 170496 160012 170548 160064
rect 214012 160012 214064 160064
rect 324320 160012 324372 160064
rect 332416 160012 332468 160064
rect 189816 159944 189868 159996
rect 213920 159944 213972 159996
rect 424324 159400 424376 159452
rect 449072 159400 449124 159452
rect 171876 159332 171928 159384
rect 214104 159332 214156 159384
rect 376116 159332 376168 159384
rect 455604 159332 455656 159384
rect 292212 158856 292264 158908
rect 306380 158856 306432 158908
rect 272524 158788 272576 158840
rect 306564 158788 306616 158840
rect 260288 158720 260340 158772
rect 306472 158720 306524 158772
rect 252376 158652 252428 158704
rect 272064 158652 272116 158704
rect 324412 158652 324464 158704
rect 334072 158652 334124 158704
rect 252468 158584 252520 158636
rect 265072 158584 265124 158636
rect 324320 158584 324372 158636
rect 330024 158584 330076 158636
rect 293408 157496 293460 157548
rect 306380 157496 306432 157548
rect 262864 157428 262916 157480
rect 306564 157428 306616 157480
rect 257344 157360 257396 157412
rect 306472 157360 306524 157412
rect 170404 157292 170456 157344
rect 213920 157292 213972 157344
rect 252468 157292 252520 157344
rect 267924 157292 267976 157344
rect 324412 157292 324464 157344
rect 332876 157292 332928 157344
rect 324320 157020 324372 157072
rect 325976 157020 326028 157072
rect 411904 156612 411956 156664
rect 449256 156612 449308 156664
rect 285128 156068 285180 156120
rect 307668 156068 307720 156120
rect 259000 156000 259052 156052
rect 307484 156000 307536 156052
rect 258816 155932 258868 155984
rect 307576 155932 307628 155984
rect 171784 155864 171836 155916
rect 213920 155864 213972 155916
rect 252468 155864 252520 155916
rect 278872 155864 278924 155916
rect 324320 155864 324372 155916
rect 356060 155864 356112 155916
rect 252376 155796 252428 155848
rect 274640 155796 274692 155848
rect 252468 155728 252520 155780
rect 264980 155728 265032 155780
rect 261668 155184 261720 155236
rect 306932 155184 306984 155236
rect 351276 155184 351328 155236
rect 451556 155184 451608 155236
rect 279516 154640 279568 154692
rect 307484 154640 307536 154692
rect 262956 154572 263008 154624
rect 306748 154572 306800 154624
rect 251732 154504 251784 154556
rect 277492 154504 277544 154556
rect 324320 154300 324372 154352
rect 326436 154300 326488 154352
rect 251180 154232 251232 154284
rect 254032 154232 254084 154284
rect 254768 153824 254820 153876
rect 307392 153824 307444 153876
rect 408408 153824 408460 153876
rect 426624 153824 426676 153876
rect 195244 153280 195296 153332
rect 214012 153280 214064 153332
rect 301504 153280 301556 153332
rect 307576 153280 307628 153332
rect 185584 153212 185636 153264
rect 213920 153212 213972 153264
rect 271144 153212 271196 153264
rect 307668 153212 307720 153264
rect 329196 153212 329248 153264
rect 431592 153280 431644 153332
rect 429660 153212 429712 153264
rect 431960 153212 432012 153264
rect 252008 153144 252060 153196
rect 271972 153144 272024 153196
rect 324320 153144 324372 153196
rect 339684 153144 339736 153196
rect 252468 153076 252520 153128
rect 269212 153076 269264 153128
rect 398932 152600 398984 152652
rect 420184 152600 420236 152652
rect 375196 152532 375248 152584
rect 418712 152532 418764 152584
rect 425796 152532 425848 152584
rect 455420 152532 455472 152584
rect 257436 152464 257488 152516
rect 307484 152464 307536 152516
rect 338764 152464 338816 152516
rect 400220 152464 400272 152516
rect 405648 152464 405700 152516
rect 456892 152464 456944 152516
rect 458824 152464 458876 152516
rect 580172 152464 580224 152516
rect 204904 151920 204956 151972
rect 213920 151920 213972 151972
rect 257712 151920 257764 151972
rect 306564 151920 306616 151972
rect 191104 151852 191156 151904
rect 214012 151852 214064 151904
rect 278136 151852 278188 151904
rect 307668 151852 307720 151904
rect 189816 151784 189868 151836
rect 213920 151784 213972 151836
rect 324320 151716 324372 151768
rect 341064 151716 341116 151768
rect 343824 151716 343876 151768
rect 535552 151716 535604 151768
rect 252468 151648 252520 151700
rect 270500 151648 270552 151700
rect 252376 151580 252428 151632
rect 273260 151580 273312 151632
rect 324320 151308 324372 151360
rect 327356 151308 327408 151360
rect 365628 151104 365680 151156
rect 406476 151104 406528 151156
rect 182088 151036 182140 151088
rect 206284 151036 206336 151088
rect 363696 151036 363748 151088
rect 412272 151036 412324 151088
rect 289360 150560 289412 150612
rect 307484 150560 307536 150612
rect 196716 150492 196768 150544
rect 213920 150492 213972 150544
rect 273904 150492 273956 150544
rect 307300 150492 307352 150544
rect 194048 150424 194100 150476
rect 214012 150424 214064 150476
rect 256148 150424 256200 150476
rect 307668 150424 307720 150476
rect 211804 150356 211856 150408
rect 213920 150356 213972 150408
rect 251916 150356 251968 150408
rect 281632 150356 281684 150408
rect 251548 150288 251600 150340
rect 255412 150288 255464 150340
rect 252652 149744 252704 149796
rect 262220 149744 262272 149796
rect 379428 149744 379480 149796
rect 397552 149744 397604 149796
rect 254860 149676 254912 149728
rect 306656 149676 306708 149728
rect 387248 149676 387300 149728
rect 454224 149676 454276 149728
rect 272616 149200 272668 149252
rect 307484 149200 307536 149252
rect 296260 149132 296312 149184
rect 307668 149132 307720 149184
rect 355324 149064 355376 149116
rect 420276 149064 420328 149116
rect 206376 148996 206428 149048
rect 213920 148996 213972 149048
rect 252468 148996 252520 149048
rect 276020 148996 276072 149048
rect 324412 148996 324464 149048
rect 352012 148996 352064 149048
rect 371884 148996 371936 149048
rect 435456 148996 435508 149048
rect 442724 148996 442776 149048
rect 324320 148928 324372 148980
rect 329932 148928 329984 148980
rect 431316 148724 431368 148776
rect 434168 148724 434220 148776
rect 409880 148520 409932 148572
rect 410708 148520 410760 148572
rect 426440 148520 426492 148572
rect 427452 148520 427504 148572
rect 446496 148520 446548 148572
rect 449624 148520 449676 148572
rect 387248 148384 387300 148436
rect 419448 148452 419500 148504
rect 421288 148452 421340 148504
rect 428464 148384 428516 148436
rect 435456 148384 435508 148436
rect 252008 148316 252060 148368
rect 273996 148316 274048 148368
rect 360016 148316 360068 148368
rect 400036 148316 400088 148368
rect 425152 148316 425204 148368
rect 436744 148316 436796 148368
rect 466552 148316 466604 148368
rect 522304 148316 522356 148368
rect 435548 148248 435600 148300
rect 438032 148248 438084 148300
rect 436100 148180 436152 148232
rect 443000 148180 443052 148232
rect 438676 148112 438728 148164
rect 439596 148112 439648 148164
rect 402612 147976 402664 148028
rect 403624 147976 403676 148028
rect 443644 147976 443696 148028
rect 446036 147976 446088 148028
rect 274180 147772 274232 147824
rect 307484 147772 307536 147824
rect 396816 147772 396868 147824
rect 405832 147772 405884 147824
rect 441896 147772 441948 147824
rect 442724 147772 442776 147824
rect 455972 147772 456024 147824
rect 271328 147704 271380 147756
rect 307576 147704 307628 147756
rect 377404 147704 377456 147756
rect 418896 147704 418948 147756
rect 448980 147704 449032 147756
rect 466552 147704 466604 147756
rect 260380 147636 260432 147688
rect 307668 147636 307720 147688
rect 373356 147636 373408 147688
rect 416872 147636 416924 147688
rect 429108 147636 429160 147688
rect 456064 147636 456116 147688
rect 339408 147568 339460 147620
rect 421564 147568 421616 147620
rect 421932 147568 421984 147620
rect 446404 147568 446456 147620
rect 451556 147568 451608 147620
rect 252376 147500 252428 147552
rect 276112 147500 276164 147552
rect 324320 147500 324372 147552
rect 345112 147500 345164 147552
rect 252468 147432 252520 147484
rect 277400 147432 277452 147484
rect 251180 146956 251232 147008
rect 253940 146956 253992 147008
rect 392584 146956 392636 147008
rect 400128 146956 400180 147008
rect 447784 146956 447836 147008
rect 459560 146956 459612 147008
rect 251548 146888 251600 146940
rect 263600 146888 263652 146940
rect 327724 146888 327776 146940
rect 338212 146888 338264 146940
rect 339408 146888 339460 146940
rect 395804 146888 395856 146940
rect 402980 146888 403032 146940
rect 431224 146888 431276 146940
rect 454316 146888 454368 146940
rect 381544 146412 381596 146464
rect 407764 146412 407816 146464
rect 304540 146344 304592 146396
rect 307484 146344 307536 146396
rect 331864 146344 331916 146396
rect 432604 146344 432656 146396
rect 433524 146344 433576 146396
rect 433984 146344 434036 146396
rect 460204 146344 460256 146396
rect 188344 146276 188396 146328
rect 213920 146276 213972 146328
rect 254676 146276 254728 146328
rect 307668 146276 307720 146328
rect 400128 146276 400180 146328
rect 580356 146276 580408 146328
rect 251732 146208 251784 146260
rect 259644 146208 259696 146260
rect 324320 146208 324372 146260
rect 346676 146208 346728 146260
rect 251916 146140 251968 146192
rect 266452 146140 266504 146192
rect 324412 146140 324464 146192
rect 331312 146140 331364 146192
rect 252100 146072 252152 146124
rect 270592 146072 270644 146124
rect 446772 145936 446824 145988
rect 449256 145936 449308 145988
rect 252008 145596 252060 145648
rect 268476 145596 268528 145648
rect 253388 145528 253440 145580
rect 307024 145528 307076 145580
rect 369124 145528 369176 145580
rect 423588 145528 423640 145580
rect 456064 145528 456116 145580
rect 580264 145528 580316 145580
rect 399852 145392 399904 145444
rect 403532 145392 403584 145444
rect 359464 145052 359516 145104
rect 397460 145052 397512 145104
rect 171784 144984 171836 145036
rect 213920 144984 213972 145036
rect 287980 144984 288032 145036
rect 307484 144984 307536 145036
rect 378876 144984 378928 145036
rect 417056 145392 417108 145444
rect 166264 144916 166316 144968
rect 214012 144916 214064 144968
rect 268568 144916 268620 144968
rect 307668 144916 307720 144968
rect 329196 144916 329248 144968
rect 399852 144916 399904 144968
rect 252192 144848 252244 144900
rect 267740 144848 267792 144900
rect 324412 144848 324464 144900
rect 331496 144848 331548 144900
rect 452568 144848 452620 144900
rect 467104 144848 467156 144900
rect 324320 144780 324372 144832
rect 328552 144780 328604 144832
rect 294696 144236 294748 144288
rect 307576 144236 307628 144288
rect 373264 144236 373316 144288
rect 376668 144236 376720 144288
rect 397460 144236 397512 144288
rect 264520 144168 264572 144220
rect 306564 144168 306616 144220
rect 340972 144168 341024 144220
rect 400496 144168 400548 144220
rect 252468 144032 252520 144084
rect 258080 144032 258132 144084
rect 192576 143556 192628 143608
rect 213920 143556 213972 143608
rect 293500 143556 293552 143608
rect 307484 143556 307536 143608
rect 324964 143556 325016 143608
rect 327816 143556 327868 143608
rect 252468 143488 252520 143540
rect 260932 143488 260984 143540
rect 324320 143488 324372 143540
rect 331404 143488 331456 143540
rect 449072 143420 449124 143472
rect 449532 143420 449584 143472
rect 211804 142672 211856 142724
rect 213920 142672 213972 142724
rect 251824 142672 251876 142724
rect 257344 142672 257396 142724
rect 279608 142196 279660 142248
rect 307484 142196 307536 142248
rect 189724 142128 189776 142180
rect 213920 142128 213972 142180
rect 255964 142128 256016 142180
rect 307668 142128 307720 142180
rect 331956 142128 332008 142180
rect 397552 142128 397604 142180
rect 452476 142128 452528 142180
rect 498844 142128 498896 142180
rect 251732 142060 251784 142112
rect 259460 142060 259512 142112
rect 324412 142060 324464 142112
rect 332784 142060 332836 142112
rect 365168 142060 365220 142112
rect 397460 142060 397512 142112
rect 324320 141788 324372 141840
rect 327264 141788 327316 141840
rect 252376 141380 252428 141432
rect 264244 141380 264296 141432
rect 301688 140904 301740 140956
rect 307668 140904 307720 140956
rect 206376 140836 206428 140888
rect 213920 140836 213972 140888
rect 290556 140836 290608 140888
rect 307576 140836 307628 140888
rect 196624 140768 196676 140820
rect 214012 140768 214064 140820
rect 257620 140768 257672 140820
rect 307668 140768 307720 140820
rect 343824 140768 343876 140820
rect 346400 140768 346452 140820
rect 324320 140700 324372 140752
rect 337476 140700 337528 140752
rect 451924 140428 451976 140480
rect 455604 140428 455656 140480
rect 194508 140020 194560 140072
rect 215944 140020 215996 140072
rect 335636 140020 335688 140072
rect 376668 140020 376720 140072
rect 286324 139544 286376 139596
rect 306564 139544 306616 139596
rect 251732 139476 251784 139528
rect 255596 139476 255648 139528
rect 256056 139476 256108 139528
rect 307576 139476 307628 139528
rect 182916 139408 182968 139460
rect 213920 139408 213972 139460
rect 250536 139408 250588 139460
rect 307668 139408 307720 139460
rect 251732 139340 251784 139392
rect 280160 139340 280212 139392
rect 354036 139340 354088 139392
rect 354680 139340 354732 139392
rect 397460 139340 397512 139392
rect 252468 139272 252520 139324
rect 260840 139272 260892 139324
rect 324320 139272 324372 139324
rect 354864 139272 354916 139324
rect 452108 138864 452160 138916
rect 458364 138864 458416 138916
rect 282276 138116 282328 138168
rect 307668 138116 307720 138168
rect 253204 138048 253256 138100
rect 307484 138048 307536 138100
rect 193956 137980 194008 138032
rect 213920 137980 213972 138032
rect 250444 137980 250496 138032
rect 307576 137980 307628 138032
rect 252468 137912 252520 137964
rect 281540 137912 281592 137964
rect 324320 137912 324372 137964
rect 347964 137912 348016 137964
rect 360108 137912 360160 137964
rect 397552 137912 397604 137964
rect 251364 137844 251416 137896
rect 269120 137844 269172 137896
rect 322940 137844 322992 137896
rect 323308 137844 323360 137896
rect 330484 137844 330536 137896
rect 391848 137844 391900 137896
rect 397460 137844 397512 137896
rect 256240 137232 256292 137284
rect 307116 137232 307168 137284
rect 210516 136688 210568 136740
rect 213920 136688 213972 136740
rect 293316 136688 293368 136740
rect 306748 136688 306800 136740
rect 171876 136620 171928 136672
rect 214104 136620 214156 136672
rect 276756 136620 276808 136672
rect 307668 136620 307720 136672
rect 252468 136552 252520 136604
rect 287704 136552 287756 136604
rect 323400 136552 323452 136604
rect 343824 136552 343876 136604
rect 251732 136484 251784 136536
rect 279424 136484 279476 136536
rect 324320 136484 324372 136536
rect 342444 136484 342496 136536
rect 300216 135464 300268 135516
rect 307668 135464 307720 135516
rect 207756 135396 207808 135448
rect 214012 135396 214064 135448
rect 298744 135396 298796 135448
rect 306932 135396 306984 135448
rect 202236 135328 202288 135380
rect 213920 135328 213972 135380
rect 280804 135328 280856 135380
rect 306564 135328 306616 135380
rect 181444 135260 181496 135312
rect 214104 135260 214156 135312
rect 267004 135260 267056 135312
rect 306748 135260 306800 135312
rect 390192 135260 390244 135312
rect 391940 135260 391992 135312
rect 397460 135260 397512 135312
rect 251456 135192 251508 135244
rect 287796 135192 287848 135244
rect 324412 135192 324464 135244
rect 335452 135192 335504 135244
rect 451924 135192 451976 135244
rect 454316 135192 454368 135244
rect 252468 135124 252520 135176
rect 271236 135124 271288 135176
rect 324320 135124 324372 135176
rect 332692 135124 332744 135176
rect 394056 134648 394108 134700
rect 396080 134648 396132 134700
rect 397460 134648 397512 134700
rect 327080 134512 327132 134564
rect 367100 134512 367152 134564
rect 387156 134512 387208 134564
rect 399024 134512 399076 134564
rect 296076 134036 296128 134088
rect 307668 134036 307720 134088
rect 174636 133968 174688 134020
rect 214012 133968 214064 134020
rect 290464 133968 290516 134020
rect 307484 133968 307536 134020
rect 170404 133900 170456 133952
rect 213920 133900 213972 133952
rect 289268 133900 289320 133952
rect 307576 133900 307628 133952
rect 251364 133832 251416 133884
rect 290648 133832 290700 133884
rect 324320 133832 324372 133884
rect 357532 133832 357584 133884
rect 452200 133832 452252 133884
rect 482284 133832 482336 133884
rect 252376 133764 252428 133816
rect 282368 133764 282420 133816
rect 252468 133696 252520 133748
rect 269948 133696 270000 133748
rect 321652 133152 321704 133204
rect 357440 133152 357492 133204
rect 297456 132608 297508 132660
rect 307668 132608 307720 132660
rect 207664 132540 207716 132592
rect 214012 132540 214064 132592
rect 282460 132540 282512 132592
rect 307484 132540 307536 132592
rect 391296 132540 391348 132592
rect 394608 132540 394660 132592
rect 397552 132540 397604 132592
rect 173164 132472 173216 132524
rect 213920 132472 213972 132524
rect 269856 132472 269908 132524
rect 307576 132472 307628 132524
rect 392584 132472 392636 132524
rect 397460 132472 397512 132524
rect 252468 132404 252520 132456
rect 300124 132404 300176 132456
rect 449992 132404 450044 132456
rect 472624 132404 472676 132456
rect 251548 132336 251600 132388
rect 265624 132336 265676 132388
rect 252008 131792 252060 131844
rect 279516 131792 279568 131844
rect 265716 131724 265768 131776
rect 301504 131724 301556 131776
rect 337476 131724 337528 131776
rect 398748 131724 398800 131776
rect 303068 131248 303120 131300
rect 307484 131248 307536 131300
rect 287704 131180 287756 131232
rect 307576 131180 307628 131232
rect 264428 131112 264480 131164
rect 307668 131112 307720 131164
rect 252376 131044 252428 131096
rect 304264 131044 304316 131096
rect 324412 131044 324464 131096
rect 356244 131044 356296 131096
rect 360844 131044 360896 131096
rect 252468 130976 252520 131028
rect 274088 130976 274140 131028
rect 324320 130976 324372 131028
rect 339592 130976 339644 131028
rect 252468 130500 252520 130552
rect 257528 130500 257580 130552
rect 449164 130024 449216 130076
rect 449440 130024 449492 130076
rect 257344 129956 257396 130008
rect 307576 129956 307628 130008
rect 292028 129888 292080 129940
rect 307668 129888 307720 129940
rect 273996 129820 274048 129872
rect 307484 129820 307536 129872
rect 395896 129820 395948 129872
rect 398288 129820 398340 129872
rect 184204 129752 184256 129804
rect 213920 129752 213972 129804
rect 304356 129752 304408 129804
rect 307116 129752 307168 129804
rect 360936 129752 360988 129804
rect 397552 129752 397604 129804
rect 252468 129684 252520 129736
rect 284944 129684 284996 129736
rect 324412 129684 324464 129736
rect 343732 129684 343784 129736
rect 362224 129684 362276 129736
rect 385684 129684 385736 129736
rect 397460 129684 397512 129736
rect 452568 129684 452620 129736
rect 465080 129684 465132 129736
rect 251456 129616 251508 129668
rect 268384 129616 268436 129668
rect 252376 129548 252428 129600
rect 267096 129548 267148 129600
rect 324320 129412 324372 129464
rect 327080 129412 327132 129464
rect 285036 128392 285088 128444
rect 306564 128392 306616 128444
rect 186964 128324 187016 128376
rect 213920 128324 213972 128376
rect 268476 128324 268528 128376
rect 307116 128324 307168 128376
rect 251640 128256 251692 128308
rect 295984 128256 296036 128308
rect 324320 128256 324372 128308
rect 349344 128256 349396 128308
rect 392676 128256 392728 128308
rect 452108 128256 452160 128308
rect 458272 128256 458324 128308
rect 252468 128188 252520 128240
rect 264336 128188 264388 128240
rect 324412 128188 324464 128240
rect 329840 128188 329892 128240
rect 385684 127576 385736 127628
rect 397460 127576 397512 127628
rect 252192 127440 252244 127492
rect 257712 127440 257764 127492
rect 297548 127100 297600 127152
rect 307116 127100 307168 127152
rect 264244 127032 264296 127084
rect 307668 127032 307720 127084
rect 170496 126964 170548 127016
rect 213920 126964 213972 127016
rect 260196 126964 260248 127016
rect 306748 126964 306800 127016
rect 252468 126896 252520 126948
rect 293224 126896 293276 126948
rect 342996 126896 343048 126948
rect 343640 126896 343692 126948
rect 397552 126896 397604 126948
rect 452568 126896 452620 126948
rect 476212 126896 476264 126948
rect 252100 126828 252152 126880
rect 275376 126828 275428 126880
rect 377956 126828 378008 126880
rect 397460 126828 397512 126880
rect 251364 126216 251416 126268
rect 300308 126216 300360 126268
rect 203616 125672 203668 125724
rect 213920 125672 213972 125724
rect 284944 125672 284996 125724
rect 307668 125672 307720 125724
rect 200764 125604 200816 125656
rect 214012 125604 214064 125656
rect 275284 125604 275336 125656
rect 306748 125604 306800 125656
rect 324320 125536 324372 125588
rect 347872 125536 347924 125588
rect 353944 125536 353996 125588
rect 397460 125536 397512 125588
rect 452568 125536 452620 125588
rect 464344 125536 464396 125588
rect 251916 125332 251968 125384
rect 256240 125332 256292 125384
rect 252468 124992 252520 125044
rect 258908 124992 258960 125044
rect 252284 124856 252336 124908
rect 302976 124856 303028 124908
rect 451280 124720 451332 124772
rect 454224 124720 454276 124772
rect 302884 124312 302936 124364
rect 307668 124312 307720 124364
rect 171968 124244 172020 124296
rect 214012 124244 214064 124296
rect 291936 124244 291988 124296
rect 306748 124244 306800 124296
rect 167644 124176 167696 124228
rect 213920 124176 213972 124228
rect 258724 124176 258776 124228
rect 307116 124176 307168 124228
rect 252376 124108 252428 124160
rect 283564 124108 283616 124160
rect 252468 124040 252520 124092
rect 263048 124040 263100 124092
rect 251180 123496 251232 123548
rect 253296 123496 253348 123548
rect 338212 123428 338264 123480
rect 397368 123428 397420 123480
rect 395436 123224 395488 123276
rect 397460 123224 397512 123276
rect 300124 122952 300176 123004
rect 307116 122952 307168 123004
rect 183008 122884 183060 122936
rect 214012 122884 214064 122936
rect 289176 122884 289228 122936
rect 306564 122884 306616 122936
rect 166356 122816 166408 122868
rect 213920 122816 213972 122868
rect 260104 122816 260156 122868
rect 307668 122816 307720 122868
rect 252468 122748 252520 122800
rect 287888 122748 287940 122800
rect 324320 122748 324372 122800
rect 345020 122748 345072 122800
rect 252008 122680 252060 122732
rect 264612 122680 264664 122732
rect 452568 122612 452620 122664
rect 459560 122612 459612 122664
rect 251364 122476 251416 122528
rect 254584 122476 254636 122528
rect 395344 122272 395396 122324
rect 397460 122272 397512 122324
rect 287796 121592 287848 121644
rect 307668 121592 307720 121644
rect 189908 121524 189960 121576
rect 213920 121524 213972 121576
rect 283564 121524 283616 121576
rect 307484 121524 307536 121576
rect 169024 121456 169076 121508
rect 214012 121456 214064 121508
rect 264336 121456 264388 121508
rect 307576 121456 307628 121508
rect 252468 121388 252520 121440
rect 280896 121388 280948 121440
rect 324320 121388 324372 121440
rect 251824 121320 251876 121372
rect 261576 121320 261628 121372
rect 324412 121320 324464 121372
rect 338120 121320 338172 121372
rect 367008 121388 367060 121440
rect 397460 121388 397512 121440
rect 346584 121320 346636 121372
rect 370504 121320 370556 121372
rect 252376 120232 252428 120284
rect 259000 120232 259052 120284
rect 301504 120232 301556 120284
rect 306748 120232 306800 120284
rect 206468 120164 206520 120216
rect 214012 120164 214064 120216
rect 279516 120164 279568 120216
rect 307576 120164 307628 120216
rect 169300 120096 169352 120148
rect 213920 120096 213972 120148
rect 261484 120096 261536 120148
rect 307668 120096 307720 120148
rect 252468 120028 252520 120080
rect 292212 120028 292264 120080
rect 324320 120028 324372 120080
rect 346492 120028 346544 120080
rect 383016 120028 383068 120080
rect 397460 120028 397512 120080
rect 251364 119960 251416 120012
rect 272524 119960 272576 120012
rect 271420 119348 271472 119400
rect 307300 119348 307352 119400
rect 325056 119348 325108 119400
rect 333980 119348 334032 119400
rect 252284 119280 252336 119332
rect 260288 119280 260340 119332
rect 211896 118804 211948 118856
rect 214104 118804 214156 118856
rect 302976 118804 303028 118856
rect 307668 118804 307720 118856
rect 173348 118736 173400 118788
rect 213920 118736 213972 118788
rect 292120 118736 292172 118788
rect 307576 118736 307628 118788
rect 167736 118668 167788 118720
rect 214012 118668 214064 118720
rect 282368 118668 282420 118720
rect 307484 118668 307536 118720
rect 251824 118600 251876 118652
rect 293408 118600 293460 118652
rect 324320 118600 324372 118652
rect 354772 118600 354824 118652
rect 452476 118600 452528 118652
rect 484400 118600 484452 118652
rect 252468 118532 252520 118584
rect 262864 118532 262916 118584
rect 254584 117512 254636 117564
rect 307668 117512 307720 117564
rect 298836 117444 298888 117496
rect 306564 117444 306616 117496
rect 188436 117376 188488 117428
rect 214012 117376 214064 117428
rect 293224 117376 293276 117428
rect 307668 117376 307720 117428
rect 169208 117308 169260 117360
rect 213920 117308 213972 117360
rect 304448 117308 304500 117360
rect 307576 117308 307628 117360
rect 251364 117240 251416 117292
rect 261668 117240 261720 117292
rect 347228 117240 347280 117292
rect 365076 117240 365128 117292
rect 380164 117240 380216 117292
rect 397460 117240 397512 117292
rect 449348 117240 449400 117292
rect 503720 117240 503772 117292
rect 252468 117172 252520 117224
rect 258816 117172 258868 117224
rect 252008 116560 252060 116612
rect 305736 116560 305788 116612
rect 324320 116560 324372 116612
rect 347228 116560 347280 116612
rect 185676 116016 185728 116068
rect 213920 116016 213972 116068
rect 272524 116016 272576 116068
rect 306748 116016 306800 116068
rect 181536 115948 181588 116000
rect 214012 115948 214064 116000
rect 262864 115948 262916 116000
rect 307484 115948 307536 116000
rect 252284 115880 252336 115932
rect 285128 115880 285180 115932
rect 324320 115880 324372 115932
rect 342352 115880 342404 115932
rect 354588 115880 354640 115932
rect 397460 115880 397512 115932
rect 251916 115812 251968 115864
rect 262956 115812 263008 115864
rect 451556 115812 451608 115864
rect 455512 115812 455564 115864
rect 324964 115268 325016 115320
rect 332600 115268 332652 115320
rect 251824 115200 251876 115252
rect 268568 115200 268620 115252
rect 286416 115200 286468 115252
rect 307392 115200 307444 115252
rect 323584 115200 323636 115252
rect 337384 115200 337436 115252
rect 203708 114588 203760 114640
rect 214012 114588 214064 114640
rect 294604 114588 294656 114640
rect 307576 114588 307628 114640
rect 184296 114520 184348 114572
rect 213920 114520 213972 114572
rect 265624 114520 265676 114572
rect 307668 114520 307720 114572
rect 251364 114452 251416 114504
rect 265716 114452 265768 114504
rect 324320 114452 324372 114504
rect 358820 114452 358872 114504
rect 362868 114452 362920 114504
rect 397460 114452 397512 114504
rect 452476 114452 452528 114504
rect 485780 114452 485832 114504
rect 324412 114384 324464 114436
rect 351920 114384 351972 114436
rect 363604 114384 363656 114436
rect 251640 114180 251692 114232
rect 254768 114180 254820 114232
rect 252468 113772 252520 113824
rect 271144 113772 271196 113824
rect 360200 113772 360252 113824
rect 387156 113772 387208 113824
rect 295984 113296 296036 113348
rect 306564 113296 306616 113348
rect 198096 113228 198148 113280
rect 214012 113228 214064 113280
rect 279424 113228 279476 113280
rect 306932 113228 306984 113280
rect 173256 113160 173308 113212
rect 213920 113160 213972 113212
rect 268384 113160 268436 113212
rect 307668 113160 307720 113212
rect 395988 113092 396040 113144
rect 397460 113092 397512 113144
rect 456064 113092 456116 113144
rect 580172 113092 580224 113144
rect 252468 112820 252520 112872
rect 257436 112820 257488 112872
rect 252192 112480 252244 112532
rect 271328 112480 271380 112532
rect 257528 112412 257580 112464
rect 307208 112412 307260 112464
rect 251640 112208 251692 112260
rect 254860 112208 254912 112260
rect 202328 111868 202380 111920
rect 214012 111868 214064 111920
rect 301596 111868 301648 111920
rect 307668 111868 307720 111920
rect 169116 111800 169168 111852
rect 213920 111800 213972 111852
rect 271236 111800 271288 111852
rect 307484 111800 307536 111852
rect 168288 111732 168340 111784
rect 196716 111732 196768 111784
rect 387064 111732 387116 111784
rect 397460 111732 397512 111784
rect 452476 111732 452528 111784
rect 469220 111732 469272 111784
rect 390468 111664 390520 111716
rect 399576 111664 399628 111716
rect 452568 111664 452620 111716
rect 466460 111664 466512 111716
rect 251824 111256 251876 111308
rect 260380 111256 260432 111308
rect 252284 111052 252336 111104
rect 305644 111052 305696 111104
rect 345664 111052 345716 111104
rect 397552 111052 397604 111104
rect 304264 110576 304316 110628
rect 307484 110576 307536 110628
rect 263048 110508 263100 110560
rect 307576 110508 307628 110560
rect 173440 110440 173492 110492
rect 213920 110440 213972 110492
rect 253296 110440 253348 110492
rect 307668 110440 307720 110492
rect 167828 110372 167880 110424
rect 194048 110372 194100 110424
rect 251916 110372 251968 110424
rect 289360 110372 289412 110424
rect 324320 110372 324372 110424
rect 347780 110372 347832 110424
rect 378784 110372 378836 110424
rect 397460 110372 397512 110424
rect 252468 110304 252520 110356
rect 273904 110304 273956 110356
rect 452108 110304 452160 110356
rect 456892 110304 456944 110356
rect 252100 110236 252152 110288
rect 256148 110236 256200 110288
rect 300400 109148 300452 109200
rect 307484 109148 307536 109200
rect 174728 109080 174780 109132
rect 214012 109080 214064 109132
rect 275376 109080 275428 109132
rect 307576 109080 307628 109132
rect 170588 109012 170640 109064
rect 213920 109012 213972 109064
rect 258816 109012 258868 109064
rect 307668 109012 307720 109064
rect 395344 109012 395396 109064
rect 397736 109012 397788 109064
rect 168104 108944 168156 108996
rect 189816 108944 189868 108996
rect 252376 108944 252428 108996
rect 296260 108944 296312 108996
rect 324412 108944 324464 108996
rect 366364 108944 366416 108996
rect 252468 108876 252520 108928
rect 272616 108876 272668 108928
rect 324320 108876 324372 108928
rect 340144 108876 340196 108928
rect 249156 107856 249208 107908
rect 307668 107856 307720 107908
rect 296168 107788 296220 107840
rect 307576 107788 307628 107840
rect 170680 107720 170732 107772
rect 214012 107720 214064 107772
rect 273904 107720 273956 107772
rect 307668 107720 307720 107772
rect 166448 107652 166500 107704
rect 213920 107652 213972 107704
rect 363604 107652 363656 107704
rect 397460 107652 397512 107704
rect 252100 107584 252152 107636
rect 274180 107584 274232 107636
rect 323308 107584 323360 107636
rect 367744 107584 367796 107636
rect 252008 106904 252060 106956
rect 308404 106904 308456 106956
rect 376024 106904 376076 106956
rect 397644 106904 397696 106956
rect 274088 106428 274140 106480
rect 307668 106428 307720 106480
rect 204996 106360 205048 106412
rect 214012 106360 214064 106412
rect 285128 106360 285180 106412
rect 307576 106360 307628 106412
rect 194048 106292 194100 106344
rect 213920 106292 213972 106344
rect 252468 106224 252520 106276
rect 304540 106224 304592 106276
rect 324320 106224 324372 106276
rect 356152 106224 356204 106276
rect 363788 106224 363840 106276
rect 251916 106156 251968 106208
rect 294696 106156 294748 106208
rect 251364 106088 251416 106140
rect 254676 106088 254728 106140
rect 182824 105544 182876 105596
rect 216036 105544 216088 105596
rect 365076 105544 365128 105596
rect 397460 105544 397512 105596
rect 211988 105000 212040 105052
rect 213920 105000 213972 105052
rect 294788 105000 294840 105052
rect 307668 105000 307720 105052
rect 198188 104932 198240 104984
rect 214012 104932 214064 104984
rect 196808 104864 196860 104916
rect 213920 104864 213972 104916
rect 304632 104864 304684 104916
rect 307576 104864 307628 104916
rect 452568 104864 452620 104916
rect 454224 104864 454276 104916
rect 251916 104796 251968 104848
rect 308496 104796 308548 104848
rect 324320 104796 324372 104848
rect 335544 104796 335596 104848
rect 378968 104796 379020 104848
rect 397552 104796 397604 104848
rect 252468 104728 252520 104780
rect 287980 104728 288032 104780
rect 252284 104116 252336 104168
rect 293500 104116 293552 104168
rect 324504 104116 324556 104168
rect 329104 104116 329156 104168
rect 293408 103640 293460 103692
rect 307668 103640 307720 103692
rect 195336 103572 195388 103624
rect 214012 103572 214064 103624
rect 287888 103572 287940 103624
rect 307484 103572 307536 103624
rect 191196 103504 191248 103556
rect 213920 103504 213972 103556
rect 262956 103504 263008 103556
rect 307576 103504 307628 103556
rect 252468 103436 252520 103488
rect 286416 103436 286468 103488
rect 321652 103436 321704 103488
rect 374644 103436 374696 103488
rect 382096 103436 382148 103488
rect 397552 103436 397604 103488
rect 252008 103368 252060 103420
rect 264520 103368 264572 103420
rect 452568 103028 452620 103080
rect 454132 103028 454184 103080
rect 252376 102960 252428 103012
rect 257528 102960 257580 103012
rect 167920 102756 167972 102808
rect 214656 102756 214708 102808
rect 303528 102348 303580 102400
rect 308404 102348 308456 102400
rect 294696 102280 294748 102332
rect 307668 102280 307720 102332
rect 209044 102212 209096 102264
rect 214012 102212 214064 102264
rect 287980 102212 288032 102264
rect 307484 102212 307536 102264
rect 189816 102144 189868 102196
rect 213920 102144 213972 102196
rect 257436 102144 257488 102196
rect 307576 102144 307628 102196
rect 252468 102076 252520 102128
rect 271420 102076 271472 102128
rect 324320 102076 324372 102128
rect 351368 102076 351420 102128
rect 388444 102076 388496 102128
rect 397552 102076 397604 102128
rect 324412 102008 324464 102060
rect 335360 102008 335412 102060
rect 393228 102008 393280 102060
rect 397644 102008 397696 102060
rect 166540 101396 166592 101448
rect 214564 101396 214616 101448
rect 252100 101396 252152 101448
rect 297364 101396 297416 101448
rect 327080 101396 327132 101448
rect 394056 101396 394108 101448
rect 257528 100920 257580 100972
rect 307668 100920 307720 100972
rect 252008 100852 252060 100904
rect 255964 100852 256016 100904
rect 296260 100784 296312 100836
rect 307576 100784 307628 100836
rect 196716 100716 196768 100768
rect 213920 100716 213972 100768
rect 301780 100716 301832 100768
rect 306748 100716 306800 100768
rect 251732 100648 251784 100700
rect 301688 100648 301740 100700
rect 324320 100648 324372 100700
rect 345756 100648 345808 100700
rect 452568 100648 452620 100700
rect 477500 100648 477552 100700
rect 252468 100580 252520 100632
rect 279608 100580 279660 100632
rect 252376 100512 252428 100564
rect 270040 100512 270092 100564
rect 374644 99968 374696 100020
rect 397552 99968 397604 100020
rect 192668 99424 192720 99476
rect 213920 99424 213972 99476
rect 303160 99424 303212 99476
rect 307668 99424 307720 99476
rect 167828 99356 167880 99408
rect 214012 99356 214064 99408
rect 297364 99356 297416 99408
rect 307576 99356 307628 99408
rect 576124 99356 576176 99408
rect 580172 99356 580224 99408
rect 251548 99288 251600 99340
rect 257620 99288 257672 99340
rect 251824 99152 251876 99204
rect 290556 99152 290608 99204
rect 251180 99084 251232 99136
rect 253388 99084 253440 99136
rect 452292 98880 452344 98932
rect 454040 98880 454092 98932
rect 332600 98608 332652 98660
rect 391940 98608 391992 98660
rect 172060 98064 172112 98116
rect 214012 98064 214064 98116
rect 300308 98064 300360 98116
rect 307576 98064 307628 98116
rect 164884 97996 164936 98048
rect 213920 97996 213972 98048
rect 283656 97996 283708 98048
rect 307668 97996 307720 98048
rect 399024 97792 399076 97844
rect 399668 97792 399720 97844
rect 252192 97588 252244 97640
rect 256056 97588 256108 97640
rect 453304 97248 453356 97300
rect 467840 97248 467892 97300
rect 255964 96772 256016 96824
rect 307668 96772 307720 96824
rect 251916 96704 251968 96756
rect 307576 96704 307628 96756
rect 209136 96636 209188 96688
rect 213920 96636 213972 96688
rect 249064 96636 249116 96688
rect 307668 96636 307720 96688
rect 356796 96636 356848 96688
rect 397552 96636 397604 96688
rect 174544 96568 174596 96620
rect 321468 96568 321520 96620
rect 299296 95888 299348 95940
rect 314660 95888 314712 95940
rect 378048 95276 378100 95328
rect 419356 95276 419408 95328
rect 441896 95276 441948 95328
rect 460940 95276 460992 95328
rect 211160 95208 211212 95260
rect 213920 95208 213972 95260
rect 298928 95208 298980 95260
rect 307668 95208 307720 95260
rect 342904 95208 342956 95260
rect 400680 95208 400732 95260
rect 448980 95208 449032 95260
rect 480352 95208 480404 95260
rect 193864 95140 193916 95192
rect 322940 95140 322992 95192
rect 356704 95140 356756 95192
rect 422576 95140 422628 95192
rect 438676 95140 438728 95192
rect 525064 95140 525116 95192
rect 202144 95072 202196 95124
rect 321652 95072 321704 95124
rect 368296 95072 368348 95124
rect 447048 95072 447100 95124
rect 63408 95004 63460 95056
rect 196808 95004 196860 95056
rect 276664 95004 276716 95056
rect 325700 95004 325752 95056
rect 326344 95004 326396 95056
rect 371976 95004 372028 95056
rect 430948 95004 431000 95056
rect 438124 95004 438176 95056
rect 438676 95004 438728 95056
rect 438768 95004 438820 95056
rect 459652 95004 459704 95056
rect 436744 94936 436796 94988
rect 463700 94936 463752 94988
rect 425796 94868 425848 94920
rect 458824 94868 458876 94920
rect 395804 94800 395856 94852
rect 432236 94800 432288 94852
rect 438768 94800 438820 94852
rect 441252 94732 441304 94784
rect 317420 94460 317472 94512
rect 344284 94460 344336 94512
rect 115848 94052 115900 94104
rect 169300 94052 169352 94104
rect 113180 93984 113232 94036
rect 181444 93984 181496 94036
rect 126520 93916 126572 93968
rect 200764 93916 200816 93968
rect 94964 93848 95016 93900
rect 170680 93848 170732 93900
rect 66168 93780 66220 93832
rect 198188 93780 198240 93832
rect 308404 93780 308456 93832
rect 321744 93780 321796 93832
rect 353300 93780 353352 93832
rect 387248 93780 387300 93832
rect 399484 93780 399536 93832
rect 405188 93780 405240 93832
rect 447692 93780 447744 93832
rect 476120 93780 476172 93832
rect 387156 93712 387208 93764
rect 416780 93712 416832 93764
rect 417424 93712 417476 93764
rect 458180 93712 458232 93764
rect 391204 93644 391256 93696
rect 407120 93644 407172 93696
rect 423864 93644 423916 93696
rect 456800 93644 456852 93696
rect 393964 93576 394016 93628
rect 403256 93576 403308 93628
rect 435364 93576 435416 93628
rect 457444 93576 457496 93628
rect 382924 93508 382976 93560
rect 440608 93508 440660 93560
rect 443184 93508 443236 93560
rect 459744 93508 459796 93560
rect 130752 93372 130804 93424
rect 171784 93372 171836 93424
rect 151728 93304 151780 93356
rect 195244 93304 195296 93356
rect 113824 93236 113876 93288
rect 173348 93236 173400 93288
rect 97264 93168 97316 93220
rect 174728 93168 174780 93220
rect 121460 93100 121512 93152
rect 214932 93100 214984 93152
rect 318800 93100 318852 93152
rect 353300 93100 353352 93152
rect 416780 92828 416832 92880
rect 418068 92828 418120 92880
rect 418896 92488 418948 92540
rect 420644 92488 420696 92540
rect 422944 92488 422996 92540
rect 424508 92488 424560 92540
rect 447784 92488 447836 92540
rect 449624 92488 449676 92540
rect 98184 92420 98236 92472
rect 121460 92420 121512 92472
rect 125784 92420 125836 92472
rect 189724 92420 189776 92472
rect 192484 92420 192536 92472
rect 321560 92420 321612 92472
rect 382188 92420 382240 92472
rect 410984 92420 411036 92472
rect 120356 92352 120408 92404
rect 182916 92352 182968 92404
rect 404544 92352 404596 92404
rect 462320 92352 462372 92404
rect 116768 92284 116820 92336
rect 171876 92284 171928 92336
rect 375288 92284 375340 92336
rect 416136 92284 416188 92336
rect 432880 92284 432932 92336
rect 461032 92284 461084 92336
rect 152096 92216 152148 92268
rect 191104 92216 191156 92268
rect 386328 92216 386380 92268
rect 405740 92216 405792 92268
rect 407120 92216 407172 92268
rect 576124 92216 576176 92268
rect 133144 92148 133196 92200
rect 167920 92148 167972 92200
rect 135720 92080 135772 92132
rect 166540 92080 166592 92132
rect 405740 91740 405792 91792
rect 406476 91740 406528 91792
rect 107384 91196 107436 91248
rect 119344 91196 119396 91248
rect 98644 91128 98696 91180
rect 116584 91128 116636 91180
rect 87144 91060 87196 91112
rect 134524 91060 134576 91112
rect 416136 91060 416188 91112
rect 418988 91060 419040 91112
rect 67272 90992 67324 91044
rect 214564 90992 214616 91044
rect 369768 90992 369820 91044
rect 437388 90992 437440 91044
rect 67456 90924 67508 90976
rect 209044 90924 209096 90976
rect 340880 90924 340932 90976
rect 398196 90924 398248 90976
rect 415492 90924 415544 90976
rect 416688 90924 416740 90976
rect 462412 90924 462464 90976
rect 129464 90856 129516 90908
rect 192576 90856 192628 90908
rect 426440 90856 426492 90908
rect 427728 90856 427780 90908
rect 470692 90856 470744 90908
rect 110144 90788 110196 90840
rect 169208 90788 169260 90840
rect 124036 90720 124088 90772
rect 171968 90720 172020 90772
rect 151544 90652 151596 90704
rect 185584 90652 185636 90704
rect 216588 90380 216640 90432
rect 317512 90380 317564 90432
rect 192484 90312 192536 90364
rect 307300 90312 307352 90364
rect 311164 90312 311216 90364
rect 340880 90312 340932 90364
rect 403624 90312 403676 90364
rect 428372 90312 428424 90364
rect 66076 89632 66128 89684
rect 209136 89632 209188 89684
rect 409144 89632 409196 89684
rect 500224 89632 500276 89684
rect 117136 89564 117188 89616
rect 206468 89564 206520 89616
rect 413560 89564 413612 89616
rect 467932 89564 467984 89616
rect 99748 89496 99800 89548
rect 173440 89496 173492 89548
rect 110328 89428 110380 89480
rect 181536 89428 181588 89480
rect 151360 89360 151412 89412
rect 204904 89360 204956 89412
rect 132224 89292 132276 89344
rect 166264 89292 166316 89344
rect 310520 88952 310572 89004
rect 397460 88952 397512 89004
rect 408500 88952 408552 89004
rect 409696 88952 409748 89004
rect 427820 88952 427872 89004
rect 429016 88952 429068 89004
rect 75368 88272 75420 88324
rect 211160 88272 211212 88324
rect 401600 88272 401652 88324
rect 402612 88272 402664 88324
rect 549260 88272 549312 88324
rect 86408 88204 86460 88256
rect 164884 88204 164936 88256
rect 316040 88204 316092 88256
rect 454224 88204 454276 88256
rect 105728 88136 105780 88188
rect 184296 88136 184348 88188
rect 400864 88136 400916 88188
rect 401324 88136 401376 88188
rect 494060 88136 494112 88188
rect 134800 88068 134852 88120
rect 188344 88068 188396 88120
rect 119896 88000 119948 88052
rect 169024 88000 169076 88052
rect 121368 87932 121420 87984
rect 166356 87932 166408 87984
rect 179236 87592 179288 87644
rect 267832 87592 267884 87644
rect 355324 87592 355376 87644
rect 62028 86912 62080 86964
rect 189816 86912 189868 86964
rect 416688 86912 416740 86964
rect 418804 86912 418856 86964
rect 418988 86912 419040 86964
rect 580172 86912 580224 86964
rect 112444 86844 112496 86896
rect 211896 86844 211948 86896
rect 103336 86776 103388 86828
rect 184204 86776 184256 86828
rect 118056 86708 118108 86760
rect 193956 86708 194008 86760
rect 102968 86640 103020 86692
rect 173256 86640 173308 86692
rect 122840 86572 122892 86624
rect 167644 86572 167696 86624
rect 299388 86300 299440 86352
rect 320824 86300 320876 86352
rect 328460 86300 328512 86352
rect 374644 86300 374696 86352
rect 242900 86232 242952 86284
rect 294052 86232 294104 86284
rect 312544 86232 312596 86284
rect 401600 86232 401652 86284
rect 67548 85484 67600 85536
rect 191196 85484 191248 85536
rect 90640 85416 90692 85468
rect 211988 85416 212040 85468
rect 111064 85348 111116 85400
rect 174636 85348 174688 85400
rect 121920 85280 121972 85332
rect 183008 85280 183060 85332
rect 2780 85212 2832 85264
rect 4804 85212 4856 85264
rect 115296 85212 115348 85264
rect 167736 85212 167788 85264
rect 104716 84124 104768 84176
rect 213276 84124 213328 84176
rect 313740 84124 313792 84176
rect 466552 84124 466604 84176
rect 101956 84056 102008 84108
rect 202328 84056 202380 84108
rect 96528 83988 96580 84040
rect 170588 83988 170640 84040
rect 95148 83920 95200 83972
rect 166448 83920 166500 83972
rect 118608 83852 118660 83904
rect 189908 83852 189960 83904
rect 125416 83784 125468 83836
rect 196624 83784 196676 83836
rect 238024 83512 238076 83564
rect 251272 83512 251324 83564
rect 199384 83444 199436 83496
rect 271144 83444 271196 83496
rect 313280 82832 313332 82884
rect 313740 82832 313792 82884
rect 64788 82764 64840 82816
rect 308404 82764 308456 82816
rect 108856 82696 108908 82748
rect 207664 82696 207716 82748
rect 238760 82696 238812 82748
rect 295340 82696 295392 82748
rect 450176 82696 450228 82748
rect 125508 82628 125560 82680
rect 203616 82628 203668 82680
rect 108948 82560 109000 82612
rect 185676 82560 185728 82612
rect 97908 82492 97960 82544
rect 170496 82492 170548 82544
rect 93768 81336 93820 81388
rect 204996 81336 205048 81388
rect 126888 81268 126940 81320
rect 211804 81268 211856 81320
rect 111708 81200 111760 81252
rect 188436 81200 188488 81252
rect 100668 81132 100720 81184
rect 169116 81132 169168 81184
rect 107476 81064 107528 81116
rect 173164 81064 173216 81116
rect 185584 80656 185636 80708
rect 307208 80656 307260 80708
rect 336832 80656 336884 80708
rect 427820 80656 427872 80708
rect 92388 79976 92440 80028
rect 194048 79976 194100 80028
rect 309784 79976 309836 80028
rect 310428 79976 310480 80028
rect 419632 79976 419684 80028
rect 115848 79908 115900 79960
rect 210516 79908 210568 79960
rect 122748 79840 122800 79892
rect 213184 79840 213236 79892
rect 89628 79772 89680 79824
rect 167828 79772 167880 79824
rect 276664 79296 276716 79348
rect 310428 79296 310480 79348
rect 99288 78616 99340 78668
rect 186964 78616 187016 78668
rect 245660 78616 245712 78668
rect 411260 78616 411312 78668
rect 86868 78548 86920 78600
rect 172060 78548 172112 78600
rect 124128 78480 124180 78532
rect 206376 78480 206428 78532
rect 134524 78412 134576 78464
rect 192668 78412 192720 78464
rect 334716 77256 334768 77308
rect 336832 77256 336884 77308
rect 116584 77188 116636 77240
rect 214748 77188 214800 77240
rect 285588 77188 285640 77240
rect 286876 77188 286928 77240
rect 433340 77188 433392 77240
rect 113088 77120 113140 77172
rect 202236 77120 202288 77172
rect 75920 76576 75972 76628
rect 285128 76576 285180 76628
rect 63500 76508 63552 76560
rect 303068 76508 303120 76560
rect 85488 75828 85540 75880
rect 196716 75828 196768 75880
rect 119344 75760 119396 75812
rect 203708 75760 203760 75812
rect 139400 75216 139452 75268
rect 323584 75216 323636 75268
rect 23480 75148 23532 75200
rect 297548 75148 297600 75200
rect 67640 74468 67692 74520
rect 195336 74468 195388 74520
rect 177764 73924 177816 73976
rect 347044 73924 347096 73976
rect 35900 73856 35952 73908
rect 268476 73856 268528 73908
rect 20720 73788 20772 73840
rect 297364 73788 297416 73840
rect 346400 73788 346452 73840
rect 451556 73788 451608 73840
rect 104808 73108 104860 73160
rect 198096 73108 198148 73160
rect 438860 73108 438912 73160
rect 471980 73108 472032 73160
rect 580172 73108 580224 73160
rect 124220 72496 124272 72548
rect 250536 72496 250588 72548
rect 247684 72428 247736 72480
rect 418896 72428 418948 72480
rect 3424 71680 3476 71732
rect 44824 71680 44876 71732
rect 88340 71068 88392 71120
rect 300216 71068 300268 71120
rect 303620 71068 303672 71120
rect 396816 71068 396868 71120
rect 69020 71000 69072 71052
rect 304632 71000 304684 71052
rect 271144 69776 271196 69828
rect 451740 69776 451792 69828
rect 74540 69708 74592 69760
rect 282460 69708 282512 69760
rect 64880 69640 64932 69692
rect 305920 69640 305972 69692
rect 89720 68280 89772 68332
rect 249156 68280 249208 68332
rect 184940 66988 184992 67040
rect 315304 66988 315356 67040
rect 100760 66920 100812 66972
rect 275376 66920 275428 66972
rect 62120 66852 62172 66904
rect 304448 66852 304500 66904
rect 324964 66852 325016 66904
rect 451372 66852 451424 66904
rect 110420 65560 110472 65612
rect 263048 65560 263100 65612
rect 80060 65492 80112 65544
rect 279516 65492 279568 65544
rect 284208 64812 284260 64864
rect 447784 64812 447836 64864
rect 241520 64268 241572 64320
rect 284208 64268 284260 64320
rect 38660 64200 38712 64252
rect 285036 64200 285088 64252
rect 33140 64132 33192 64184
rect 301780 64132 301832 64184
rect 70400 62840 70452 62892
rect 269856 62840 269908 62892
rect 53840 62772 53892 62824
rect 293408 62772 293460 62824
rect 198004 61480 198056 61532
rect 273260 61480 273312 61532
rect 354036 61480 354088 61532
rect 95240 61412 95292 61464
rect 280804 61412 280856 61464
rect 71780 61344 71832 61396
rect 274088 61344 274140 61396
rect 345020 61344 345072 61396
rect 408500 61344 408552 61396
rect 460204 60664 460256 60716
rect 580172 60664 580224 60716
rect 99380 60052 99432 60104
rect 267004 60052 267056 60104
rect 269120 60052 269172 60104
rect 363604 60052 363656 60104
rect 11060 59984 11112 60036
rect 303160 59984 303212 60036
rect 355324 59984 355376 60036
rect 416780 59984 416832 60036
rect 3056 59304 3108 59356
rect 62764 59304 62816 59356
rect 350540 59304 350592 59356
rect 434720 59304 434772 59356
rect 266452 58760 266504 58812
rect 350540 58760 350592 58812
rect 106280 58692 106332 58744
rect 276756 58692 276808 58744
rect 85580 58624 85632 58676
rect 296168 58624 296220 58676
rect 341524 57944 341576 57996
rect 345020 57944 345072 57996
rect 103520 57264 103572 57316
rect 300400 57264 300452 57316
rect 13820 57196 13872 57248
rect 284944 57196 284996 57248
rect 296168 57196 296220 57248
rect 435364 57196 435416 57248
rect 255320 55972 255372 56024
rect 269764 55972 269816 56024
rect 110512 55904 110564 55956
rect 293316 55904 293368 55956
rect 19340 55836 19392 55888
rect 260196 55836 260248 55888
rect 4068 55156 4120 55208
rect 251180 55156 251232 55208
rect 262128 54544 262180 54596
rect 381544 54544 381596 54596
rect 56600 54476 56652 54528
rect 264428 54476 264480 54528
rect 3424 53796 3476 53848
rect 4068 53796 4120 53848
rect 281448 53728 281500 53780
rect 395436 53728 395488 53780
rect 73160 53116 73212 53168
rect 292120 53116 292172 53168
rect 19432 53048 19484 53100
rect 283656 53048 283708 53100
rect 280160 52436 280212 52488
rect 281448 52436 281500 52488
rect 244924 51824 244976 51876
rect 409144 51824 409196 51876
rect 45560 51756 45612 51808
rect 273996 51756 274048 51808
rect 29000 51688 29052 51740
rect 296260 51688 296312 51740
rect 51080 50396 51132 50448
rect 262956 50396 263008 50448
rect 284944 50396 284996 50448
rect 342996 50396 343048 50448
rect 67640 50328 67692 50380
rect 297456 50328 297508 50380
rect 342352 50328 342404 50380
rect 405740 50328 405792 50380
rect 77300 49036 77352 49088
rect 296076 49036 296128 49088
rect 2780 48968 2832 49020
rect 286324 48968 286376 49020
rect 298100 48968 298152 49020
rect 337476 48968 337528 49020
rect 342904 48968 342956 49020
rect 444380 48968 444432 49020
rect 291844 48288 291896 48340
rect 298100 48288 298152 48340
rect 216036 47676 216088 47728
rect 292580 47676 292632 47728
rect 373356 47676 373408 47728
rect 92480 47608 92532 47660
rect 298744 47608 298796 47660
rect 60740 47540 60792 47592
rect 294788 47540 294840 47592
rect 271696 46860 271748 46912
rect 398104 46860 398156 46912
rect 399576 46860 399628 46912
rect 580172 46860 580224 46912
rect 26240 46248 26292 46300
rect 257528 46248 257580 46300
rect 42800 46180 42852 46232
rect 292028 46180 292080 46232
rect 248420 45568 248472 45620
rect 271696 45568 271748 45620
rect 3516 45500 3568 45552
rect 48964 45500 49016 45552
rect 59360 44888 59412 44940
rect 298836 44888 298888 44940
rect 44180 44820 44232 44872
rect 287980 44820 288032 44872
rect 81440 43460 81492 43512
rect 289268 43460 289320 43512
rect 295340 43460 295392 43512
rect 329288 43460 329340 43512
rect 6920 43392 6972 43444
rect 300308 43392 300360 43444
rect 177856 42168 177908 42220
rect 337476 42168 337528 42220
rect 118700 42100 118752 42152
rect 301596 42100 301648 42152
rect 44272 42032 44324 42084
rect 262864 42032 262916 42084
rect 342260 41352 342312 41404
rect 422944 41352 422996 41404
rect 338028 41284 338080 41336
rect 359464 41284 359516 41336
rect 85672 40740 85724 40792
rect 290464 40740 290516 40792
rect 322940 40740 322992 40792
rect 342260 40740 342312 40792
rect 46940 40672 46992 40724
rect 257436 40672 257488 40724
rect 259460 40672 259512 40724
rect 336740 40672 336792 40724
rect 338028 40672 338080 40724
rect 121460 39448 121512 39500
rect 271236 39448 271288 39500
rect 256056 39380 256108 39432
rect 445852 39380 445904 39432
rect 37280 39312 37332 39364
rect 307116 39312 307168 39364
rect 209688 38564 209740 38616
rect 324320 38564 324372 38616
rect 324964 38564 325016 38616
rect 364984 38564 365036 38616
rect 365628 38564 365680 38616
rect 451280 38564 451332 38616
rect 128360 37952 128412 38004
rect 216680 37952 216732 38004
rect 251180 37952 251232 38004
rect 365076 37952 365128 38004
rect 27620 37884 27672 37936
rect 279424 37884 279476 37936
rect 329840 37884 329892 37936
rect 365628 37884 365680 37936
rect 240784 36660 240836 36712
rect 407212 36660 407264 36712
rect 11152 36592 11204 36644
rect 255964 36592 256016 36644
rect 35992 36524 36044 36576
rect 305828 36524 305880 36576
rect 179420 35300 179472 35352
rect 254676 35300 254728 35352
rect 207020 35232 207072 35284
rect 345756 35232 345808 35284
rect 48320 35164 48372 35216
rect 272524 35164 272576 35216
rect 292028 35164 292080 35216
rect 398840 35164 398892 35216
rect 427728 35164 427780 35216
rect 464620 35164 464672 35216
rect 254676 34484 254728 34536
rect 256056 34484 256108 34536
rect 143540 33872 143592 33924
rect 331956 33872 332008 33924
rect 30380 33804 30432 33856
rect 265624 33804 265676 33856
rect 52460 33736 52512 33788
rect 304356 33736 304408 33788
rect 349804 33736 349856 33788
rect 438124 33736 438176 33788
rect 3516 33056 3568 33108
rect 35164 33056 35216 33108
rect 337476 33056 337528 33108
rect 449992 33056 450044 33108
rect 464620 33056 464672 33108
rect 579896 33056 579948 33108
rect 91100 32376 91152 32428
rect 264336 32376 264388 32428
rect 309876 32376 309928 32428
rect 324964 32376 325016 32428
rect 336740 31764 336792 31816
rect 337476 31764 337528 31816
rect 320824 31696 320876 31748
rect 396908 31696 396960 31748
rect 320180 31220 320232 31272
rect 320824 31220 320876 31272
rect 201500 31152 201552 31204
rect 336004 31152 336056 31204
rect 66260 31084 66312 31136
rect 302976 31084 303028 31136
rect 5540 31016 5592 31068
rect 251916 31016 251968 31068
rect 98000 29588 98052 29640
rect 260104 29588 260156 29640
rect 317512 28908 317564 28960
rect 318708 28908 318760 28960
rect 391296 28908 391348 28960
rect 86960 28296 87012 28348
rect 287796 28296 287848 28348
rect 93860 28228 93912 28280
rect 305644 28228 305696 28280
rect 309140 27616 309192 27668
rect 318708 27616 318760 27668
rect 200120 27548 200172 27600
rect 311900 27548 311952 27600
rect 312544 27548 312596 27600
rect 117320 26936 117372 26988
rect 282276 26936 282328 26988
rect 78680 26868 78732 26920
rect 305736 26868 305788 26920
rect 336832 26188 336884 26240
rect 443000 26188 443052 26240
rect 179328 25644 179380 25696
rect 299480 25644 299532 25696
rect 300768 25644 300820 25696
rect 82820 25576 82872 25628
rect 273904 25576 273956 25628
rect 4160 25508 4212 25560
rect 298928 25508 298980 25560
rect 305644 25508 305696 25560
rect 378876 25508 378928 25560
rect 300768 24760 300820 24812
rect 369124 24760 369176 24812
rect 113180 24080 113232 24132
rect 250444 24080 250496 24132
rect 176568 23400 176620 23452
rect 331220 23400 331272 23452
rect 331220 22924 331272 22976
rect 332048 22924 332100 22976
rect 52552 22788 52604 22840
rect 293224 22788 293276 22840
rect 12440 22720 12492 22772
rect 268384 22720 268436 22772
rect 1308 22040 1360 22092
rect 249800 22040 249852 22092
rect 314660 22040 314712 22092
rect 392584 22040 392636 22092
rect 20 21564 72 21616
rect 1308 21564 1360 21616
rect 281540 21428 281592 21480
rect 314660 21428 314712 21480
rect 111800 21360 111852 21412
rect 307024 21360 307076 21412
rect 3516 20612 3568 20664
rect 22744 20612 22796 20664
rect 274640 20612 274692 20664
rect 275836 20612 275888 20664
rect 420920 20612 420972 20664
rect 498844 20612 498896 20664
rect 579896 20612 579948 20664
rect 102140 20000 102192 20052
rect 300124 20000 300176 20052
rect 57980 19932 58032 19984
rect 287888 19932 287940 19984
rect 176476 19252 176528 19304
rect 244280 19252 244332 19304
rect 244924 19252 244976 19304
rect 289728 19252 289780 19304
rect 396724 19252 396776 19304
rect 188988 18640 189040 18692
rect 260840 18640 260892 18692
rect 93952 18572 94004 18624
rect 283564 18572 283616 18624
rect 263600 17960 263652 18012
rect 289728 17960 289780 18012
rect 210424 17348 210476 17400
rect 96620 17280 96672 17332
rect 258816 17280 258868 17332
rect 259552 17280 259604 17332
rect 377404 17280 377456 17332
rect 104900 17212 104952 17264
rect 289176 17212 289228 17264
rect 179512 15988 179564 16040
rect 294880 15988 294932 16040
rect 296168 15988 296220 16040
rect 50160 15920 50212 15972
rect 257344 15920 257396 15972
rect 275928 15920 275980 15972
rect 277952 15920 278004 15972
rect 449900 15920 449952 15972
rect 69848 15852 69900 15904
rect 282368 15852 282420 15904
rect 266360 15104 266412 15156
rect 385684 15104 385736 15156
rect 108120 14492 108172 14544
rect 253296 14492 253348 14544
rect 84200 14424 84252 14476
rect 301504 14424 301556 14476
rect 271788 13744 271840 13796
rect 360936 13744 360988 13796
rect 249984 13200 250036 13252
rect 266360 13200 266412 13252
rect 177948 13132 178000 13184
rect 284944 13132 284996 13184
rect 109040 13064 109092 13116
rect 258724 13064 258776 13116
rect 348424 13064 348476 13116
rect 449072 13064 449124 13116
rect 270776 12452 270828 12504
rect 271788 12452 271840 12504
rect 285680 12384 285732 12436
rect 286968 12384 287020 12436
rect 450084 12384 450136 12436
rect 256700 11840 256752 11892
rect 285680 11840 285732 11892
rect 28448 11772 28500 11824
rect 264244 11772 264296 11824
rect 34520 11704 34572 11756
rect 294604 11704 294656 11756
rect 183560 10956 183612 11008
rect 349160 10956 349212 11008
rect 349804 10956 349856 11008
rect 345296 10888 345348 10940
rect 345756 10888 345808 10940
rect 400864 10888 400916 10940
rect 120632 10276 120684 10328
rect 253204 10276 253256 10328
rect 287980 9596 288032 9648
rect 429844 9596 429896 9648
rect 123484 9052 123536 9104
rect 275284 9052 275336 9104
rect 119896 8984 119948 9036
rect 291936 8984 291988 9036
rect 23020 8916 23072 8968
rect 295984 8916 296036 8968
rect 349436 8236 349488 8288
rect 349712 8236 349764 8288
rect 412640 8236 412692 8288
rect 309876 8168 309928 8220
rect 356796 8168 356848 8220
rect 115204 7624 115256 7676
rect 304264 7624 304316 7676
rect 4068 7556 4120 7608
rect 249064 7556 249116 7608
rect 293684 7556 293736 7608
rect 309232 7556 309284 7608
rect 309876 7556 309928 7608
rect 327080 7556 327132 7608
rect 349712 7556 349764 7608
rect 3516 6808 3568 6860
rect 31024 6808 31076 6860
rect 324964 6808 325016 6860
rect 414020 6808 414072 6860
rect 418804 6808 418856 6860
rect 580172 6808 580224 6860
rect 347044 6740 347096 6792
rect 348424 6740 348476 6792
rect 175188 6264 175240 6316
rect 302056 6264 302108 6316
rect 116400 6196 116452 6248
rect 302884 6196 302936 6248
rect 60832 6128 60884 6180
rect 287704 6128 287756 6180
rect 324412 5516 324464 5568
rect 324964 5516 325016 5568
rect 77392 4904 77444 4956
rect 261484 4836 261536 4888
rect 56048 4768 56100 4820
rect 254584 4768 254636 4820
rect 289728 4768 289780 4820
rect 395344 4768 395396 4820
rect 215944 4088 215996 4140
rect 247592 4088 247644 4140
rect 291844 4088 291896 4140
rect 298468 4088 298520 4140
rect 302056 4088 302108 4140
rect 329196 4088 329248 4140
rect 351184 4088 351236 4140
rect 351644 4088 351696 4140
rect 403624 4088 403676 4140
rect 282184 4020 282236 4072
rect 291384 4020 291436 4072
rect 292028 4020 292080 4072
rect 305644 4020 305696 4072
rect 306748 4020 306800 4072
rect 278688 3952 278740 4004
rect 288992 3952 289044 4004
rect 289728 3952 289780 4004
rect 286600 3816 286652 3868
rect 289084 3816 289136 3868
rect 132960 3612 133012 3664
rect 203524 3612 203576 3664
rect 52460 3544 52512 3596
rect 53380 3544 53432 3596
rect 85580 3544 85632 3596
rect 86500 3544 86552 3596
rect 103336 3544 103388 3596
rect 214564 3544 214616 3596
rect 242992 3544 243044 3596
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 41880 3476 41932 3528
rect 192484 3476 192536 3528
rect 235816 3476 235868 3528
rect 238024 3476 238076 3528
rect 242900 3476 242952 3528
rect 244096 3476 244148 3528
rect 276664 3476 276716 3528
rect 25320 3408 25372 3460
rect 185584 3408 185636 3460
rect 206284 3408 206336 3460
rect 268844 3408 268896 3460
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 135260 3340 135312 3392
rect 136456 3340 136508 3392
rect 277124 3272 277176 3324
rect 278044 3544 278096 3596
rect 299572 3544 299624 3596
rect 300768 3544 300820 3596
rect 309048 3544 309100 3596
rect 311164 3544 311216 3596
rect 316040 3544 316092 3596
rect 317328 3544 317380 3596
rect 322112 3544 322164 3596
rect 327080 3544 327132 3596
rect 284300 3476 284352 3528
rect 284944 3476 284996 3528
rect 298008 3476 298060 3528
rect 315028 3476 315080 3528
rect 315304 3476 315356 3528
rect 316224 3476 316276 3528
rect 331864 3612 331916 3664
rect 340972 3612 341024 3664
rect 342168 3612 342220 3664
rect 327724 3544 327776 3596
rect 336004 3544 336056 3596
rect 344560 3544 344612 3596
rect 305552 3408 305604 3460
rect 332600 3476 332652 3528
rect 333888 3476 333940 3528
rect 340972 3476 341024 3528
rect 341524 3476 341576 3528
rect 349252 3476 349304 3528
rect 350448 3476 350500 3528
rect 355324 3408 355376 3460
rect 324320 3340 324372 3392
rect 325608 3340 325660 3392
rect 271144 3000 271196 3052
rect 276020 3000 276072 3052
rect 1676 2932 1728 2984
rect 3424 2932 3476 2984
rect 40684 2048 40736 2100
rect 294696 2048 294748 2100
<< obsm1 >>
rect 68800 95100 164756 174600
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 702574 8156 703520
rect 8116 702568 8168 702574
rect 8116 702510 8168 702516
rect 24320 700330 24348 703520
rect 40512 702642 40540 703520
rect 63408 702840 63460 702846
rect 63408 702782 63460 702788
rect 53748 702704 53800 702710
rect 53748 702646 53800 702652
rect 40500 702636 40552 702642
rect 40500 702578 40552 702584
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 39304 700324 39356 700330
rect 39304 700266 39356 700272
rect 52368 700324 52420 700330
rect 52368 700266 52420 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 7564 683188 7616 683194
rect 7564 683130 7616 683136
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3148 554736 3200 554742
rect 3148 554678 3200 554684
rect 3160 553897 3188 554678
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 7576 529242 7604 683130
rect 18604 656940 18656 656946
rect 18604 656882 18656 656888
rect 17224 632120 17276 632126
rect 17224 632062 17276 632068
rect 17236 617574 17264 632062
rect 17224 617568 17276 617574
rect 17224 617510 17276 617516
rect 17224 600364 17276 600370
rect 17224 600306 17276 600312
rect 8944 587920 8996 587926
rect 8944 587862 8996 587868
rect 7564 529236 7616 529242
rect 7564 529178 7616 529184
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3424 516112 3476 516118
rect 3424 516054 3476 516060
rect 3436 514865 3464 516054
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 8208 477556 8260 477562
rect 8208 477498 8260 477504
rect 3882 475688 3938 475697
rect 3882 475623 3938 475632
rect 3896 475386 3924 475623
rect 3884 475380 3936 475386
rect 3884 475322 3936 475328
rect 4804 475380 4856 475386
rect 4804 475322 4856 475328
rect 3424 462664 3476 462670
rect 3422 462632 3424 462641
rect 3476 462632 3478 462641
rect 3422 462567 3478 462576
rect 3424 449608 3476 449614
rect 3422 449576 3424 449585
rect 3476 449576 3478 449585
rect 3422 449511 3478 449520
rect 4816 428466 4844 475322
rect 4804 428460 4856 428466
rect 4804 428402 4856 428408
rect 4066 423600 4122 423609
rect 4066 423535 4122 423544
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 4080 404530 4108 423535
rect 4804 416832 4856 416838
rect 4804 416774 4856 416780
rect 4068 404524 4120 404530
rect 4068 404466 4120 404472
rect 3976 398132 4028 398138
rect 3976 398074 4028 398080
rect 3988 397497 4016 398074
rect 3974 397488 4030 397497
rect 3974 397423 4030 397432
rect 2964 373312 3016 373318
rect 2964 373254 3016 373260
rect 2976 371385 3004 373254
rect 2962 371376 3018 371385
rect 2962 371311 3018 371320
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 2832 358456 2834 358465
rect 2778 358391 2834 358400
rect 3332 345704 3384 345710
rect 3332 345646 3384 345652
rect 3344 345409 3372 345646
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3148 320136 3200 320142
rect 3148 320078 3200 320084
rect 3160 319297 3188 320078
rect 3146 319288 3202 319297
rect 3146 319223 3202 319232
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3238 293176 3294 293185
rect 3238 293111 3294 293120
rect 3252 291854 3280 293111
rect 3240 291848 3292 291854
rect 3240 291790 3292 291796
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3988 258738 4016 397423
rect 4816 358494 4844 416774
rect 4804 358488 4856 358494
rect 4804 358430 4856 358436
rect 4068 292596 4120 292602
rect 4068 292538 4120 292544
rect 3976 258732 4028 258738
rect 3976 258674 4028 258680
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3344 238746 3372 241023
rect 3436 240106 3464 254079
rect 3424 240100 3476 240106
rect 3424 240042 3476 240048
rect 3332 238740 3384 238746
rect 3332 238682 3384 238688
rect 3424 229764 3476 229770
rect 3424 229706 3476 229712
rect 1308 214600 1360 214606
rect 1308 214542 1360 214548
rect 1320 22098 1348 214542
rect 3436 201929 3464 229706
rect 3516 216164 3568 216170
rect 3516 216106 3568 216112
rect 3528 214985 3556 216106
rect 3514 214976 3570 214985
rect 3514 214911 3570 214920
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111580 3476 111586
rect 3424 111522 3476 111528
rect 3436 110673 3464 111522
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 2780 85264 2832 85270
rect 2780 85206 2832 85212
rect 2792 84697 2820 85206
rect 2778 84688 2834 84697
rect 2778 84623 2834 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 4080 55214 4108 292538
rect 8220 267782 8248 477498
rect 8956 462670 8984 587862
rect 15108 585404 15160 585410
rect 15108 585346 15160 585352
rect 8944 462664 8996 462670
rect 8944 462606 8996 462612
rect 8944 460964 8996 460970
rect 8944 460906 8996 460912
rect 8956 449614 8984 460906
rect 8944 449608 8996 449614
rect 8944 449550 8996 449556
rect 9588 404524 9640 404530
rect 9588 404466 9640 404472
rect 9600 294642 9628 404466
rect 15120 373318 15148 585346
rect 17236 475386 17264 600306
rect 17224 475380 17276 475386
rect 17224 475322 17276 475328
rect 18616 402898 18644 656882
rect 39316 620294 39344 700266
rect 39304 620288 39356 620294
rect 39304 620230 39356 620236
rect 51080 620288 51132 620294
rect 51080 620230 51132 620236
rect 51092 619682 51120 620230
rect 51080 619676 51132 619682
rect 51080 619618 51132 619624
rect 52276 619676 52328 619682
rect 52276 619618 52328 619624
rect 40684 618316 40736 618322
rect 40684 618258 40736 618264
rect 38568 596216 38620 596222
rect 38568 596158 38620 596164
rect 38476 589552 38528 589558
rect 38476 589494 38528 589500
rect 35808 589416 35860 589422
rect 35808 589358 35860 589364
rect 31024 586628 31076 586634
rect 31024 586570 31076 586576
rect 22744 565888 22796 565894
rect 22744 565830 22796 565836
rect 21364 527128 21416 527134
rect 21364 527070 21416 527076
rect 21376 526454 21404 527070
rect 21364 526448 21416 526454
rect 21364 526390 21416 526396
rect 18604 402892 18656 402898
rect 18604 402834 18656 402840
rect 15108 373312 15160 373318
rect 15108 373254 15160 373260
rect 9588 294636 9640 294642
rect 9588 294578 9640 294584
rect 17224 291848 17276 291854
rect 17224 291790 17276 291796
rect 13084 290488 13136 290494
rect 13084 290430 13136 290436
rect 8208 267776 8260 267782
rect 8208 267718 8260 267724
rect 8944 263628 8996 263634
rect 8944 263570 8996 263576
rect 4804 253224 4856 253230
rect 4804 253166 4856 253172
rect 4816 85270 4844 253166
rect 8956 216170 8984 263570
rect 8944 216164 8996 216170
rect 8944 216106 8996 216112
rect 8944 175976 8996 175982
rect 8944 175918 8996 175924
rect 8956 111586 8984 175918
rect 13096 150414 13124 290430
rect 17236 244186 17264 291790
rect 21376 260846 21404 526390
rect 22756 404326 22784 565830
rect 27528 564460 27580 564466
rect 27528 564402 27580 564408
rect 25688 410576 25740 410582
rect 25688 410518 25740 410524
rect 25700 409902 25728 410518
rect 25688 409896 25740 409902
rect 25688 409838 25740 409844
rect 26148 409896 26200 409902
rect 26148 409838 26200 409844
rect 22744 404320 22796 404326
rect 22744 404262 22796 404268
rect 22744 303680 22796 303686
rect 22744 303622 22796 303628
rect 21364 260840 21416 260846
rect 21364 260782 21416 260788
rect 18604 257372 18656 257378
rect 18604 257314 18656 257320
rect 17224 244180 17276 244186
rect 17224 244122 17276 244128
rect 14464 213240 14516 213246
rect 14464 213182 14516 213188
rect 13084 150408 13136 150414
rect 13084 150350 13136 150356
rect 8944 111580 8996 111586
rect 8944 111522 8996 111528
rect 14476 97986 14504 213182
rect 18616 137970 18644 257314
rect 18604 137964 18656 137970
rect 18604 137906 18656 137912
rect 14464 97980 14516 97986
rect 14464 97922 14516 97928
rect 4804 85264 4856 85270
rect 4804 85206 4856 85212
rect 20720 73840 20772 73846
rect 20720 73782 20772 73788
rect 16578 72448 16634 72457
rect 16578 72383 16634 72392
rect 11060 60036 11112 60042
rect 11060 59978 11112 59984
rect 4068 55208 4120 55214
rect 4068 55150 4120 55156
rect 4080 53854 4108 55150
rect 3424 53848 3476 53854
rect 3424 53790 3476 53796
rect 4068 53848 4120 53854
rect 4068 53790 4120 53796
rect 2780 49020 2832 49026
rect 2780 48962 2832 48968
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1320 21622 1348 22034
rect 20 21616 72 21622
rect 20 21558 72 21564
rect 1308 21616 1360 21622
rect 1308 21558 1360 21564
rect 32 16574 60 21558
rect 2792 16574 2820 48962
rect 32 16546 152 16574
rect 2792 16546 2912 16574
rect 124 354 152 16546
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1688 480 1716 2926
rect 2884 480 2912 16546
rect 3436 2990 3464 53790
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 6920 43444 6972 43450
rect 6920 43386 6972 43392
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 5540 31068 5592 31074
rect 5540 31010 5592 31016
rect 4160 25560 4212 25566
rect 4160 25502 4212 25508
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3528 19417 3556 20606
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 4172 16574 4200 25502
rect 5552 16574 5580 31010
rect 6932 16574 6960 43386
rect 8298 24168 8354 24177
rect 8298 24103 8354 24112
rect 8312 16574 8340 24103
rect 4172 16546 5304 16574
rect 5552 16546 6040 16574
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3528 6497 3556 6802
rect 3514 6488 3570 6497
rect 3514 6423 3570 6432
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 4080 480 4108 7550
rect 5276 480 5304 16546
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 9678 10296 9734 10305
rect 9678 10231 9734 10240
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 10231
rect 11072 3534 11100 59978
rect 13820 57248 13872 57254
rect 13820 57190 13872 57196
rect 11152 36644 11204 36650
rect 11152 36586 11204 36592
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 36586
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12452 16574 12480 22714
rect 13832 16574 13860 57190
rect 16592 16574 16620 72383
rect 19340 55888 19392 55894
rect 19340 55830 19392 55836
rect 17958 29608 18014 29617
rect 17958 29543 18014 29552
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 16592 16546 17080 16574
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 16302 2680 16358 2689
rect 16302 2615 16358 2624
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 354 16018 480
rect 16316 354 16344 2615
rect 17052 480 17080 16546
rect 15906 326 16344 354
rect 15906 -960 16018 326
rect 17010 -960 17122 480
rect 17972 354 18000 29543
rect 19352 6914 19380 55830
rect 19432 53100 19484 53106
rect 19432 53042 19484 53048
rect 19444 16574 19472 53042
rect 20732 16574 20760 73782
rect 22756 20670 22784 303622
rect 26160 245614 26188 409838
rect 26148 245608 26200 245614
rect 26148 245550 26200 245556
rect 27540 233918 27568 564402
rect 31036 398138 31064 586570
rect 35164 585200 35216 585206
rect 35164 585142 35216 585148
rect 35176 554742 35204 585142
rect 35716 555484 35768 555490
rect 35716 555426 35768 555432
rect 35164 554736 35216 554742
rect 35164 554678 35216 554684
rect 33048 525088 33100 525094
rect 33048 525030 33100 525036
rect 31668 467900 31720 467906
rect 31668 467842 31720 467848
rect 31024 398132 31076 398138
rect 31024 398074 31076 398080
rect 31024 279472 31076 279478
rect 31024 279414 31076 279420
rect 27528 233912 27580 233918
rect 27528 233854 27580 233860
rect 23480 75200 23532 75206
rect 23480 75142 23532 75148
rect 22744 20664 22796 20670
rect 22744 20606 22796 20612
rect 23492 16574 23520 75142
rect 29000 51740 29052 51746
rect 29000 51682 29052 51688
rect 26240 46300 26292 46306
rect 26240 46242 26292 46248
rect 19444 16546 20208 16574
rect 20732 16546 21864 16574
rect 23492 16546 24256 16574
rect 19352 6886 19472 6914
rect 19444 480 19472 6886
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23032 480 23060 8910
rect 24228 480 24256 16546
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25332 480 25360 3402
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 46242
rect 27620 37936 27672 37942
rect 27620 37878 27672 37884
rect 27632 16574 27660 37878
rect 29012 16574 29040 51682
rect 30380 33856 30432 33862
rect 30380 33798 30432 33804
rect 30392 16574 30420 33798
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 27724 480 27752 16546
rect 28448 11824 28500 11830
rect 28448 11766 28500 11772
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 11766
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31036 6866 31064 279414
rect 31680 231742 31708 467842
rect 32956 423700 33008 423706
rect 32956 423642 33008 423648
rect 32968 232966 32996 423642
rect 33060 318102 33088 525030
rect 34428 451308 34480 451314
rect 34428 451250 34480 451256
rect 33048 318096 33100 318102
rect 33048 318038 33100 318044
rect 34440 313954 34468 451250
rect 34428 313948 34480 313954
rect 34428 313890 34480 313896
rect 35728 302938 35756 555426
rect 35716 302932 35768 302938
rect 35716 302874 35768 302880
rect 35716 267844 35768 267850
rect 35716 267786 35768 267792
rect 35728 234598 35756 267786
rect 35820 244254 35848 589358
rect 37188 547936 37240 547942
rect 37188 547878 37240 547884
rect 37096 464364 37148 464370
rect 37096 464306 37148 464312
rect 37108 396030 37136 464306
rect 37096 396024 37148 396030
rect 37096 395966 37148 395972
rect 37004 376780 37056 376786
rect 37004 376722 37056 376728
rect 37016 253910 37044 376722
rect 36820 253904 36872 253910
rect 36820 253846 36872 253852
rect 37004 253904 37056 253910
rect 37004 253846 37056 253852
rect 36832 253230 36860 253846
rect 36820 253224 36872 253230
rect 36820 253166 36872 253172
rect 35808 244248 35860 244254
rect 35808 244190 35860 244196
rect 37108 238814 37136 395966
rect 37096 238808 37148 238814
rect 37096 238750 37148 238756
rect 37200 235890 37228 547878
rect 38488 399498 38516 589494
rect 38476 399492 38528 399498
rect 38476 399434 38528 399440
rect 38580 252521 38608 596158
rect 39948 592068 40000 592074
rect 39948 592010 40000 592016
rect 39856 552084 39908 552090
rect 39856 552026 39908 552032
rect 39764 308508 39816 308514
rect 39764 308450 39816 308456
rect 38566 252512 38622 252521
rect 38566 252447 38622 252456
rect 37188 235884 37240 235890
rect 37188 235826 37240 235832
rect 35164 234592 35216 234598
rect 35164 234534 35216 234540
rect 35716 234592 35768 234598
rect 35716 234534 35768 234540
rect 32956 232960 33008 232966
rect 32956 232902 33008 232908
rect 31668 231736 31720 231742
rect 31668 231678 31720 231684
rect 31758 68232 31814 68241
rect 31758 68167 31814 68176
rect 31772 16574 31800 68167
rect 33140 64184 33192 64190
rect 33140 64126 33192 64132
rect 33152 16574 33180 64126
rect 35176 33114 35204 234534
rect 39776 233170 39804 308450
rect 39868 300150 39896 552026
rect 39856 300144 39908 300150
rect 39856 300086 39908 300092
rect 39960 290494 39988 592010
rect 40696 542434 40724 618258
rect 46204 605872 46256 605878
rect 46204 605814 46256 605820
rect 45468 592136 45520 592142
rect 45468 592078 45520 592084
rect 41328 590844 41380 590850
rect 41328 590786 41380 590792
rect 40684 542428 40736 542434
rect 40684 542370 40736 542376
rect 41236 538280 41288 538286
rect 41236 538222 41288 538228
rect 41144 466472 41196 466478
rect 41144 466414 41196 466420
rect 41156 397458 41184 466414
rect 41144 397452 41196 397458
rect 41144 397394 41196 397400
rect 41248 363662 41276 538222
rect 41340 398206 41368 590786
rect 42706 588024 42762 588033
rect 42706 587959 42762 587968
rect 42616 444440 42668 444446
rect 42616 444382 42668 444388
rect 41328 398200 41380 398206
rect 41328 398142 41380 398148
rect 41328 397452 41380 397458
rect 41328 397394 41380 397400
rect 41236 363656 41288 363662
rect 41236 363598 41288 363604
rect 41248 309806 41276 363598
rect 41236 309800 41288 309806
rect 41236 309742 41288 309748
rect 39948 290488 40000 290494
rect 39948 290430 40000 290436
rect 41236 284368 41288 284374
rect 41236 284310 41288 284316
rect 39948 278792 40000 278798
rect 39948 278734 40000 278740
rect 39764 233164 39816 233170
rect 39764 233106 39816 233112
rect 39960 202162 39988 278734
rect 41248 209778 41276 284310
rect 41340 273970 41368 397394
rect 42628 365022 42656 444382
rect 42616 365016 42668 365022
rect 42616 364958 42668 364964
rect 41328 273964 41380 273970
rect 41328 273906 41380 273912
rect 41328 270564 41380 270570
rect 41328 270506 41380 270512
rect 41236 209772 41288 209778
rect 41236 209714 41288 209720
rect 39948 202156 40000 202162
rect 39948 202098 40000 202104
rect 41340 187134 41368 270506
rect 42720 240786 42748 587959
rect 44822 586664 44878 586673
rect 44822 586599 44878 586608
rect 44088 586560 44140 586566
rect 44088 586502 44140 586508
rect 43994 585304 44050 585313
rect 43994 585239 44050 585248
rect 42800 542428 42852 542434
rect 42800 542370 42852 542376
rect 42812 466478 42840 542370
rect 43904 529236 43956 529242
rect 43904 529178 43956 529184
rect 43916 528630 43944 529178
rect 43904 528624 43956 528630
rect 43904 528566 43956 528572
rect 42800 466472 42852 466478
rect 42800 466414 42852 466420
rect 43812 456816 43864 456822
rect 43812 456758 43864 456764
rect 43824 311166 43852 456758
rect 43916 353258 43944 528566
rect 44008 394058 44036 585239
rect 43996 394052 44048 394058
rect 43996 393994 44048 394000
rect 43996 357468 44048 357474
rect 43996 357410 44048 357416
rect 43904 353252 43956 353258
rect 43904 353194 43956 353200
rect 43812 311160 43864 311166
rect 43812 311102 43864 311108
rect 43812 289876 43864 289882
rect 43812 289818 43864 289824
rect 42708 240780 42760 240786
rect 42708 240722 42760 240728
rect 42800 215280 42852 215286
rect 42800 215222 42852 215228
rect 42812 214606 42840 215222
rect 42800 214600 42852 214606
rect 42800 214542 42852 214548
rect 43824 209098 43852 289818
rect 43904 289128 43956 289134
rect 43904 289070 43956 289076
rect 43812 209092 43864 209098
rect 43812 209034 43864 209040
rect 43916 197305 43944 289070
rect 44008 244186 44036 357410
rect 43996 244180 44048 244186
rect 43996 244122 44048 244128
rect 44100 215286 44128 586502
rect 44836 345710 44864 586599
rect 45376 481704 45428 481710
rect 45376 481646 45428 481652
rect 45284 349852 45336 349858
rect 45284 349794 45336 349800
rect 44824 345704 44876 345710
rect 44824 345646 44876 345652
rect 44824 297424 44876 297430
rect 44824 297366 44876 297372
rect 44088 215280 44140 215286
rect 44088 215222 44140 215228
rect 43902 197296 43958 197305
rect 43902 197231 43958 197240
rect 41328 187128 41380 187134
rect 41328 187070 41380 187076
rect 35900 73908 35952 73914
rect 35900 73850 35952 73856
rect 35164 33108 35216 33114
rect 35164 33050 35216 33056
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 31024 6860 31076 6866
rect 31024 6802 31076 6808
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 34520 11756 34572 11762
rect 34520 11698 34572 11704
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 11698
rect 35912 6914 35940 73850
rect 44836 71738 44864 297366
rect 45296 267714 45324 349794
rect 45388 305658 45416 481646
rect 45480 399566 45508 592078
rect 46216 404394 46244 605814
rect 48136 590776 48188 590782
rect 48136 590718 48188 590724
rect 46848 585472 46900 585478
rect 46848 585414 46900 585420
rect 46572 441652 46624 441658
rect 46572 441594 46624 441600
rect 46204 404388 46256 404394
rect 46204 404330 46256 404336
rect 45468 399560 45520 399566
rect 45468 399502 45520 399508
rect 45468 396840 45520 396846
rect 45468 396782 45520 396788
rect 45376 305652 45428 305658
rect 45376 305594 45428 305600
rect 45284 267708 45336 267714
rect 45284 267650 45336 267656
rect 45480 237182 45508 396782
rect 46584 295322 46612 441594
rect 46756 414044 46808 414050
rect 46756 413986 46808 413992
rect 46664 394120 46716 394126
rect 46664 394062 46716 394068
rect 46572 295316 46624 295322
rect 46572 295258 46624 295264
rect 46676 238066 46704 394062
rect 46664 238060 46716 238066
rect 46664 238002 46716 238008
rect 46768 237386 46796 413986
rect 46860 303006 46888 585414
rect 48044 484424 48096 484430
rect 48044 484366 48096 484372
rect 48056 308446 48084 484366
rect 48148 402354 48176 590718
rect 50344 588328 50396 588334
rect 50344 588270 50396 588276
rect 49608 586900 49660 586906
rect 49608 586842 49660 586848
rect 49516 586832 49568 586838
rect 49516 586774 49568 586780
rect 48228 585268 48280 585274
rect 48228 585210 48280 585216
rect 48136 402348 48188 402354
rect 48136 402290 48188 402296
rect 48136 396772 48188 396778
rect 48136 396714 48188 396720
rect 48044 308440 48096 308446
rect 48044 308382 48096 308388
rect 46848 303000 46900 303006
rect 46848 302942 46900 302948
rect 48044 287088 48096 287094
rect 48044 287030 48096 287036
rect 46848 276072 46900 276078
rect 46848 276014 46900 276020
rect 46756 237380 46808 237386
rect 46756 237322 46808 237328
rect 45468 237176 45520 237182
rect 45468 237118 45520 237124
rect 46860 189990 46888 276014
rect 48056 211886 48084 287030
rect 48148 235822 48176 396714
rect 48240 240106 48268 585210
rect 48964 527196 49016 527202
rect 48964 527138 49016 527144
rect 48976 404258 49004 527138
rect 49424 463752 49476 463758
rect 49424 463694 49476 463700
rect 48964 404252 49016 404258
rect 48964 404194 49016 404200
rect 49436 355434 49464 463694
rect 49424 355428 49476 355434
rect 49424 355370 49476 355376
rect 49424 347064 49476 347070
rect 49424 347006 49476 347012
rect 48964 267776 49016 267782
rect 48964 267718 49016 267724
rect 48228 240100 48280 240106
rect 48228 240042 48280 240048
rect 48240 239426 48268 240042
rect 48228 239420 48280 239426
rect 48228 239362 48280 239368
rect 48976 238882 49004 267718
rect 49436 266354 49464 347006
rect 49528 337414 49556 586774
rect 49516 337408 49568 337414
rect 49516 337350 49568 337356
rect 49620 315314 49648 586842
rect 50356 410582 50384 588270
rect 50988 585540 51040 585546
rect 50988 585482 51040 585488
rect 50436 501016 50488 501022
rect 50436 500958 50488 500964
rect 50344 410576 50396 410582
rect 50344 410518 50396 410524
rect 50448 404462 50476 500958
rect 50712 420980 50764 420986
rect 50712 420922 50764 420928
rect 50436 404456 50488 404462
rect 50436 404398 50488 404404
rect 49608 315308 49660 315314
rect 49608 315250 49660 315256
rect 50724 296750 50752 420922
rect 50896 400920 50948 400926
rect 50896 400862 50948 400868
rect 50804 378888 50856 378894
rect 50804 378830 50856 378836
rect 50712 296744 50764 296750
rect 50712 296686 50764 296692
rect 49608 290488 49660 290494
rect 49608 290430 49660 290436
rect 49620 289950 49648 290430
rect 49608 289944 49660 289950
rect 49608 289886 49660 289892
rect 49424 266348 49476 266354
rect 49424 266290 49476 266296
rect 49516 263696 49568 263702
rect 49516 263638 49568 263644
rect 48964 238876 49016 238882
rect 48964 238818 49016 238824
rect 48136 235816 48188 235822
rect 48136 235758 48188 235764
rect 48044 211880 48096 211886
rect 48044 211822 48096 211828
rect 49528 208350 49556 263638
rect 49620 224942 49648 289886
rect 50724 284306 50752 296686
rect 50712 284300 50764 284306
rect 50712 284242 50764 284248
rect 50816 247042 50844 378830
rect 50804 247036 50856 247042
rect 50804 246978 50856 246984
rect 50908 238542 50936 400862
rect 51000 367810 51028 585482
rect 52184 450560 52236 450566
rect 52184 450502 52236 450508
rect 51080 428460 51132 428466
rect 51080 428402 51132 428408
rect 51092 427854 51120 428402
rect 51080 427848 51132 427854
rect 51080 427790 51132 427796
rect 52092 427848 52144 427854
rect 52092 427790 52144 427796
rect 52104 388550 52132 427790
rect 52092 388544 52144 388550
rect 52092 388486 52144 388492
rect 52196 369238 52224 450502
rect 52288 402490 52316 619618
rect 52276 402484 52328 402490
rect 52276 402426 52328 402432
rect 52380 385014 52408 700266
rect 53564 594856 53616 594862
rect 53564 594798 53616 594804
rect 53472 430636 53524 430642
rect 53472 430578 53524 430584
rect 52368 385008 52420 385014
rect 52368 384950 52420 384956
rect 52380 373994 52408 384950
rect 52288 373966 52408 373994
rect 52184 369232 52236 369238
rect 52184 369174 52236 369180
rect 50988 367804 51040 367810
rect 50988 367746 51040 367752
rect 50988 285728 51040 285734
rect 50988 285670 51040 285676
rect 50896 238536 50948 238542
rect 50896 238478 50948 238484
rect 49608 224936 49660 224942
rect 49608 224878 49660 224884
rect 49516 208344 49568 208350
rect 49516 208286 49568 208292
rect 46848 189984 46900 189990
rect 46848 189926 46900 189932
rect 51000 186969 51028 285670
rect 52184 280220 52236 280226
rect 52184 280162 52236 280168
rect 52196 195294 52224 280162
rect 52288 249762 52316 373966
rect 52368 370524 52420 370530
rect 52368 370466 52420 370472
rect 52276 249756 52328 249762
rect 52276 249698 52328 249704
rect 52380 233102 52408 370466
rect 53484 366382 53512 430578
rect 53576 400994 53604 594798
rect 53656 568608 53708 568614
rect 53656 568550 53708 568556
rect 53564 400988 53616 400994
rect 53564 400930 53616 400936
rect 53472 366376 53524 366382
rect 53472 366318 53524 366324
rect 53564 298784 53616 298790
rect 53564 298726 53616 298732
rect 52460 298104 52512 298110
rect 52460 298046 52512 298052
rect 52472 297430 52500 298046
rect 52460 297424 52512 297430
rect 52460 297366 52512 297372
rect 53472 267776 53524 267782
rect 53472 267718 53524 267724
rect 52368 233096 52420 233102
rect 52368 233038 52420 233044
rect 53484 217297 53512 267718
rect 53576 241466 53604 298726
rect 53668 298110 53696 568550
rect 53760 407794 53788 702646
rect 63132 607232 63184 607238
rect 63132 607174 63184 607180
rect 54944 593428 54996 593434
rect 54944 593370 54996 593376
rect 54484 532024 54536 532030
rect 54484 531966 54536 531972
rect 53840 525768 53892 525774
rect 53840 525710 53892 525716
rect 53852 525094 53880 525710
rect 53840 525088 53892 525094
rect 53840 525030 53892 525036
rect 53748 407788 53800 407794
rect 53748 407730 53800 407736
rect 53760 369170 53788 407730
rect 53748 369164 53800 369170
rect 53748 369106 53800 369112
rect 53748 354000 53800 354006
rect 53748 353942 53800 353948
rect 53656 298104 53708 298110
rect 53656 298046 53708 298052
rect 53656 277432 53708 277438
rect 53656 277374 53708 277380
rect 53564 241460 53616 241466
rect 53564 241402 53616 241408
rect 53470 217288 53526 217297
rect 53470 217223 53526 217232
rect 53668 203658 53696 277374
rect 53760 258058 53788 353942
rect 54496 270570 54524 531966
rect 54956 396914 54984 593370
rect 55036 591320 55088 591326
rect 55036 591262 55088 591268
rect 55048 525774 55076 591262
rect 60004 590912 60056 590918
rect 60004 590854 60056 590860
rect 56324 590708 56376 590714
rect 56324 590650 56376 590656
rect 56232 588124 56284 588130
rect 56232 588066 56284 588072
rect 55128 571396 55180 571402
rect 55128 571338 55180 571344
rect 55036 525768 55088 525774
rect 55036 525710 55088 525716
rect 55036 524340 55088 524346
rect 55036 524282 55088 524288
rect 54944 396908 54996 396914
rect 54944 396850 54996 396856
rect 54944 352572 54996 352578
rect 54944 352514 54996 352520
rect 54852 276004 54904 276010
rect 54852 275946 54904 275952
rect 54864 275913 54892 275946
rect 54850 275904 54906 275913
rect 54850 275839 54906 275848
rect 54484 270564 54536 270570
rect 54484 270506 54536 270512
rect 54852 263628 54904 263634
rect 54852 263570 54904 263576
rect 53748 258052 53800 258058
rect 53748 257994 53800 258000
rect 53760 257378 53788 257994
rect 53748 257372 53800 257378
rect 53748 257314 53800 257320
rect 54758 238368 54814 238377
rect 54758 238303 54814 238312
rect 54772 237318 54800 238303
rect 54760 237312 54812 237318
rect 54760 237254 54812 237260
rect 54864 224874 54892 263570
rect 54956 237250 54984 352514
rect 55048 238746 55076 524282
rect 55140 276010 55168 571338
rect 56244 403714 56272 588066
rect 56232 403708 56284 403714
rect 56232 403650 56284 403656
rect 56336 403646 56364 590650
rect 59084 589348 59136 589354
rect 59084 589290 59136 589296
rect 57704 588260 57756 588266
rect 57704 588202 57756 588208
rect 57244 586696 57296 586702
rect 57244 586638 57296 586644
rect 56506 583944 56562 583953
rect 56506 583879 56562 583888
rect 56520 545834 56548 583879
rect 56508 545828 56560 545834
rect 56508 545770 56560 545776
rect 56416 488572 56468 488578
rect 56416 488514 56468 488520
rect 56324 403640 56376 403646
rect 56324 403582 56376 403588
rect 56428 287054 56456 488514
rect 56336 287026 56456 287054
rect 56336 280838 56364 287026
rect 56324 280832 56376 280838
rect 56324 280774 56376 280780
rect 55128 276004 55180 276010
rect 55128 275946 55180 275952
rect 56232 273284 56284 273290
rect 56232 273226 56284 273232
rect 55128 262268 55180 262274
rect 55128 262210 55180 262216
rect 55036 238740 55088 238746
rect 55036 238682 55088 238688
rect 54944 237244 54996 237250
rect 54944 237186 54996 237192
rect 54852 224868 54904 224874
rect 54852 224810 54904 224816
rect 53656 203652 53708 203658
rect 53656 203594 53708 203600
rect 52184 195288 52236 195294
rect 52184 195230 52236 195236
rect 55140 194002 55168 262210
rect 56244 227662 56272 273226
rect 56336 228546 56364 280774
rect 56520 277394 56548 545770
rect 57256 524346 57284 586638
rect 57612 579692 57664 579698
rect 57612 579634 57664 579640
rect 57244 524340 57296 524346
rect 57244 524282 57296 524288
rect 57624 402286 57652 579634
rect 57716 405074 57744 588202
rect 58990 584080 59046 584089
rect 58990 584015 59046 584024
rect 59004 532030 59032 584015
rect 59096 556170 59124 589290
rect 59268 588192 59320 588198
rect 59268 588134 59320 588140
rect 59176 575544 59228 575550
rect 59176 575486 59228 575492
rect 59084 556164 59136 556170
rect 59084 556106 59136 556112
rect 59096 555490 59124 556106
rect 59084 555484 59136 555490
rect 59084 555426 59136 555432
rect 59084 535492 59136 535498
rect 59084 535434 59136 535440
rect 58992 532024 59044 532030
rect 58992 531966 59044 531972
rect 57796 504552 57848 504558
rect 57796 504494 57848 504500
rect 57704 405068 57756 405074
rect 57704 405010 57756 405016
rect 57612 402280 57664 402286
rect 57612 402222 57664 402228
rect 57808 313274 57836 504494
rect 57888 491360 57940 491366
rect 57888 491302 57940 491308
rect 57796 313268 57848 313274
rect 57796 313210 57848 313216
rect 57244 292664 57296 292670
rect 57244 292606 57296 292612
rect 56428 277366 56548 277394
rect 56428 276690 56456 277366
rect 56416 276684 56468 276690
rect 56416 276626 56468 276632
rect 56428 267734 56456 276626
rect 56508 273964 56560 273970
rect 56508 273906 56560 273912
rect 56520 273290 56548 273906
rect 56508 273284 56560 273290
rect 56508 273226 56560 273232
rect 56428 267706 56548 267734
rect 56416 251864 56468 251870
rect 56416 251806 56468 251812
rect 56324 228540 56376 228546
rect 56324 228482 56376 228488
rect 56232 227656 56284 227662
rect 56232 227598 56284 227604
rect 56428 195265 56456 251806
rect 56414 195256 56470 195265
rect 56414 195191 56470 195200
rect 55128 193996 55180 194002
rect 55128 193938 55180 193944
rect 56520 192545 56548 267706
rect 56506 192536 56562 192545
rect 56506 192471 56562 192480
rect 50986 186960 51042 186969
rect 50986 186895 51042 186904
rect 48964 184272 49016 184278
rect 48964 184214 49016 184220
rect 44824 71732 44876 71738
rect 44824 71674 44876 71680
rect 38660 64252 38712 64258
rect 38660 64194 38712 64200
rect 37280 39364 37332 39370
rect 37280 39306 37332 39312
rect 35992 36576 36044 36582
rect 35992 36518 36044 36524
rect 36004 16574 36032 36518
rect 37292 16574 37320 39306
rect 38672 16574 38700 64194
rect 45560 51808 45612 51814
rect 45560 51750 45612 51756
rect 42800 46232 42852 46238
rect 42800 46174 42852 46180
rect 36004 16546 36768 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 35912 6886 36032 6914
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 40684 2100 40736 2106
rect 40684 2042 40736 2048
rect 40696 480 40724 2042
rect 41892 480 41920 3470
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42812 354 42840 46174
rect 44180 44872 44232 44878
rect 44180 44814 44232 44820
rect 44192 6914 44220 44814
rect 44272 42084 44324 42090
rect 44272 42026 44324 42032
rect 44284 16574 44312 42026
rect 45572 16574 45600 51750
rect 48976 45558 49004 184214
rect 57256 164218 57284 292606
rect 57796 258120 57848 258126
rect 57796 258062 57848 258068
rect 57702 251152 57758 251161
rect 57702 251087 57758 251096
rect 57716 249898 57744 251087
rect 57704 249892 57756 249898
rect 57704 249834 57756 249840
rect 57716 222086 57744 249834
rect 57704 222080 57756 222086
rect 57704 222022 57756 222028
rect 57808 200870 57836 258062
rect 57900 238610 57928 491302
rect 58992 471708 59044 471714
rect 58992 471650 59044 471656
rect 59004 464370 59032 471650
rect 58992 464364 59044 464370
rect 58992 464306 59044 464312
rect 58992 411324 59044 411330
rect 58992 411266 59044 411272
rect 58622 392048 58678 392057
rect 58622 391983 58678 391992
rect 58636 278798 58664 391983
rect 59004 329118 59032 411266
rect 59096 393281 59124 535434
rect 59082 393272 59138 393281
rect 59082 393207 59138 393216
rect 59096 392057 59124 393207
rect 59082 392048 59138 392057
rect 59082 391983 59138 391992
rect 58992 329112 59044 329118
rect 58992 329054 59044 329060
rect 59188 316742 59216 575486
rect 59280 320142 59308 588134
rect 60016 450566 60044 590854
rect 60556 587988 60608 587994
rect 60556 587930 60608 587936
rect 60462 511864 60518 511873
rect 60462 511799 60518 511808
rect 60004 450560 60056 450566
rect 60004 450502 60056 450508
rect 60372 448588 60424 448594
rect 60372 448530 60424 448536
rect 60384 387802 60412 448530
rect 60372 387796 60424 387802
rect 60372 387738 60424 387744
rect 60476 374678 60504 511799
rect 60568 402422 60596 587930
rect 60740 585336 60792 585342
rect 60740 585278 60792 585284
rect 60752 579698 60780 585278
rect 61382 585168 61438 585177
rect 61382 585103 61438 585112
rect 60740 579692 60792 579698
rect 60740 579634 60792 579640
rect 60646 579184 60702 579193
rect 60646 579119 60702 579128
rect 60556 402416 60608 402422
rect 60556 402358 60608 402364
rect 60556 387796 60608 387802
rect 60556 387738 60608 387744
rect 60568 387122 60596 387738
rect 60556 387116 60608 387122
rect 60556 387058 60608 387064
rect 60464 374672 60516 374678
rect 60464 374614 60516 374620
rect 59268 320136 59320 320142
rect 59268 320078 59320 320084
rect 59280 319462 59308 320078
rect 59268 319456 59320 319462
rect 59268 319398 59320 319404
rect 59176 316736 59228 316742
rect 59176 316678 59228 316684
rect 59268 315308 59320 315314
rect 59268 315250 59320 315256
rect 59280 314702 59308 315250
rect 59268 314696 59320 314702
rect 59268 314638 59320 314644
rect 59084 300892 59136 300898
rect 59084 300834 59136 300840
rect 58716 292800 58768 292806
rect 58716 292742 58768 292748
rect 58624 278792 58676 278798
rect 58624 278734 58676 278740
rect 57888 238604 57940 238610
rect 57888 238546 57940 238552
rect 57796 200864 57848 200870
rect 57796 200806 57848 200812
rect 58728 189038 58756 292742
rect 59096 267646 59124 300834
rect 59176 270564 59228 270570
rect 59176 270506 59228 270512
rect 59084 267640 59136 267646
rect 59084 267582 59136 267588
rect 59084 247104 59136 247110
rect 59084 247046 59136 247052
rect 59096 225622 59124 247046
rect 59188 230450 59216 270506
rect 59280 238950 59308 314638
rect 60464 296064 60516 296070
rect 60464 296006 60516 296012
rect 60372 262336 60424 262342
rect 60372 262278 60424 262284
rect 59268 238944 59320 238950
rect 59268 238886 59320 238892
rect 59176 230444 59228 230450
rect 59176 230386 59228 230392
rect 59084 225616 59136 225622
rect 59084 225558 59136 225564
rect 60384 215218 60412 262278
rect 60476 239018 60504 296006
rect 60568 262206 60596 387058
rect 60556 262200 60608 262206
rect 60556 262142 60608 262148
rect 60556 255332 60608 255338
rect 60556 255274 60608 255280
rect 60464 239012 60516 239018
rect 60464 238954 60516 238960
rect 60372 215212 60424 215218
rect 60372 215154 60424 215160
rect 58716 189032 58768 189038
rect 58716 188974 58768 188980
rect 60568 182918 60596 255274
rect 60660 238513 60688 579119
rect 60738 572384 60794 572393
rect 60738 572319 60794 572328
rect 60752 571402 60780 572319
rect 60740 571396 60792 571402
rect 60740 571338 60792 571344
rect 60738 568984 60794 568993
rect 60738 568919 60794 568928
rect 60752 568614 60780 568919
rect 60740 568608 60792 568614
rect 60740 568550 60792 568556
rect 60738 565584 60794 565593
rect 60738 565519 60794 565528
rect 60752 564466 60780 565519
rect 60740 564460 60792 564466
rect 60740 564402 60792 564408
rect 60740 556164 60792 556170
rect 60740 556106 60792 556112
rect 60752 555393 60780 556106
rect 60738 555384 60794 555393
rect 60738 555319 60794 555328
rect 60738 552664 60794 552673
rect 60738 552599 60794 552608
rect 60752 552090 60780 552599
rect 60740 552084 60792 552090
rect 60740 552026 60792 552032
rect 60738 549264 60794 549273
rect 60738 549199 60794 549208
rect 60752 547942 60780 549199
rect 60740 547936 60792 547942
rect 60740 547878 60792 547884
rect 60738 545864 60794 545873
rect 60738 545799 60740 545808
rect 60792 545799 60794 545808
rect 60740 545770 60792 545776
rect 60738 542464 60794 542473
rect 60738 542399 60740 542408
rect 60792 542399 60794 542408
rect 60740 542370 60792 542376
rect 60738 539064 60794 539073
rect 60738 538999 60794 539008
rect 60752 538286 60780 538999
rect 60740 538280 60792 538286
rect 60740 538222 60792 538228
rect 60738 532264 60794 532273
rect 60738 532199 60794 532208
rect 60752 532030 60780 532199
rect 60740 532024 60792 532030
rect 60740 531966 60792 531972
rect 60738 528864 60794 528873
rect 60738 528799 60794 528808
rect 60752 528630 60780 528799
rect 60740 528624 60792 528630
rect 60740 528566 60792 528572
rect 60740 525768 60792 525774
rect 60740 525710 60792 525716
rect 60752 525473 60780 525710
rect 60738 525464 60794 525473
rect 60738 525399 60794 525408
rect 60738 492144 60794 492153
rect 60738 492079 60794 492088
rect 60752 491366 60780 492079
rect 60740 491360 60792 491366
rect 60740 491302 60792 491308
rect 60738 488744 60794 488753
rect 60738 488679 60794 488688
rect 60752 488578 60780 488679
rect 60740 488572 60792 488578
rect 60740 488514 60792 488520
rect 60738 485344 60794 485353
rect 60738 485279 60794 485288
rect 60752 484430 60780 485279
rect 60740 484424 60792 484430
rect 60740 484366 60792 484372
rect 60738 481944 60794 481953
rect 60738 481879 60794 481888
rect 60752 481710 60780 481879
rect 60740 481704 60792 481710
rect 60740 481646 60792 481652
rect 60738 478544 60794 478553
rect 60738 478479 60794 478488
rect 60752 477562 60780 478479
rect 60740 477556 60792 477562
rect 60740 477498 60792 477504
rect 60738 468344 60794 468353
rect 60738 468279 60794 468288
rect 60752 467906 60780 468279
rect 60740 467900 60792 467906
rect 60740 467842 60792 467848
rect 60738 464944 60794 464953
rect 60738 464879 60794 464888
rect 60752 463758 60780 464879
rect 60740 463752 60792 463758
rect 60740 463694 60792 463700
rect 60738 458144 60794 458153
rect 60738 458079 60794 458088
rect 60752 456822 60780 458079
rect 60740 456816 60792 456822
rect 60740 456758 60792 456764
rect 60738 452024 60794 452033
rect 60738 451959 60794 451968
rect 60752 451314 60780 451959
rect 60740 451308 60792 451314
rect 60740 451250 60792 451256
rect 60738 445224 60794 445233
rect 60738 445159 60794 445168
rect 60752 444446 60780 445159
rect 60740 444440 60792 444446
rect 60740 444382 60792 444388
rect 60738 441824 60794 441833
rect 60738 441759 60794 441768
rect 60752 441658 60780 441759
rect 60740 441652 60792 441658
rect 60740 441594 60792 441600
rect 60738 431624 60794 431633
rect 60738 431559 60794 431568
rect 60752 430642 60780 431559
rect 60740 430636 60792 430642
rect 60740 430578 60792 430584
rect 60738 428224 60794 428233
rect 60738 428159 60794 428168
rect 60752 427854 60780 428159
rect 60740 427848 60792 427854
rect 60740 427790 60792 427796
rect 60738 424824 60794 424833
rect 60738 424759 60794 424768
rect 60752 423706 60780 424759
rect 60740 423700 60792 423706
rect 60740 423642 60792 423648
rect 60738 421424 60794 421433
rect 60738 421359 60794 421368
rect 60752 420986 60780 421359
rect 60740 420980 60792 420986
rect 60740 420922 60792 420928
rect 61014 418024 61070 418033
rect 61014 417959 61070 417968
rect 61028 416838 61056 417959
rect 61016 416832 61068 416838
rect 61016 416774 61068 416780
rect 60830 414624 60886 414633
rect 60830 414559 60886 414568
rect 60844 414050 60872 414559
rect 60832 414044 60884 414050
rect 60832 413986 60884 413992
rect 61396 411330 61424 585103
rect 61476 584588 61528 584594
rect 61476 584530 61528 584536
rect 61488 516118 61516 584530
rect 61566 575784 61622 575793
rect 61566 575719 61622 575728
rect 61580 575550 61608 575719
rect 61568 575544 61620 575550
rect 61568 575486 61620 575492
rect 61566 535664 61622 535673
rect 61566 535599 61622 535608
rect 61580 535498 61608 535599
rect 61568 535492 61620 535498
rect 61568 535434 61620 535440
rect 61476 516112 61528 516118
rect 61476 516054 61528 516060
rect 61474 508464 61530 508473
rect 61474 508399 61530 508408
rect 61488 448594 61516 508399
rect 63144 505073 63172 607174
rect 63316 603152 63368 603158
rect 63316 603094 63368 603100
rect 63224 586764 63276 586770
rect 63224 586706 63276 586712
rect 62302 505064 62358 505073
rect 62302 504999 62358 505008
rect 63130 505064 63186 505073
rect 63130 504999 63186 505008
rect 62316 504558 62344 504999
rect 62304 504552 62356 504558
rect 62304 504494 62356 504500
rect 62026 502344 62082 502353
rect 62026 502279 62082 502288
rect 61934 498944 61990 498953
rect 61934 498879 61990 498888
rect 61842 448624 61898 448633
rect 61476 448588 61528 448594
rect 61842 448559 61898 448568
rect 61476 448530 61528 448536
rect 61384 411324 61436 411330
rect 61384 411266 61436 411272
rect 60738 407824 60794 407833
rect 60738 407759 60740 407768
rect 60792 407759 60794 407768
rect 60740 407730 60792 407736
rect 61856 394670 61884 448559
rect 61948 405006 61976 498879
rect 61936 405000 61988 405006
rect 61936 404942 61988 404948
rect 61844 394664 61896 394670
rect 61844 394606 61896 394612
rect 61844 269136 61896 269142
rect 61844 269078 61896 269084
rect 61660 254040 61712 254046
rect 61660 253982 61712 253988
rect 60646 238504 60702 238513
rect 60646 238439 60702 238448
rect 61672 229090 61700 253982
rect 61752 241528 61804 241534
rect 61752 241470 61804 241476
rect 61764 231810 61792 241470
rect 61752 231804 61804 231810
rect 61752 231746 61804 231752
rect 61660 229084 61712 229090
rect 61660 229026 61712 229032
rect 61856 207670 61884 269078
rect 61948 262138 61976 404942
rect 62040 398834 62068 502279
rect 62762 495544 62818 495553
rect 62762 495479 62818 495488
rect 62040 398806 62160 398834
rect 62132 398138 62160 398806
rect 62120 398132 62172 398138
rect 62120 398074 62172 398080
rect 62028 394664 62080 394670
rect 62028 394606 62080 394612
rect 62040 393990 62068 394606
rect 62028 393984 62080 393990
rect 62028 393926 62080 393932
rect 61936 262132 61988 262138
rect 61936 262074 61988 262080
rect 61936 253972 61988 253978
rect 61936 253914 61988 253920
rect 61948 235618 61976 253914
rect 62040 252550 62068 393926
rect 62776 383654 62804 495479
rect 63130 461544 63186 461553
rect 63130 461479 63186 461488
rect 63144 460970 63172 461479
rect 63132 460964 63184 460970
rect 63132 460906 63184 460912
rect 63144 401062 63172 460906
rect 63236 436801 63264 586706
rect 63222 436792 63278 436801
rect 63222 436727 63278 436736
rect 63328 414633 63356 603094
rect 63420 471753 63448 702782
rect 72988 702778 73016 703520
rect 72976 702772 73028 702778
rect 72976 702714 73028 702720
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 618934 88380 702406
rect 105464 699718 105492 703520
rect 130384 702500 130436 702506
rect 130384 702442 130436 702448
rect 102784 699712 102836 699718
rect 102784 699654 102836 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 88340 618928 88392 618934
rect 88340 618870 88392 618876
rect 63500 605872 63552 605878
rect 63500 605814 63552 605820
rect 63512 579193 63540 605814
rect 86224 604512 86276 604518
rect 86224 604454 86276 604460
rect 80704 599004 80756 599010
rect 80704 598946 80756 598952
rect 77484 589416 77536 589422
rect 77484 589358 77536 589364
rect 67916 585540 67968 585546
rect 67916 585482 67968 585488
rect 67928 584868 67956 585482
rect 71136 585404 71188 585410
rect 71136 585346 71188 585352
rect 71148 584868 71176 585346
rect 74354 585304 74410 585313
rect 74354 585239 74410 585248
rect 74368 584868 74396 585239
rect 77496 584882 77524 589358
rect 80716 586673 80744 598946
rect 86236 590918 86264 604454
rect 102796 596834 102824 699654
rect 119344 605940 119396 605946
rect 119344 605882 119396 605888
rect 112444 601724 112496 601730
rect 112444 601666 112496 601672
rect 90364 596828 90416 596834
rect 90364 596770 90416 596776
rect 102784 596828 102836 596834
rect 102784 596770 102836 596776
rect 86224 590912 86276 590918
rect 86224 590854 86276 590860
rect 86500 590912 86552 590918
rect 86500 590854 86552 590860
rect 83372 586900 83424 586906
rect 83372 586842 83424 586848
rect 80702 586664 80758 586673
rect 80702 586599 80758 586608
rect 80716 586514 80744 586599
rect 80624 586486 80744 586514
rect 80624 584882 80652 586486
rect 77496 584854 77602 584882
rect 80178 584854 80652 584882
rect 83384 584868 83412 586842
rect 86512 584882 86540 590854
rect 90376 588266 90404 596770
rect 92940 595468 92992 595474
rect 92940 595410 92992 595416
rect 92952 590850 92980 595410
rect 92940 590844 92992 590850
rect 92940 590786 92992 590792
rect 90364 588260 90416 588266
rect 90364 588202 90416 588208
rect 90376 586514 90404 588202
rect 90192 586486 90404 586514
rect 90192 584882 90220 586486
rect 86512 584854 86618 584882
rect 89838 584854 90220 584882
rect 92952 584882 92980 590786
rect 106188 589960 106240 589966
rect 106188 589902 106240 589908
rect 106200 589558 106228 589902
rect 105820 589552 105872 589558
rect 105820 589494 105872 589500
rect 106188 589552 106240 589558
rect 106188 589494 106240 589500
rect 99380 589484 99432 589490
rect 99380 589426 99432 589432
rect 96252 586832 96304 586838
rect 96252 586774 96304 586780
rect 92952 584854 93058 584882
rect 96264 584868 96292 586774
rect 99392 584882 99420 589426
rect 102692 585472 102744 585478
rect 102692 585414 102744 585420
rect 99392 584854 99498 584882
rect 102704 584868 102732 585414
rect 105832 584882 105860 589494
rect 112456 588198 112484 601666
rect 119356 593473 119384 605882
rect 127624 594108 127676 594114
rect 127624 594050 127676 594056
rect 118698 593464 118754 593473
rect 118698 593399 118754 593408
rect 119342 593464 119398 593473
rect 119342 593399 119398 593408
rect 112444 588192 112496 588198
rect 112444 588134 112496 588140
rect 109132 585268 109184 585274
rect 109132 585210 109184 585216
rect 105832 584854 105938 584882
rect 109144 584868 109172 585210
rect 112456 584882 112484 588134
rect 115570 586800 115626 586809
rect 115570 586735 115626 586744
rect 112378 584854 112484 584882
rect 115584 584868 115612 586735
rect 118712 584882 118740 593399
rect 127636 592142 127664 594050
rect 127624 592136 127676 592142
rect 127624 592078 127676 592084
rect 122012 586832 122064 586838
rect 122012 586774 122064 586780
rect 118712 584854 118818 584882
rect 122024 584868 122052 586774
rect 125232 586560 125284 586566
rect 125232 586502 125284 586508
rect 127636 586514 127664 592078
rect 130396 588130 130424 702442
rect 137848 700330 137876 703520
rect 154132 700330 154160 703520
rect 170324 702434 170352 703520
rect 202800 702710 202828 703520
rect 218992 702846 219020 703520
rect 218980 702840 219032 702846
rect 218980 702782 219032 702788
rect 202788 702704 202840 702710
rect 202788 702646 202840 702652
rect 217324 702636 217376 702642
rect 217324 702578 217376 702584
rect 210424 702568 210476 702574
rect 210424 702510 210476 702516
rect 169772 702406 170352 702434
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 154120 700324 154172 700330
rect 154120 700266 154172 700272
rect 169772 614786 169800 702406
rect 185584 619676 185636 619682
rect 185584 619618 185636 619624
rect 169760 614780 169812 614786
rect 169760 614722 169812 614728
rect 178684 611380 178736 611386
rect 178684 611322 178736 611328
rect 169024 607368 169076 607374
rect 169024 607310 169076 607316
rect 166264 604580 166316 604586
rect 166264 604522 166316 604528
rect 134524 600432 134576 600438
rect 134524 600374 134576 600380
rect 130384 588124 130436 588130
rect 130384 588066 130436 588072
rect 130396 586514 130424 588066
rect 125244 584868 125272 586502
rect 127636 586486 127756 586514
rect 130396 586486 130608 586514
rect 127728 584882 127756 586486
rect 130580 584882 130608 586486
rect 134246 585168 134302 585177
rect 134246 585103 134302 585112
rect 134260 584882 134288 585103
rect 134536 584882 134564 600374
rect 140228 597916 140280 597922
rect 140228 597858 140280 597864
rect 140240 596174 140268 597858
rect 153844 596352 153896 596358
rect 153844 596294 153896 596300
rect 143540 596216 143592 596222
rect 140240 596146 140636 596174
rect 143592 596164 143856 596174
rect 143540 596158 143856 596164
rect 143552 596146 143856 596158
rect 140608 594862 140636 596146
rect 140596 594856 140648 594862
rect 140596 594798 140648 594804
rect 137468 586764 137520 586770
rect 137468 586706 137520 586712
rect 137480 585274 137508 586706
rect 137468 585268 137520 585274
rect 137468 585210 137520 585216
rect 127728 584854 127834 584882
rect 130580 584854 131054 584882
rect 134260 584868 134564 584882
rect 137480 584868 137508 585210
rect 140608 584882 140636 594798
rect 143828 593366 143856 596146
rect 143816 593360 143868 593366
rect 143816 593302 143868 593308
rect 143828 584882 143856 593302
rect 153856 587994 153884 596294
rect 163228 592068 163280 592074
rect 163228 592010 163280 592016
rect 159916 590776 159968 590782
rect 159916 590718 159968 590724
rect 156786 588024 156842 588033
rect 153844 587988 153896 587994
rect 156786 587959 156842 587968
rect 153844 587930 153896 587936
rect 147128 586628 147180 586634
rect 147128 586570 147180 586576
rect 134274 584854 134564 584868
rect 140608 584854 140714 584882
rect 143828 584854 143934 584882
rect 147140 584868 147168 586570
rect 150348 585336 150400 585342
rect 150348 585278 150400 585284
rect 150360 584868 150388 585278
rect 153856 584882 153884 587930
rect 153594 584854 153884 584882
rect 156800 584868 156828 587959
rect 159928 584882 159956 590718
rect 163240 587994 163268 592010
rect 163228 587988 163280 587994
rect 163228 587930 163280 587936
rect 159928 584854 160034 584882
rect 163240 584868 163268 587930
rect 166276 586702 166304 604522
rect 169036 593434 169064 607310
rect 178696 596174 178724 611322
rect 178604 596146 178724 596174
rect 169024 593428 169076 593434
rect 169024 593370 169076 593376
rect 169576 593428 169628 593434
rect 169576 593370 169628 593376
rect 166264 586696 166316 586702
rect 166264 586638 166316 586644
rect 166276 586514 166304 586638
rect 166276 586486 166488 586514
rect 166460 584868 166488 586486
rect 169588 584882 169616 593370
rect 178604 592249 178632 596146
rect 178590 592240 178646 592249
rect 178590 592175 178646 592184
rect 172888 587920 172940 587926
rect 172888 587862 172940 587868
rect 169588 584854 169694 584882
rect 172900 584868 172928 587862
rect 175462 585168 175518 585177
rect 175462 585103 175518 585112
rect 175476 584868 175504 585103
rect 178604 584882 178632 592175
rect 181904 586628 181956 586634
rect 181904 586570 181956 586576
rect 178604 584854 178710 584882
rect 181916 584868 181944 586570
rect 185596 585342 185624 619618
rect 191104 610020 191156 610026
rect 191104 609962 191156 609968
rect 188250 592104 188306 592113
rect 188250 592039 188306 592048
rect 185124 585336 185176 585342
rect 185124 585278 185176 585284
rect 185584 585336 185636 585342
rect 185584 585278 185636 585284
rect 185136 584868 185164 585278
rect 188264 584882 188292 592039
rect 191116 590714 191144 609962
rect 207572 608728 207624 608734
rect 207572 608670 207624 608676
rect 204352 603220 204404 603226
rect 204352 603162 204404 603168
rect 191104 590708 191156 590714
rect 191104 590650 191156 590656
rect 191472 590708 191524 590714
rect 191472 590650 191524 590656
rect 197268 590708 197320 590714
rect 197268 590650 197320 590656
rect 191484 584882 191512 590650
rect 197280 588334 197308 590650
rect 197268 588328 197320 588334
rect 197268 588270 197320 588276
rect 194784 588056 194836 588062
rect 194784 587998 194836 588004
rect 188264 584854 188370 584882
rect 191484 584854 191590 584882
rect 194796 584868 194824 587998
rect 197280 587586 197308 588270
rect 197268 587580 197320 587586
rect 197268 587522 197320 587528
rect 198004 587580 198056 587586
rect 198004 587522 198056 587528
rect 198016 584868 198044 587522
rect 201224 586696 201276 586702
rect 201224 586638 201276 586644
rect 201236 584868 201264 586638
rect 204364 584882 204392 603162
rect 207584 584882 207612 608670
rect 210436 586401 210464 702510
rect 214104 588124 214156 588130
rect 214104 588066 214156 588072
rect 210422 586392 210478 586401
rect 210422 586327 210478 586336
rect 210882 586392 210938 586401
rect 210882 586327 210938 586336
rect 204364 584854 204470 584882
rect 207584 584854 207690 584882
rect 210896 584868 210924 586327
rect 214116 584868 214144 588066
rect 217336 586770 217364 702578
rect 235184 700398 235212 703520
rect 245660 702772 245712 702778
rect 245660 702714 245712 702720
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 220728 620288 220780 620294
rect 220728 620230 220780 620236
rect 220740 596154 220768 620230
rect 236644 618928 236696 618934
rect 236644 618870 236696 618876
rect 229100 617568 229152 617574
rect 229100 617510 229152 617516
rect 227628 616140 227680 616146
rect 227628 616082 227680 616088
rect 223028 610088 223080 610094
rect 223028 610030 223080 610036
rect 220728 596148 220780 596154
rect 220728 596090 220780 596096
rect 217324 586764 217376 586770
rect 217324 586706 217376 586712
rect 217232 586696 217284 586702
rect 217232 586638 217284 586644
rect 217244 585138 217272 586638
rect 217336 586514 217364 586706
rect 220740 586673 220768 596090
rect 220542 586664 220598 586673
rect 220542 586599 220598 586608
rect 220726 586664 220782 586673
rect 220726 586599 220782 586608
rect 217336 586486 217456 586514
rect 217232 585132 217284 585138
rect 217232 585074 217284 585080
rect 217428 584882 217456 586486
rect 217350 584854 217456 584882
rect 220556 584868 220584 586599
rect 223040 584882 223068 610030
rect 227640 585410 227668 616082
rect 229112 615494 229140 617510
rect 229112 615466 229508 615494
rect 229480 614174 229508 615466
rect 229468 614168 229520 614174
rect 229468 614110 229520 614116
rect 226340 585404 226392 585410
rect 226340 585346 226392 585352
rect 227628 585404 227680 585410
rect 227628 585346 227680 585352
rect 223040 584854 223146 584882
rect 226352 584868 226380 585346
rect 229480 584882 229508 614110
rect 232688 608660 232740 608666
rect 232688 608602 232740 608608
rect 232700 584882 232728 608602
rect 236656 597514 236684 618870
rect 236000 597508 236052 597514
rect 236000 597450 236052 597456
rect 236644 597508 236696 597514
rect 236644 597450 236696 597456
rect 236012 596222 236040 597450
rect 236000 596216 236052 596222
rect 236000 596158 236052 596164
rect 229480 584854 229586 584882
rect 232700 584854 232806 584882
rect 236012 584868 236040 596158
rect 244924 586832 244976 586838
rect 244924 586774 244976 586780
rect 239220 586696 239272 586702
rect 239220 586638 239272 586644
rect 239232 584868 239260 586638
rect 243084 586628 243136 586634
rect 243084 586570 243136 586576
rect 64786 584624 64842 584633
rect 64722 584582 64786 584610
rect 64786 584559 64842 584568
rect 242466 584310 243032 584338
rect 243004 580582 243032 584310
rect 242992 580576 243044 580582
rect 242992 580518 243044 580524
rect 242992 579692 243044 579698
rect 242992 579634 243044 579640
rect 63498 579184 63554 579193
rect 63498 579119 63554 579128
rect 243004 567194 243032 579634
rect 242912 567166 243032 567194
rect 63406 471744 63462 471753
rect 63406 471679 63408 471688
rect 63460 471679 63462 471688
rect 63408 471650 63460 471656
rect 63420 471619 63448 471650
rect 63406 435024 63462 435033
rect 63406 434959 63462 434968
rect 63314 414624 63370 414633
rect 63314 414559 63370 414568
rect 63222 411360 63278 411369
rect 63222 411295 63278 411304
rect 63132 401056 63184 401062
rect 63132 400998 63184 401004
rect 62684 383626 62804 383654
rect 62684 376786 62712 383626
rect 62672 376780 62724 376786
rect 62672 376722 62724 376728
rect 62684 376174 62712 376722
rect 62672 376168 62724 376174
rect 62672 376110 62724 376116
rect 63236 348430 63264 411295
rect 63316 398132 63368 398138
rect 63316 398074 63368 398080
rect 63224 348424 63276 348430
rect 63224 348366 63276 348372
rect 62764 294160 62816 294166
rect 62764 294102 62816 294108
rect 62028 252544 62080 252550
rect 62028 252486 62080 252492
rect 61936 235612 61988 235618
rect 61936 235554 61988 235560
rect 61844 207664 61896 207670
rect 61844 207606 61896 207612
rect 60556 182912 60608 182918
rect 60556 182854 60608 182860
rect 57244 164212 57296 164218
rect 57244 164154 57296 164160
rect 62028 121508 62080 121514
rect 62028 121450 62080 121456
rect 62040 86970 62068 121450
rect 62028 86964 62080 86970
rect 62028 86906 62080 86912
rect 62120 66904 62172 66910
rect 62120 66846 62172 66852
rect 53840 62824 53892 62830
rect 53840 62766 53892 62772
rect 51080 50448 51132 50454
rect 51080 50390 51132 50396
rect 48964 45552 49016 45558
rect 48964 45494 49016 45500
rect 46940 40724 46992 40730
rect 46940 40666 46992 40672
rect 46952 16574 46980 40666
rect 48320 35216 48372 35222
rect 48320 35158 48372 35164
rect 48332 16574 48360 35158
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 44192 6886 44312 6914
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50160 15972 50212 15978
rect 50160 15914 50212 15920
rect 50172 480 50200 15914
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 50390
rect 52460 33788 52512 33794
rect 52460 33730 52512 33736
rect 52472 3602 52500 33730
rect 52552 22840 52604 22846
rect 52552 22782 52604 22788
rect 52460 3596 52512 3602
rect 52460 3538 52512 3544
rect 52564 480 52592 22782
rect 53852 16574 53880 62766
rect 56600 54528 56652 54534
rect 56600 54470 56652 54476
rect 56612 16574 56640 54470
rect 60740 47592 60792 47598
rect 60740 47534 60792 47540
rect 59360 44940 59412 44946
rect 59360 44882 59412 44888
rect 57980 19984 58032 19990
rect 57980 19926 58032 19932
rect 57992 16574 58020 19926
rect 53852 16546 54984 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 53380 3596 53432 3602
rect 53380 3538 53432 3544
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3538
rect 54956 480 54984 16546
rect 56048 4820 56100 4826
rect 56048 4762 56100 4768
rect 56060 480 56088 4762
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 44882
rect 60752 16574 60780 47534
rect 62132 16574 62160 66846
rect 62776 59362 62804 294102
rect 63328 260778 63356 398074
rect 63316 260772 63368 260778
rect 63316 260714 63368 260720
rect 62856 258732 62908 258738
rect 62856 258674 62908 258680
rect 62868 238241 62896 258674
rect 63420 256018 63448 434959
rect 63498 418024 63554 418033
rect 63498 417959 63554 417968
rect 63512 384334 63540 417959
rect 140594 405104 140650 405113
rect 64078 405062 64736 405090
rect 64708 398886 64736 405062
rect 66272 405062 66654 405090
rect 68284 405068 68336 405074
rect 64878 404424 64934 404433
rect 64878 404359 64934 404368
rect 64696 398880 64748 398886
rect 64696 398822 64748 398828
rect 63500 384328 63552 384334
rect 63500 384270 63552 384276
rect 64604 288448 64656 288454
rect 64604 288390 64656 288396
rect 63408 256012 63460 256018
rect 63408 255954 63460 255960
rect 63224 247172 63276 247178
rect 63224 247114 63276 247120
rect 62854 238232 62910 238241
rect 62854 238167 62910 238176
rect 63236 191146 63264 247114
rect 63420 242214 63448 255954
rect 64512 252612 64564 252618
rect 64512 252554 64564 252560
rect 63408 242208 63460 242214
rect 63408 242150 63460 242156
rect 63316 241596 63368 241602
rect 63316 241538 63368 241544
rect 63328 221474 63356 241538
rect 64524 229838 64552 252554
rect 64512 229832 64564 229838
rect 64512 229774 64564 229780
rect 63316 221468 63368 221474
rect 63316 221410 63368 221416
rect 64616 220182 64644 288390
rect 64708 239086 64736 398822
rect 64892 289134 64920 404359
rect 66272 383518 66300 405062
rect 68284 405010 68336 405016
rect 69032 405062 69874 405090
rect 71792 405062 73094 405090
rect 66904 403708 66956 403714
rect 66904 403650 66956 403656
rect 66260 383512 66312 383518
rect 66260 383454 66312 383460
rect 66916 367062 66944 403650
rect 67272 383512 67324 383518
rect 67272 383454 67324 383460
rect 67284 382974 67312 383454
rect 67272 382968 67324 382974
rect 67272 382910 67324 382916
rect 66904 367056 66956 367062
rect 66904 366998 66956 367004
rect 66904 333260 66956 333266
rect 66904 333202 66956 333208
rect 65982 297392 66038 297401
rect 65982 297327 66038 297336
rect 64880 289128 64932 289134
rect 64880 289070 64932 289076
rect 64788 270632 64840 270638
rect 64788 270574 64840 270580
rect 64696 239080 64748 239086
rect 64696 239022 64748 239028
rect 64604 220176 64656 220182
rect 64604 220118 64656 220124
rect 63224 191140 63276 191146
rect 63224 191082 63276 191088
rect 63408 127016 63460 127022
rect 63408 126958 63460 126964
rect 63420 95062 63448 126958
rect 63408 95056 63460 95062
rect 63408 94998 63460 95004
rect 64800 82822 64828 270574
rect 65800 248668 65852 248674
rect 65800 248610 65852 248616
rect 65812 233889 65840 248610
rect 65996 246974 66024 297327
rect 66168 273352 66220 273358
rect 66168 273294 66220 273300
rect 66076 271924 66128 271930
rect 66076 271866 66128 271872
rect 65984 246968 66036 246974
rect 65984 246910 66036 246916
rect 65798 233880 65854 233889
rect 65798 233815 65854 233824
rect 66088 205018 66116 271866
rect 66076 205012 66128 205018
rect 66076 204954 66128 204960
rect 66180 181393 66208 273294
rect 66916 252618 66944 333202
rect 66904 252612 66956 252618
rect 66904 252554 66956 252560
rect 67284 241641 67312 382910
rect 68296 358970 68324 405010
rect 68284 358964 68336 358970
rect 68284 358906 68336 358912
rect 68296 352578 68324 358906
rect 68284 352572 68336 352578
rect 68284 352514 68336 352520
rect 68652 340196 68704 340202
rect 68652 340138 68704 340144
rect 68284 309800 68336 309806
rect 68284 309742 68336 309748
rect 67456 299532 67508 299538
rect 67456 299474 67508 299480
rect 67364 295996 67416 296002
rect 67364 295938 67416 295944
rect 67376 278905 67404 295938
rect 67468 279478 67496 299474
rect 68296 291825 68324 309742
rect 68468 298240 68520 298246
rect 68468 298182 68520 298188
rect 68480 291854 68508 298182
rect 68664 291938 68692 340138
rect 69032 308514 69060 405062
rect 71136 401056 71188 401062
rect 71136 400998 71188 401004
rect 71044 399492 71096 399498
rect 71044 399434 71096 399440
rect 69112 380180 69164 380186
rect 69112 380122 69164 380128
rect 69020 308508 69072 308514
rect 69020 308450 69072 308456
rect 68744 303000 68796 303006
rect 68744 302942 68796 302948
rect 68572 291910 68692 291938
rect 68468 291848 68520 291854
rect 68282 291816 68338 291825
rect 68468 291790 68520 291796
rect 68282 291751 68338 291760
rect 67730 291136 67786 291145
rect 67730 291071 67786 291080
rect 67638 290456 67694 290465
rect 67638 290391 67694 290400
rect 67652 289882 67680 290391
rect 67744 289950 67772 291071
rect 67732 289944 67784 289950
rect 67732 289886 67784 289892
rect 67640 289876 67692 289882
rect 67640 289818 67692 289824
rect 67730 289776 67786 289785
rect 67730 289711 67786 289720
rect 67744 289134 67772 289711
rect 67732 289128 67784 289134
rect 67638 289096 67694 289105
rect 67732 289070 67784 289076
rect 67638 289031 67694 289040
rect 67652 288454 67680 289031
rect 67640 288448 67692 288454
rect 67640 288390 67692 288396
rect 67638 287736 67694 287745
rect 67638 287671 67694 287680
rect 67652 287094 67680 287671
rect 67640 287088 67692 287094
rect 67640 287030 67692 287036
rect 67730 287056 67786 287065
rect 67730 286991 67786 287000
rect 67744 285734 67772 286991
rect 67732 285728 67784 285734
rect 67732 285670 67784 285676
rect 68006 284880 68062 284889
rect 68006 284815 68062 284824
rect 67640 284368 67692 284374
rect 67638 284336 67640 284345
rect 67692 284336 67694 284345
rect 67638 284271 67694 284280
rect 67732 284300 67784 284306
rect 67732 284242 67784 284248
rect 67744 282985 67772 284242
rect 68020 283665 68048 284815
rect 68006 283656 68062 283665
rect 68006 283591 68062 283600
rect 67730 282976 67786 282985
rect 67730 282911 67786 282920
rect 68572 281625 68600 291910
rect 68652 291848 68704 291854
rect 68652 291790 68704 291796
rect 68664 285025 68692 291790
rect 68756 285705 68784 302942
rect 69020 295384 69072 295390
rect 69020 295326 69072 295332
rect 68926 290864 68982 290873
rect 68926 290799 68982 290808
rect 68940 286385 68968 290799
rect 68926 286376 68982 286385
rect 68926 286311 68982 286320
rect 68742 285696 68798 285705
rect 68742 285631 68798 285640
rect 68650 285016 68706 285025
rect 68650 284951 68706 284960
rect 68926 283656 68982 283665
rect 68926 283591 68982 283600
rect 68558 281616 68614 281625
rect 68558 281551 68614 281560
rect 67638 280936 67694 280945
rect 67638 280871 67694 280880
rect 67652 280838 67680 280871
rect 67640 280832 67692 280838
rect 67640 280774 67692 280780
rect 67638 280256 67694 280265
rect 67638 280191 67640 280200
rect 67692 280191 67694 280200
rect 67640 280162 67692 280168
rect 67638 279576 67694 279585
rect 67638 279511 67694 279520
rect 67652 279478 67680 279511
rect 67456 279472 67508 279478
rect 67456 279414 67508 279420
rect 67640 279472 67692 279478
rect 67640 279414 67692 279420
rect 67362 278896 67418 278905
rect 67362 278831 67418 278840
rect 67640 278724 67692 278730
rect 67640 278666 67692 278672
rect 67652 278225 67680 278666
rect 67638 278216 67694 278225
rect 67638 278151 67694 278160
rect 67638 277536 67694 277545
rect 67638 277471 67694 277480
rect 67652 277438 67680 277471
rect 67640 277432 67692 277438
rect 67640 277374 67692 277380
rect 67730 276856 67786 276865
rect 67730 276791 67786 276800
rect 67640 276684 67692 276690
rect 67640 276626 67692 276632
rect 67652 276185 67680 276626
rect 67638 276176 67694 276185
rect 67638 276111 67694 276120
rect 67744 276078 67772 276791
rect 67732 276072 67784 276078
rect 67732 276014 67784 276020
rect 67640 276004 67692 276010
rect 67640 275946 67692 275952
rect 67652 275505 67680 275946
rect 67638 275496 67694 275505
rect 67638 275431 67694 275440
rect 68282 274816 68338 274825
rect 68282 274751 68338 274760
rect 67638 274136 67694 274145
rect 67638 274071 67694 274080
rect 67652 273290 67680 274071
rect 67822 273456 67878 273465
rect 67822 273391 67878 273400
rect 67836 273358 67864 273391
rect 67824 273352 67876 273358
rect 67824 273294 67876 273300
rect 67640 273284 67692 273290
rect 67640 273226 67692 273232
rect 67638 272776 67694 272785
rect 67638 272711 67694 272720
rect 67454 272096 67510 272105
rect 67454 272031 67510 272040
rect 67362 250336 67418 250345
rect 67362 250271 67418 250280
rect 67270 241632 67326 241641
rect 67270 241567 67326 241576
rect 67376 220250 67404 250271
rect 67364 220244 67416 220250
rect 67364 220186 67416 220192
rect 67468 192574 67496 272031
rect 67652 271930 67680 272711
rect 67640 271924 67692 271930
rect 67640 271866 67692 271872
rect 67730 271416 67786 271425
rect 67730 271351 67786 271360
rect 67638 270736 67694 270745
rect 67638 270671 67694 270680
rect 67652 270570 67680 270671
rect 67744 270638 67772 271351
rect 67732 270632 67784 270638
rect 67732 270574 67784 270580
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 67732 270496 67784 270502
rect 67732 270438 67784 270444
rect 67638 270056 67694 270065
rect 67638 269991 67694 270000
rect 67652 269142 67680 269991
rect 67744 269385 67772 270438
rect 67730 269376 67786 269385
rect 67730 269311 67786 269320
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 67730 268696 67786 268705
rect 67730 268631 67786 268640
rect 67638 268016 67694 268025
rect 67638 267951 67694 267960
rect 67652 267850 67680 267951
rect 67640 267844 67692 267850
rect 67640 267786 67692 267792
rect 67744 267782 67772 268631
rect 67732 267776 67784 267782
rect 67732 267718 67784 267724
rect 67640 267708 67692 267714
rect 67640 267650 67692 267656
rect 67652 267345 67680 267650
rect 67732 267640 67784 267646
rect 67732 267582 67784 267588
rect 67638 267336 67694 267345
rect 67638 267271 67694 267280
rect 67744 266665 67772 267582
rect 67730 266656 67786 266665
rect 67730 266591 67786 266600
rect 67640 266348 67692 266354
rect 67640 266290 67692 266296
rect 67652 265305 67680 266290
rect 67638 265296 67694 265305
rect 67638 265231 67694 265240
rect 67730 264616 67786 264625
rect 67730 264551 67786 264560
rect 67638 263936 67694 263945
rect 67638 263871 67694 263880
rect 67652 263702 67680 263871
rect 67640 263696 67692 263702
rect 67640 263638 67692 263644
rect 67744 263634 67772 264551
rect 67732 263628 67784 263634
rect 67732 263570 67784 263576
rect 67730 263256 67786 263265
rect 67730 263191 67786 263200
rect 67638 262576 67694 262585
rect 67638 262511 67694 262520
rect 67652 262274 67680 262511
rect 67744 262342 67772 263191
rect 67732 262336 67784 262342
rect 67732 262278 67784 262284
rect 67640 262268 67692 262274
rect 67640 262210 67692 262216
rect 67732 262200 67784 262206
rect 67732 262142 67784 262148
rect 67640 262132 67692 262138
rect 67640 262074 67692 262080
rect 67652 261225 67680 262074
rect 67744 261905 67772 262142
rect 67730 261896 67786 261905
rect 67730 261831 67786 261840
rect 67638 261216 67694 261225
rect 67638 261151 67694 261160
rect 67640 260840 67692 260846
rect 67640 260782 67692 260788
rect 67652 260545 67680 260782
rect 67732 260772 67784 260778
rect 67732 260714 67784 260720
rect 67638 260536 67694 260545
rect 67638 260471 67694 260480
rect 67744 259865 67772 260714
rect 67730 259856 67786 259865
rect 67730 259791 67786 259800
rect 67730 259176 67786 259185
rect 67730 259111 67786 259120
rect 67744 258126 67772 259111
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 67640 258052 67692 258058
rect 67640 257994 67692 258000
rect 67652 257825 67680 257994
rect 67638 257816 67694 257825
rect 67638 257751 67694 257760
rect 67730 256456 67786 256465
rect 67730 256391 67786 256400
rect 67640 256012 67692 256018
rect 67640 255954 67692 255960
rect 67652 255785 67680 255954
rect 67638 255776 67694 255785
rect 67638 255711 67694 255720
rect 67744 255338 67772 256391
rect 67732 255332 67784 255338
rect 67732 255274 67784 255280
rect 67638 255096 67694 255105
rect 67638 255031 67694 255040
rect 67652 254046 67680 255031
rect 67730 254416 67786 254425
rect 67730 254351 67786 254360
rect 67640 254040 67692 254046
rect 67640 253982 67692 253988
rect 67744 253978 67772 254351
rect 67732 253972 67784 253978
rect 67732 253914 67784 253920
rect 67640 253904 67692 253910
rect 67640 253846 67692 253852
rect 67652 253745 67680 253846
rect 67638 253736 67694 253745
rect 67638 253671 67694 253680
rect 67548 252612 67600 252618
rect 67548 252554 67600 252560
rect 67560 252385 67588 252554
rect 67640 252544 67692 252550
rect 67640 252486 67692 252492
rect 67546 252376 67602 252385
rect 67546 252311 67602 252320
rect 67652 251705 67680 252486
rect 68296 251870 68324 274751
rect 68284 251864 68336 251870
rect 68284 251806 68336 251812
rect 67638 251696 67694 251705
rect 67638 251631 67694 251640
rect 67638 251016 67694 251025
rect 67638 250951 67694 250960
rect 67652 249898 67680 250951
rect 67640 249892 67692 249898
rect 67640 249834 67692 249840
rect 67640 249756 67692 249762
rect 67640 249698 67692 249704
rect 67652 249665 67680 249698
rect 67638 249656 67694 249665
rect 67638 249591 67694 249600
rect 68006 248976 68062 248985
rect 68006 248911 68062 248920
rect 68020 248674 68048 248911
rect 68008 248668 68060 248674
rect 68008 248610 68060 248616
rect 67638 248296 67694 248305
rect 67638 248231 67694 248240
rect 67652 247178 67680 248231
rect 67730 247616 67786 247625
rect 67730 247551 67786 247560
rect 67640 247172 67692 247178
rect 67640 247114 67692 247120
rect 67744 247110 67772 247551
rect 67732 247104 67784 247110
rect 67732 247046 67784 247052
rect 67640 247036 67692 247042
rect 67640 246978 67692 246984
rect 67652 246945 67680 246978
rect 68100 246968 68152 246974
rect 67638 246936 67694 246945
rect 68100 246910 68152 246916
rect 67638 246871 67694 246880
rect 68112 246265 68140 246910
rect 68098 246256 68154 246265
rect 68098 246191 68154 246200
rect 67640 245608 67692 245614
rect 67638 245576 67640 245585
rect 67692 245576 67694 245585
rect 67638 245511 67694 245520
rect 67546 244896 67602 244905
rect 67546 244831 67602 244840
rect 67560 206310 67588 244831
rect 67640 244248 67692 244254
rect 67638 244216 67640 244225
rect 67692 244216 67694 244225
rect 67638 244151 67694 244160
rect 67732 244180 67784 244186
rect 67732 244122 67784 244128
rect 67744 243545 67772 244122
rect 67730 243536 67786 243545
rect 67730 243471 67786 243480
rect 67730 242856 67786 242865
rect 67730 242791 67786 242800
rect 67638 242176 67694 242185
rect 67638 242111 67694 242120
rect 67652 241602 67680 242111
rect 67640 241596 67692 241602
rect 67640 241538 67692 241544
rect 67744 241534 67772 242791
rect 67732 241528 67784 241534
rect 67638 241496 67694 241505
rect 67732 241470 67784 241476
rect 67638 241431 67640 241440
rect 67692 241431 67694 241440
rect 67640 241402 67692 241408
rect 67638 240816 67694 240825
rect 67638 240751 67640 240760
rect 67692 240751 67694 240760
rect 67640 240722 67692 240728
rect 67652 235278 67680 240722
rect 67640 235272 67692 235278
rect 67640 235214 67692 235220
rect 68940 210361 68968 283591
rect 69032 265441 69060 295326
rect 69124 288425 69152 380122
rect 70400 360256 70452 360262
rect 70400 360198 70452 360204
rect 70032 294704 70084 294710
rect 70032 294646 70084 294652
rect 70044 291924 70072 294646
rect 70412 294030 70440 360198
rect 71056 303754 71084 399434
rect 71148 360262 71176 400998
rect 71136 360256 71188 360262
rect 71136 360198 71188 360204
rect 70492 303748 70544 303754
rect 70492 303690 70544 303696
rect 71044 303748 71096 303754
rect 71044 303690 71096 303696
rect 70400 294024 70452 294030
rect 70400 293966 70452 293972
rect 70504 291938 70532 303690
rect 71792 295390 71820 405062
rect 75920 404524 75972 404530
rect 75920 404466 75972 404472
rect 75932 402966 75960 404466
rect 75920 402960 75972 402966
rect 75920 402902 75972 402908
rect 73804 402484 73856 402490
rect 73804 402426 73856 402432
rect 73068 307828 73120 307834
rect 73068 307770 73120 307776
rect 72976 298172 73028 298178
rect 72976 298114 73028 298120
rect 71780 295384 71832 295390
rect 71780 295326 71832 295332
rect 71962 295352 72018 295361
rect 72988 295322 73016 298114
rect 73080 295361 73108 307770
rect 73066 295352 73122 295361
rect 71962 295287 72018 295296
rect 72976 295316 73028 295322
rect 71044 294024 71096 294030
rect 71044 293966 71096 293972
rect 71056 291938 71084 293966
rect 70504 291910 70702 291938
rect 71056 291910 71346 291938
rect 71976 291924 72004 295287
rect 73066 295287 73122 295296
rect 72976 295258 73028 295264
rect 73252 294976 73304 294982
rect 73252 294918 73304 294924
rect 72608 294636 72660 294642
rect 72608 294578 72660 294584
rect 72620 291924 72648 294578
rect 73264 291924 73292 294918
rect 73816 294846 73844 402426
rect 76300 400926 76328 405076
rect 79336 405062 79534 405090
rect 81452 405062 82754 405090
rect 79336 402898 79364 405062
rect 79324 402892 79376 402898
rect 79324 402834 79376 402840
rect 76288 400920 76340 400926
rect 76288 400862 76340 400868
rect 75920 399560 75972 399566
rect 75920 399502 75972 399508
rect 75184 398200 75236 398206
rect 75184 398142 75236 398148
rect 74632 329112 74684 329118
rect 74632 329054 74684 329060
rect 74540 301028 74592 301034
rect 74540 300970 74592 300976
rect 73896 295316 73948 295322
rect 73896 295258 73948 295264
rect 73804 294840 73856 294846
rect 73804 294782 73856 294788
rect 73908 291924 73936 295258
rect 74552 291924 74580 300970
rect 74644 294982 74672 329054
rect 75196 306374 75224 398142
rect 75276 329112 75328 329118
rect 75276 329054 75328 329060
rect 75288 328506 75316 329054
rect 75276 328500 75328 328506
rect 75276 328442 75328 328448
rect 75932 307834 75960 399502
rect 79336 385694 79364 402834
rect 80702 402248 80758 402257
rect 80702 402183 80758 402192
rect 79324 385688 79376 385694
rect 79324 385630 79376 385636
rect 78588 341556 78640 341562
rect 78588 341498 78640 341504
rect 78600 309097 78628 341498
rect 79324 311228 79376 311234
rect 79324 311170 79376 311176
rect 77942 309088 77998 309097
rect 77942 309023 77998 309032
rect 78586 309088 78642 309097
rect 78586 309023 78642 309032
rect 77956 307873 77984 309023
rect 77942 307864 77998 307873
rect 75920 307828 75972 307834
rect 77942 307799 77998 307808
rect 75920 307770 75972 307776
rect 75196 306346 75316 306374
rect 74632 294976 74684 294982
rect 74632 294918 74684 294924
rect 75184 294296 75236 294302
rect 75288 294273 75316 306346
rect 76656 305720 76708 305726
rect 76656 305662 76708 305668
rect 75184 294238 75236 294244
rect 75274 294264 75330 294273
rect 75196 291924 75224 294238
rect 75274 294199 75330 294208
rect 75826 294264 75882 294273
rect 75826 294199 75882 294208
rect 75840 291924 75868 294199
rect 76472 294024 76524 294030
rect 76472 293966 76524 293972
rect 76484 291924 76512 293966
rect 76668 291938 76696 305662
rect 77956 294030 77984 307799
rect 79232 300960 79284 300966
rect 79232 300902 79284 300908
rect 78404 294092 78456 294098
rect 78404 294034 78456 294040
rect 77944 294024 77996 294030
rect 77944 293966 77996 293972
rect 77758 292768 77814 292777
rect 77758 292703 77814 292712
rect 76668 291910 77142 291938
rect 77772 291924 77800 292703
rect 78416 291924 78444 294034
rect 79048 293548 79100 293554
rect 79048 293490 79100 293496
rect 79060 292670 79088 293490
rect 79048 292664 79100 292670
rect 79048 292606 79100 292612
rect 79060 291924 79088 292606
rect 79244 291938 79272 300902
rect 79336 293554 79364 311170
rect 80060 306740 80112 306746
rect 80060 306682 80112 306688
rect 79324 293548 79376 293554
rect 79324 293490 79376 293496
rect 80072 291938 80100 306682
rect 80716 296041 80744 402183
rect 81452 318782 81480 405062
rect 82820 402416 82872 402422
rect 82820 402358 82872 402364
rect 82832 322930 82860 402358
rect 83464 402348 83516 402354
rect 83464 402290 83516 402296
rect 83476 364410 83504 402290
rect 84842 400888 84898 400897
rect 84842 400823 84898 400832
rect 83464 364404 83516 364410
rect 83464 364346 83516 364352
rect 81532 322924 81584 322930
rect 81532 322866 81584 322872
rect 82820 322924 82872 322930
rect 82820 322866 82872 322872
rect 81440 318776 81492 318782
rect 81440 318718 81492 318724
rect 81440 303816 81492 303822
rect 81440 303758 81492 303764
rect 80702 296032 80758 296041
rect 80702 295967 80758 295976
rect 81452 294030 81480 303758
rect 81440 294024 81492 294030
rect 81440 293966 81492 293972
rect 80980 292664 81032 292670
rect 80980 292606 81032 292612
rect 79244 291910 79718 291938
rect 80072 291910 80362 291938
rect 80992 291924 81020 292606
rect 81544 291938 81572 322866
rect 83476 306746 83504 364346
rect 83464 306740 83516 306746
rect 83464 306682 83516 306688
rect 84200 298308 84252 298314
rect 84200 298250 84252 298256
rect 83556 296948 83608 296954
rect 83556 296890 83608 296896
rect 82912 295520 82964 295526
rect 82912 295462 82964 295468
rect 81900 294024 81952 294030
rect 81900 293966 81952 293972
rect 81912 291938 81940 293966
rect 81544 291910 81650 291938
rect 81912 291910 82294 291938
rect 82924 291924 82952 295462
rect 83568 291924 83596 296890
rect 84212 291924 84240 298250
rect 84856 296070 84884 400823
rect 85960 396846 85988 405076
rect 88352 405062 89194 405090
rect 86224 400988 86276 400994
rect 86224 400930 86276 400936
rect 85948 396840 86000 396846
rect 85948 396782 86000 396788
rect 86236 311030 86264 400930
rect 88352 394126 88380 405062
rect 88982 399528 89038 399537
rect 88982 399463 89038 399472
rect 88340 394120 88392 394126
rect 88340 394062 88392 394068
rect 87604 319456 87656 319462
rect 87604 319398 87656 319404
rect 87616 315314 87644 319398
rect 87604 315308 87656 315314
rect 87604 315250 87656 315256
rect 85580 311024 85632 311030
rect 85580 310966 85632 310972
rect 86224 311024 86276 311030
rect 86224 310966 86276 310972
rect 85592 306374 85620 310966
rect 86236 310554 86264 310966
rect 86224 310548 86276 310554
rect 86224 310490 86276 310496
rect 88432 307352 88484 307358
rect 88432 307294 88484 307300
rect 85592 306346 86540 306374
rect 84844 296064 84896 296070
rect 84844 296006 84896 296012
rect 84844 294840 84896 294846
rect 84844 294782 84896 294788
rect 84856 291924 84884 294782
rect 85488 294228 85540 294234
rect 85488 294170 85540 294176
rect 85500 291924 85528 294170
rect 86512 291938 86540 306346
rect 88340 305108 88392 305114
rect 88340 305050 88392 305056
rect 86960 299600 87012 299606
rect 86960 299542 87012 299548
rect 86972 291938 87000 299542
rect 88352 294030 88380 305050
rect 88444 302326 88472 307294
rect 88996 305114 89024 399463
rect 89720 396908 89772 396914
rect 89720 396850 89772 396856
rect 89732 307358 89760 396850
rect 92400 375358 92428 405076
rect 95620 396778 95648 405076
rect 98840 400897 98868 405076
rect 98826 400888 98882 400897
rect 98826 400823 98882 400832
rect 102060 398682 102088 405076
rect 104164 403640 104216 403646
rect 104164 403582 104216 403588
rect 104990 403608 105046 403617
rect 102784 401668 102836 401674
rect 102784 401610 102836 401616
rect 100024 398676 100076 398682
rect 100024 398618 100076 398624
rect 102048 398676 102100 398682
rect 102048 398618 102100 398624
rect 95608 396772 95660 396778
rect 95608 396714 95660 396720
rect 95884 392624 95936 392630
rect 95884 392566 95936 392572
rect 92388 375352 92440 375358
rect 92388 375294 92440 375300
rect 93768 375352 93820 375358
rect 93768 375294 93820 375300
rect 90364 374672 90416 374678
rect 90364 374614 90416 374620
rect 89720 307352 89772 307358
rect 89720 307294 89772 307300
rect 90376 307018 90404 374614
rect 93780 374066 93808 375294
rect 93768 374060 93820 374066
rect 93768 374002 93820 374008
rect 91744 357604 91796 357610
rect 91744 357546 91796 357552
rect 89720 307012 89772 307018
rect 89720 306954 89772 306960
rect 90364 307012 90416 307018
rect 90364 306954 90416 306960
rect 88984 305108 89036 305114
rect 88984 305050 89036 305056
rect 88432 302320 88484 302326
rect 88432 302262 88484 302268
rect 88340 294024 88392 294030
rect 88340 293966 88392 293972
rect 88064 292732 88116 292738
rect 88064 292674 88116 292680
rect 86158 291922 86448 291938
rect 86158 291916 86460 291922
rect 86158 291910 86408 291916
rect 86512 291910 86802 291938
rect 86972 291910 87446 291938
rect 88076 291924 88104 292674
rect 88444 291938 88472 302262
rect 89076 294024 89128 294030
rect 89076 293966 89128 293972
rect 89088 291938 89116 293966
rect 89732 291938 89760 306954
rect 90376 306406 90404 306954
rect 90364 306400 90416 306406
rect 90364 306342 90416 306348
rect 90272 302252 90324 302258
rect 90272 302194 90324 302200
rect 90284 291938 90312 302194
rect 91100 300212 91152 300218
rect 91100 300154 91152 300160
rect 91112 291938 91140 300154
rect 91756 294234 91784 357546
rect 93780 308514 93808 374002
rect 95148 362228 95200 362234
rect 95148 362170 95200 362176
rect 93768 308508 93820 308514
rect 93768 308450 93820 308456
rect 95160 306374 95188 362170
rect 95068 306346 95188 306374
rect 95896 306374 95924 392566
rect 98644 384328 98696 384334
rect 98644 384270 98696 384276
rect 96620 365016 96672 365022
rect 96620 364958 96672 364964
rect 96632 364478 96660 364958
rect 96620 364472 96672 364478
rect 96620 364414 96672 364420
rect 95896 306346 96016 306374
rect 93216 297016 93268 297022
rect 93216 296958 93268 296964
rect 91744 294228 91796 294234
rect 91744 294170 91796 294176
rect 91928 294228 91980 294234
rect 91928 294170 91980 294176
rect 88444 291910 88734 291938
rect 89088 291910 89378 291938
rect 89732 291910 90022 291938
rect 90284 291910 90666 291938
rect 91112 291910 91310 291938
rect 91940 291924 91968 294170
rect 92572 292800 92624 292806
rect 92572 292742 92624 292748
rect 92584 292641 92612 292742
rect 92570 292632 92626 292641
rect 92570 292567 92626 292576
rect 92584 291924 92612 292567
rect 93228 291924 93256 296958
rect 93860 296880 93912 296886
rect 93860 296822 93912 296828
rect 93872 291924 93900 296822
rect 95068 295390 95096 306346
rect 95148 296812 95200 296818
rect 95148 296754 95200 296760
rect 94504 295384 94556 295390
rect 94504 295326 94556 295332
rect 95056 295384 95108 295390
rect 95056 295326 95108 295332
rect 94516 291924 94544 295326
rect 95160 291924 95188 296754
rect 95792 294636 95844 294642
rect 95792 294578 95844 294584
rect 95804 291924 95832 294578
rect 95988 292602 96016 306346
rect 96632 294166 96660 364414
rect 98552 303884 98604 303890
rect 98552 303826 98604 303832
rect 97722 296032 97778 296041
rect 97722 295967 97778 295976
rect 97736 295497 97764 295967
rect 97722 295488 97778 295497
rect 97722 295423 97778 295432
rect 96620 294160 96672 294166
rect 96620 294102 96672 294108
rect 95976 292596 96028 292602
rect 95976 292538 96028 292544
rect 95988 291938 96016 292538
rect 96632 291938 96660 294102
rect 95988 291910 96462 291938
rect 96632 291910 97106 291938
rect 97736 291924 97764 295423
rect 98368 293548 98420 293554
rect 98368 293490 98420 293496
rect 98380 292602 98408 293490
rect 98368 292596 98420 292602
rect 98368 292538 98420 292544
rect 98380 291924 98408 292538
rect 98564 291938 98592 303826
rect 98656 293554 98684 384270
rect 100036 370530 100064 398618
rect 100024 370524 100076 370530
rect 100024 370466 100076 370472
rect 101404 365764 101456 365770
rect 101404 365706 101456 365712
rect 98734 364984 98790 364993
rect 98734 364919 98790 364928
rect 98748 303890 98776 364919
rect 98736 303884 98788 303890
rect 98736 303826 98788 303832
rect 101416 298110 101444 365706
rect 102140 306468 102192 306474
rect 102140 306410 102192 306416
rect 102152 303006 102180 306410
rect 102140 303000 102192 303006
rect 102140 302942 102192 302948
rect 101496 299668 101548 299674
rect 101496 299610 101548 299616
rect 101404 298104 101456 298110
rect 101404 298046 101456 298052
rect 100944 295452 100996 295458
rect 100944 295394 100996 295400
rect 98644 293548 98696 293554
rect 98644 293490 98696 293496
rect 99656 292868 99708 292874
rect 99656 292810 99708 292816
rect 98564 291910 99038 291938
rect 99668 291924 99696 292810
rect 100956 291924 100984 295394
rect 101416 291938 101444 298046
rect 101508 294710 101536 299610
rect 102796 296818 102824 401610
rect 103520 303952 103572 303958
rect 103520 303894 103572 303900
rect 102876 297084 102928 297090
rect 102876 297026 102928 297032
rect 102784 296812 102836 296818
rect 102784 296754 102836 296760
rect 101496 294704 101548 294710
rect 101496 294646 101548 294652
rect 102232 294160 102284 294166
rect 102232 294102 102284 294108
rect 101416 291910 101614 291938
rect 102244 291924 102272 294102
rect 102888 291924 102916 297026
rect 103532 291924 103560 303894
rect 103612 301640 103664 301646
rect 103612 301582 103664 301588
rect 103624 294030 103652 301582
rect 104176 298217 104204 403582
rect 104990 403543 105046 403552
rect 105004 304298 105032 403543
rect 105280 401674 105308 405076
rect 108500 402257 108528 405076
rect 108486 402248 108542 402257
rect 108486 402183 108542 402192
rect 105268 401668 105320 401674
rect 105268 401610 105320 401616
rect 111076 399498 111104 405076
rect 113192 405062 114310 405090
rect 111064 399492 111116 399498
rect 111064 399434 111116 399440
rect 113192 385014 113220 405062
rect 117516 402354 117544 405076
rect 120736 404394 120764 405076
rect 122852 405062 123970 405090
rect 127190 405062 127572 405090
rect 117964 404388 118016 404394
rect 117964 404330 118016 404336
rect 120724 404388 120776 404394
rect 120724 404330 120776 404336
rect 117504 402348 117556 402354
rect 117504 402290 117556 402296
rect 116582 391232 116638 391241
rect 116582 391167 116638 391176
rect 113180 385008 113232 385014
rect 113180 384950 113232 384956
rect 114468 385008 114520 385014
rect 114468 384950 114520 384956
rect 114480 384334 114508 384950
rect 114468 384328 114520 384334
rect 114468 384270 114520 384276
rect 111708 378820 111760 378826
rect 111708 378762 111760 378768
rect 110328 370524 110380 370530
rect 110328 370466 110380 370472
rect 109684 356720 109736 356726
rect 109684 356662 109736 356668
rect 106924 331900 106976 331906
rect 106924 331842 106976 331848
rect 106936 318782 106964 331842
rect 106280 318776 106332 318782
rect 106280 318718 106332 318724
rect 106924 318776 106976 318782
rect 106924 318718 106976 318724
rect 105544 316736 105596 316742
rect 105544 316678 105596 316684
rect 104992 304292 105044 304298
rect 104992 304234 105044 304240
rect 105004 303958 105032 304234
rect 104992 303952 105044 303958
rect 104992 303894 105044 303900
rect 105556 299470 105584 316678
rect 106292 306374 106320 318718
rect 109040 313268 109092 313274
rect 109040 313210 109092 313216
rect 109052 312662 109080 313210
rect 109696 312662 109724 356662
rect 109040 312656 109092 312662
rect 109040 312598 109092 312604
rect 109684 312656 109736 312662
rect 109684 312598 109736 312604
rect 106292 306346 107056 306374
rect 106188 303000 106240 303006
rect 106188 302942 106240 302948
rect 105544 299464 105596 299470
rect 105544 299406 105596 299412
rect 106096 299464 106148 299470
rect 106096 299406 106148 299412
rect 106108 298382 106136 299406
rect 106096 298376 106148 298382
rect 106096 298318 106148 298324
rect 104162 298208 104218 298217
rect 104162 298143 104218 298152
rect 103612 294024 103664 294030
rect 103612 293966 103664 293972
rect 104176 291924 104204 298143
rect 104532 294024 104584 294030
rect 104532 293966 104584 293972
rect 104544 291938 104572 293966
rect 105452 292800 105504 292806
rect 105452 292742 105504 292748
rect 104544 291910 104834 291938
rect 105464 291924 105492 292742
rect 106108 291924 106136 298318
rect 106200 292806 106228 302942
rect 106738 295624 106794 295633
rect 106738 295559 106794 295568
rect 106188 292800 106240 292806
rect 106188 292742 106240 292748
rect 106752 291924 106780 295559
rect 107028 291938 107056 306346
rect 107660 301572 107712 301578
rect 107660 301514 107712 301520
rect 107672 291938 107700 301514
rect 108672 299396 108724 299402
rect 108672 299338 108724 299344
rect 107028 291910 107410 291938
rect 107672 291910 108054 291938
rect 108684 291924 108712 299338
rect 109052 294030 109080 312598
rect 110340 302297 110368 370466
rect 109130 302288 109186 302297
rect 109130 302223 109186 302232
rect 110326 302288 110382 302297
rect 110326 302223 110382 302232
rect 109040 294024 109092 294030
rect 109040 293966 109092 293972
rect 109144 291938 109172 302223
rect 111720 299577 111748 378762
rect 113822 370560 113878 370569
rect 113822 370495 113878 370504
rect 112444 369232 112496 369238
rect 112444 369174 112496 369180
rect 111800 303068 111852 303074
rect 111800 303010 111852 303016
rect 110878 299568 110934 299577
rect 110878 299503 110934 299512
rect 111706 299568 111762 299577
rect 111706 299503 111762 299512
rect 109684 294024 109736 294030
rect 109684 293966 109736 293972
rect 109696 291938 109724 293966
rect 110892 291938 110920 299503
rect 111812 299402 111840 303010
rect 111800 299396 111852 299402
rect 111800 299338 111852 299344
rect 112456 297673 112484 369174
rect 113180 360324 113232 360330
rect 113180 360266 113232 360272
rect 112536 355360 112588 355366
rect 112536 355302 112588 355308
rect 112548 305726 112576 355302
rect 112536 305720 112588 305726
rect 112536 305662 112588 305668
rect 112904 298444 112956 298450
rect 112904 298386 112956 298392
rect 112442 297664 112498 297673
rect 112442 297599 112498 297608
rect 111892 294024 111944 294030
rect 111892 293966 111944 293972
rect 109144 291910 109342 291938
rect 109696 291910 109986 291938
rect 110630 291922 110828 291938
rect 110630 291916 110840 291922
rect 110630 291910 110788 291916
rect 86408 291858 86460 291864
rect 110892 291910 111274 291938
rect 111904 291924 111932 293966
rect 112916 291938 112944 298386
rect 112562 291910 112944 291938
rect 113192 291924 113220 360266
rect 113836 306542 113864 370495
rect 114560 308508 114612 308514
rect 114560 308450 114612 308456
rect 113272 306536 113324 306542
rect 113272 306478 113324 306484
rect 113824 306536 113876 306542
rect 113824 306478 113876 306484
rect 113284 306374 113312 306478
rect 113284 306346 114048 306374
rect 113824 295656 113876 295662
rect 113824 295598 113876 295604
rect 113836 291924 113864 295598
rect 114020 291938 114048 306346
rect 114572 294030 114600 308450
rect 114744 304360 114796 304366
rect 114744 304302 114796 304308
rect 114560 294024 114612 294030
rect 114560 293966 114612 293972
rect 114756 291938 114784 304302
rect 116596 300286 116624 391167
rect 116676 369164 116728 369170
rect 116676 369106 116728 369112
rect 116584 300280 116636 300286
rect 116584 300222 116636 300228
rect 116688 296857 116716 369106
rect 117976 362234 118004 404330
rect 121460 402280 121512 402286
rect 121460 402222 121512 402228
rect 119344 400988 119396 400994
rect 119344 400930 119396 400936
rect 118608 385688 118660 385694
rect 118608 385630 118660 385636
rect 118620 385082 118648 385630
rect 118608 385076 118660 385082
rect 118608 385018 118660 385024
rect 117964 362228 118016 362234
rect 117964 362170 118016 362176
rect 117964 356788 118016 356794
rect 117964 356730 118016 356736
rect 116768 315308 116820 315314
rect 116768 315250 116820 315256
rect 116674 296848 116730 296857
rect 116674 296783 116730 296792
rect 115388 294024 115440 294030
rect 115388 293966 115440 293972
rect 115400 291938 115428 293966
rect 116780 292942 116808 315250
rect 117976 306374 118004 356730
rect 118516 345704 118568 345710
rect 118516 345646 118568 345652
rect 118528 345030 118556 345646
rect 118516 345024 118568 345030
rect 118516 344966 118568 344972
rect 117884 306346 118004 306374
rect 117884 303686 117912 306346
rect 117872 303680 117924 303686
rect 117872 303622 117924 303628
rect 117226 297664 117282 297673
rect 117226 297599 117282 297608
rect 117240 294001 117268 297599
rect 117686 294128 117742 294137
rect 117686 294063 117742 294072
rect 117226 293992 117282 294001
rect 117226 293927 117282 293936
rect 116400 292936 116452 292942
rect 116400 292878 116452 292884
rect 116768 292936 116820 292942
rect 116768 292878 116820 292884
rect 114020 291910 114494 291938
rect 114756 291910 115138 291938
rect 115400 291910 115782 291938
rect 116412 291924 116440 292878
rect 117226 292088 117282 292097
rect 117226 292023 117282 292032
rect 117240 291938 117268 292023
rect 117070 291910 117268 291938
rect 117700 291924 117728 294063
rect 117884 291938 117912 303622
rect 118528 295594 118556 344966
rect 118516 295588 118568 295594
rect 118516 295530 118568 295536
rect 118620 291961 118648 385018
rect 119356 306374 119384 400930
rect 120724 398200 120776 398206
rect 120724 398142 120776 398148
rect 120080 367804 120132 367810
rect 120080 367746 120132 367752
rect 119356 306346 119752 306374
rect 119724 295633 119752 306346
rect 119710 295624 119766 295633
rect 119620 295588 119672 295594
rect 119710 295559 119766 295568
rect 119620 295530 119672 295536
rect 118974 293992 119030 294001
rect 118974 293927 119030 293936
rect 118606 291952 118662 291961
rect 117884 291910 118358 291938
rect 118988 291924 119016 293927
rect 119632 291924 119660 295530
rect 118606 291887 118662 291896
rect 110788 291858 110840 291864
rect 69110 288416 69166 288425
rect 69110 288351 69166 288360
rect 119724 267734 119752 295559
rect 120092 278225 120120 367746
rect 120264 305040 120316 305046
rect 120264 304982 120316 304988
rect 120170 291952 120226 291961
rect 120170 291887 120226 291896
rect 120078 278216 120134 278225
rect 120078 278151 120134 278160
rect 119724 267706 119844 267734
rect 69018 265432 69074 265441
rect 69018 265367 69074 265376
rect 69018 258496 69074 258505
rect 69018 258431 69074 258440
rect 68926 210352 68982 210361
rect 68926 210287 68982 210296
rect 67548 206304 67600 206310
rect 67548 206246 67600 206252
rect 67456 192568 67508 192574
rect 67456 192510 67508 192516
rect 66166 181384 66222 181393
rect 66166 181319 66222 181328
rect 69032 175953 69060 258431
rect 119816 249150 119844 267706
rect 120184 261905 120212 291887
rect 120276 286385 120304 304982
rect 120356 294024 120408 294030
rect 120356 293966 120408 293972
rect 120368 291854 120396 293966
rect 120356 291848 120408 291854
rect 120356 291790 120408 291796
rect 120262 286376 120318 286385
rect 120262 286311 120318 286320
rect 120170 261896 120226 261905
rect 120170 261831 120226 261840
rect 120632 251184 120684 251190
rect 120632 251126 120684 251132
rect 120644 251025 120672 251126
rect 120170 251016 120226 251025
rect 120170 250951 120226 250960
rect 120630 251016 120686 251025
rect 120630 250951 120686 250960
rect 119804 249144 119856 249150
rect 119804 249086 119856 249092
rect 119986 248704 120042 248713
rect 119986 248639 120042 248648
rect 120000 242214 120028 248639
rect 69664 242208 69716 242214
rect 69664 242150 69716 242156
rect 119988 242208 120040 242214
rect 119988 242150 120040 242156
rect 69676 219434 69704 242150
rect 120078 241496 120134 241505
rect 120078 241431 120134 241440
rect 119894 241224 119950 241233
rect 119894 241159 119950 241168
rect 119908 240666 119936 241159
rect 119646 240638 119936 240666
rect 70044 239086 70072 240108
rect 70688 239873 70716 240108
rect 70674 239864 70730 239873
rect 70674 239799 70730 239808
rect 70032 239080 70084 239086
rect 70032 239022 70084 239028
rect 71332 219434 71360 240108
rect 71688 239420 71740 239426
rect 71688 239362 71740 239368
rect 71700 238678 71728 239362
rect 71688 238672 71740 238678
rect 71688 238614 71740 238620
rect 71976 233238 72004 240108
rect 72620 238513 72648 240108
rect 73264 238542 73292 240108
rect 73908 238649 73936 240108
rect 73894 238640 73950 238649
rect 74552 238610 74580 240108
rect 75196 238754 75224 240108
rect 74736 238726 75224 238754
rect 73894 238575 73950 238584
rect 74540 238604 74592 238610
rect 74540 238546 74592 238552
rect 73252 238536 73304 238542
rect 72606 238504 72662 238513
rect 73252 238478 73304 238484
rect 72606 238439 72662 238448
rect 74552 237454 74580 238546
rect 74540 237448 74592 237454
rect 74540 237390 74592 237396
rect 71964 233232 72016 233238
rect 71964 233174 72016 233180
rect 72424 233232 72476 233238
rect 72424 233174 72476 233180
rect 69664 219428 69716 219434
rect 69664 219370 69716 219376
rect 70412 219406 71360 219434
rect 70412 196654 70440 219406
rect 70400 196648 70452 196654
rect 70400 196590 70452 196596
rect 72436 188358 72464 233174
rect 74736 215966 74764 238726
rect 75840 238474 75868 240108
rect 75828 238468 75880 238474
rect 75828 238410 75880 238416
rect 75184 237448 75236 237454
rect 75184 237390 75236 237396
rect 74724 215960 74776 215966
rect 74724 215902 74776 215908
rect 72424 188352 72476 188358
rect 72424 188294 72476 188300
rect 75196 182850 75224 237390
rect 76484 233170 76512 240108
rect 77128 237182 77156 240108
rect 77208 238060 77260 238066
rect 77208 238002 77260 238008
rect 77220 237862 77248 238002
rect 77772 237862 77800 240108
rect 77208 237856 77260 237862
rect 77208 237798 77260 237804
rect 77760 237856 77812 237862
rect 77760 237798 77812 237804
rect 77116 237176 77168 237182
rect 77116 237118 77168 237124
rect 77128 236026 77156 237118
rect 76564 236020 76616 236026
rect 76564 235962 76616 235968
rect 77116 236020 77168 236026
rect 77116 235962 77168 235968
rect 76472 233164 76524 233170
rect 76472 233106 76524 233112
rect 76576 198694 76604 235962
rect 77220 212498 77248 237798
rect 78416 231130 78444 240108
rect 79060 237454 79088 240108
rect 79704 238754 79732 240108
rect 80348 239018 80376 240108
rect 80336 239012 80388 239018
rect 80336 238954 80388 238960
rect 80992 238754 81020 240108
rect 81636 238814 81664 240108
rect 79336 238726 79732 238754
rect 80716 238726 81020 238754
rect 81624 238808 81676 238814
rect 81624 238750 81676 238756
rect 79048 237448 79100 237454
rect 79048 237390 79100 237396
rect 79336 235822 79364 238726
rect 79324 235816 79376 235822
rect 79324 235758 79376 235764
rect 78404 231124 78456 231130
rect 78404 231066 78456 231072
rect 77208 212492 77260 212498
rect 77208 212434 77260 212440
rect 79336 200802 79364 235758
rect 80716 233102 80744 238726
rect 81636 238513 81664 238750
rect 81622 238504 81678 238513
rect 80888 238468 80940 238474
rect 81622 238439 81678 238448
rect 80888 238410 80940 238416
rect 80796 237448 80848 237454
rect 80796 237390 80848 237396
rect 80704 233096 80756 233102
rect 80704 233038 80756 233044
rect 79324 200796 79376 200802
rect 79324 200738 79376 200744
rect 76564 198688 76616 198694
rect 76564 198630 76616 198636
rect 80716 185638 80744 233038
rect 80808 192506 80836 237390
rect 80900 223582 80928 238410
rect 82280 238241 82308 240108
rect 82266 238232 82322 238241
rect 82266 238167 82322 238176
rect 82924 237454 82952 240108
rect 82084 237448 82136 237454
rect 82084 237390 82136 237396
rect 82912 237448 82964 237454
rect 82912 237390 82964 237396
rect 80888 223576 80940 223582
rect 80888 223518 80940 223524
rect 82096 222018 82124 237390
rect 83568 233034 83596 240108
rect 84212 238754 84240 240108
rect 84212 238726 84332 238754
rect 84200 233980 84252 233986
rect 84200 233922 84252 233928
rect 83556 233028 83608 233034
rect 83556 232970 83608 232976
rect 82084 222012 82136 222018
rect 82084 221954 82136 221960
rect 83568 219434 83596 232970
rect 83476 219406 83596 219434
rect 83476 213246 83504 219406
rect 83464 213240 83516 213246
rect 83464 213182 83516 213188
rect 84212 204270 84240 233922
rect 84304 205630 84332 238726
rect 84856 233986 84884 240108
rect 84844 233980 84896 233986
rect 84844 233922 84896 233928
rect 85500 219434 85528 240108
rect 85580 238876 85632 238882
rect 85580 238818 85632 238824
rect 85592 238610 85620 238818
rect 85580 238604 85632 238610
rect 85580 238546 85632 238552
rect 86144 237046 86172 240108
rect 86788 238610 86816 240108
rect 87432 238754 87460 240108
rect 86972 238726 87460 238754
rect 86776 238604 86828 238610
rect 86776 238546 86828 238552
rect 86788 238066 86816 238546
rect 86776 238060 86828 238066
rect 86776 238002 86828 238008
rect 86132 237040 86184 237046
rect 86132 236982 86184 236988
rect 84396 219406 85528 219434
rect 84396 210526 84424 219406
rect 86972 213926 87000 238726
rect 88076 224330 88104 240108
rect 88720 237182 88748 240108
rect 89364 237250 89392 240108
rect 90008 238754 90036 240108
rect 89732 238726 90036 238754
rect 89352 237244 89404 237250
rect 89352 237186 89404 237192
rect 88708 237176 88760 237182
rect 88708 237118 88760 237124
rect 88064 224324 88116 224330
rect 88064 224266 88116 224272
rect 86960 213920 87012 213926
rect 86960 213862 87012 213868
rect 84384 210520 84436 210526
rect 84384 210462 84436 210468
rect 84292 205624 84344 205630
rect 84292 205566 84344 205572
rect 84200 204264 84252 204270
rect 84200 204206 84252 204212
rect 89732 202230 89760 238726
rect 90652 219434 90680 240108
rect 91296 238950 91324 240108
rect 91284 238944 91336 238950
rect 91284 238886 91336 238892
rect 91940 238814 91968 240108
rect 91928 238808 91980 238814
rect 91928 238750 91980 238756
rect 92584 219434 92612 240108
rect 93228 235929 93256 240108
rect 93872 238754 93900 240108
rect 93872 238726 94084 238754
rect 93214 235920 93270 235929
rect 93214 235855 93270 235864
rect 93766 235920 93822 235929
rect 93766 235855 93822 235864
rect 89824 219406 90680 219434
rect 92492 219406 92612 219434
rect 89824 206378 89852 219406
rect 89812 206372 89864 206378
rect 89812 206314 89864 206320
rect 89720 202224 89772 202230
rect 89720 202166 89772 202172
rect 92492 198082 92520 219406
rect 92480 198076 92532 198082
rect 92480 198018 92532 198024
rect 93780 198014 93808 235855
rect 93952 231600 94004 231606
rect 93952 231542 94004 231548
rect 93964 223514 93992 231542
rect 93952 223508 94004 223514
rect 93952 223450 94004 223456
rect 94056 199442 94084 238726
rect 94412 235884 94464 235890
rect 94412 235826 94464 235832
rect 94424 229094 94452 235826
rect 94516 231606 94544 240108
rect 95160 235890 95188 240108
rect 95148 235884 95200 235890
rect 95148 235826 95200 235832
rect 95804 234530 95832 240108
rect 95792 234524 95844 234530
rect 95792 234466 95844 234472
rect 96448 233986 96476 240108
rect 97092 238754 97120 240108
rect 96632 238726 97120 238754
rect 95240 233980 95292 233986
rect 95240 233922 95292 233928
rect 96436 233980 96488 233986
rect 96436 233922 96488 233928
rect 94504 231600 94556 231606
rect 94504 231542 94556 231548
rect 94424 229066 94544 229094
rect 94044 199436 94096 199442
rect 94044 199378 94096 199384
rect 93768 198008 93820 198014
rect 93768 197950 93820 197956
rect 94516 197334 94544 229066
rect 95252 209710 95280 233922
rect 95240 209704 95292 209710
rect 95240 209646 95292 209652
rect 94504 197328 94556 197334
rect 94504 197270 94556 197276
rect 96632 192642 96660 238726
rect 97736 219434 97764 240108
rect 98380 233102 98408 240108
rect 99024 238882 99052 240108
rect 99012 238876 99064 238882
rect 99012 238818 99064 238824
rect 98368 233096 98420 233102
rect 98368 233038 98420 233044
rect 98644 229832 98696 229838
rect 98644 229774 98696 229780
rect 96724 219406 97764 219434
rect 96724 215150 96752 219406
rect 96712 215144 96764 215150
rect 96712 215086 96764 215092
rect 98656 195974 98684 229774
rect 99668 220794 99696 240108
rect 100312 234054 100340 240108
rect 100956 238754 100984 240108
rect 100772 238726 100984 238754
rect 100300 234048 100352 234054
rect 100300 233990 100352 233996
rect 99656 220788 99708 220794
rect 99656 220730 99708 220736
rect 98644 195968 98696 195974
rect 98644 195910 98696 195916
rect 100772 194070 100800 238726
rect 101600 221542 101628 240108
rect 102244 233238 102272 240108
rect 102232 233232 102284 233238
rect 102232 233174 102284 233180
rect 101588 221536 101640 221542
rect 101588 221478 101640 221484
rect 102888 219434 102916 240108
rect 103532 238746 103560 240108
rect 103520 238740 103572 238746
rect 103520 238682 103572 238688
rect 103428 233232 103480 233238
rect 103428 233174 103480 233180
rect 102152 219406 102916 219434
rect 102152 207738 102180 219406
rect 102140 207732 102192 207738
rect 102140 207674 102192 207680
rect 100760 194064 100812 194070
rect 100760 194006 100812 194012
rect 96620 192636 96672 192642
rect 96620 192578 96672 192584
rect 80796 192500 80848 192506
rect 80796 192442 80848 192448
rect 80704 185632 80756 185638
rect 80704 185574 80756 185580
rect 100668 184952 100720 184958
rect 100668 184894 100720 184900
rect 75184 182844 75236 182850
rect 75184 182786 75236 182792
rect 99196 178220 99248 178226
rect 99196 178162 99248 178168
rect 97816 178016 97868 178022
rect 97816 177958 97868 177964
rect 97828 176769 97856 177958
rect 99208 176769 99236 178162
rect 100680 177585 100708 184894
rect 103440 184210 103468 233174
rect 104176 232966 104204 240108
rect 104820 233986 104848 240108
rect 104808 233980 104860 233986
rect 104808 233922 104860 233928
rect 104164 232960 104216 232966
rect 104164 232902 104216 232908
rect 104176 222902 104204 232902
rect 105464 227594 105492 240108
rect 106108 238754 106136 240108
rect 106108 238726 106228 238754
rect 106200 231742 106228 238726
rect 106752 237250 106780 240108
rect 107396 237386 107424 240108
rect 108040 238406 108068 240108
rect 108028 238400 108080 238406
rect 108028 238342 108080 238348
rect 107384 237380 107436 237386
rect 107384 237322 107436 237328
rect 106740 237244 106792 237250
rect 106740 237186 106792 237192
rect 106188 231736 106240 231742
rect 106188 231678 106240 231684
rect 106200 231266 106228 231678
rect 106188 231260 106240 231266
rect 106188 231202 106240 231208
rect 105452 227588 105504 227594
rect 105452 227530 105504 227536
rect 104164 222896 104216 222902
rect 104164 222838 104216 222844
rect 108684 219434 108712 240108
rect 109972 238754 110000 240108
rect 109696 238726 110000 238754
rect 109696 235822 109724 238726
rect 109684 235816 109736 235822
rect 109684 235758 109736 235764
rect 107672 219406 108712 219434
rect 107672 206922 107700 219406
rect 107660 206916 107712 206922
rect 107660 206858 107712 206864
rect 107568 189100 107620 189106
rect 107568 189042 107620 189048
rect 106188 187740 106240 187746
rect 106188 187682 106240 187688
rect 103428 184204 103480 184210
rect 103428 184146 103480 184152
rect 106200 177585 106228 187682
rect 107580 177585 107608 189042
rect 109696 184278 109724 235758
rect 110420 232212 110472 232218
rect 110420 232154 110472 232160
rect 110432 200938 110460 232154
rect 110616 219434 110644 240108
rect 111260 232218 111288 240108
rect 111248 232212 111300 232218
rect 111248 232154 111300 232160
rect 110524 219406 110644 219434
rect 110524 206990 110552 219406
rect 111904 217326 111932 240108
rect 112548 238678 112576 240108
rect 112536 238672 112588 238678
rect 112536 238614 112588 238620
rect 113192 234546 113220 240108
rect 113836 235890 113864 240108
rect 114480 238746 114508 240108
rect 114468 238740 114520 238746
rect 114468 238682 114520 238688
rect 115124 238474 115152 240108
rect 115768 238754 115796 240108
rect 115768 238726 115888 238754
rect 115112 238468 115164 238474
rect 115112 238410 115164 238416
rect 115860 237114 115888 238726
rect 115848 237108 115900 237114
rect 115848 237050 115900 237056
rect 113824 235884 113876 235890
rect 113824 235826 113876 235832
rect 113100 234518 113220 234546
rect 113100 233918 113128 234518
rect 113088 233912 113140 233918
rect 113088 233854 113140 233860
rect 111892 217320 111944 217326
rect 111892 217262 111944 217268
rect 110512 206984 110564 206990
rect 110512 206926 110564 206932
rect 111064 206984 111116 206990
rect 111064 206926 111116 206932
rect 110420 200932 110472 200938
rect 110420 200874 110472 200880
rect 109684 184272 109736 184278
rect 109684 184214 109736 184220
rect 110052 179444 110104 179450
rect 110052 179386 110104 179392
rect 100666 177576 100722 177585
rect 100666 177511 100722 177520
rect 106186 177576 106242 177585
rect 106186 177511 106242 177520
rect 107566 177576 107622 177585
rect 107566 177511 107622 177520
rect 108120 176792 108172 176798
rect 97814 176760 97870 176769
rect 97814 176695 97870 176704
rect 99194 176760 99250 176769
rect 99194 176695 99250 176704
rect 100758 176760 100814 176769
rect 100758 176695 100760 176704
rect 100812 176695 100814 176704
rect 108118 176760 108120 176769
rect 110064 176769 110092 179386
rect 108172 176760 108174 176769
rect 108118 176695 108174 176704
rect 110050 176760 110106 176769
rect 110050 176695 110106 176704
rect 100760 176666 100812 176672
rect 104624 176044 104676 176050
rect 104624 175986 104676 175992
rect 69018 175944 69074 175953
rect 69018 175879 69074 175888
rect 104636 175409 104664 175986
rect 111076 175982 111104 206926
rect 113100 191185 113128 233854
rect 115860 192681 115888 237050
rect 116412 219434 116440 240108
rect 116768 239420 116820 239426
rect 116768 239362 116820 239368
rect 116780 237386 116808 239362
rect 117056 238610 117084 240108
rect 117136 239488 117188 239494
rect 117136 239430 117188 239436
rect 117148 238746 117176 239430
rect 117228 238944 117280 238950
rect 117228 238886 117280 238892
rect 117136 238740 117188 238746
rect 117136 238682 117188 238688
rect 117240 238678 117268 238886
rect 117700 238678 117728 240108
rect 117228 238672 117280 238678
rect 117228 238614 117280 238620
rect 117688 238672 117740 238678
rect 117688 238614 117740 238620
rect 117044 238604 117096 238610
rect 117044 238546 117096 238552
rect 118344 238542 118372 240108
rect 118988 238746 119016 240108
rect 119988 239012 120040 239018
rect 119988 238954 120040 238960
rect 118976 238740 119028 238746
rect 118976 238682 119028 238688
rect 118332 238536 118384 238542
rect 118332 238478 118384 238484
rect 120000 238406 120028 238954
rect 119988 238400 120040 238406
rect 119988 238342 120040 238348
rect 116768 237380 116820 237386
rect 116768 237322 116820 237328
rect 117964 234048 118016 234054
rect 117964 233990 118016 233996
rect 115952 219406 116440 219434
rect 115952 203726 115980 219406
rect 115940 203720 115992 203726
rect 115940 203662 115992 203668
rect 117976 199510 118004 233990
rect 120092 215286 120120 241431
rect 120184 229770 120212 250951
rect 120736 237182 120764 398142
rect 121368 305720 121420 305726
rect 121368 305662 121420 305668
rect 121380 305046 121408 305662
rect 121368 305040 121420 305046
rect 121368 304982 121420 304988
rect 121472 287054 121500 402222
rect 122748 384396 122800 384402
rect 122748 384338 122800 384344
rect 122104 367804 122156 367810
rect 122104 367746 122156 367752
rect 121550 291136 121606 291145
rect 121550 291071 121606 291080
rect 121564 289950 121592 291071
rect 121642 290456 121698 290465
rect 121642 290391 121698 290400
rect 121552 289944 121604 289950
rect 121552 289886 121604 289892
rect 121656 289882 121684 290391
rect 121644 289876 121696 289882
rect 121644 289818 121696 289824
rect 121552 289808 121604 289814
rect 121550 289776 121552 289785
rect 121604 289776 121606 289785
rect 121550 289711 121606 289720
rect 121644 289740 121696 289746
rect 121644 289682 121696 289688
rect 121656 289105 121684 289682
rect 121642 289096 121698 289105
rect 121642 289031 121698 289040
rect 121552 288380 121604 288386
rect 121552 288322 121604 288328
rect 121564 287745 121592 288322
rect 121550 287736 121606 287745
rect 121550 287671 121606 287680
rect 121734 287056 121790 287065
rect 121472 287026 121684 287054
rect 121460 285660 121512 285666
rect 121460 285602 121512 285608
rect 121472 284345 121500 285602
rect 121458 284336 121514 284345
rect 121458 284271 121514 284280
rect 121458 283656 121514 283665
rect 121458 283591 121460 283600
rect 121512 283591 121514 283600
rect 121460 283562 121512 283568
rect 121550 282296 121606 282305
rect 121550 282231 121606 282240
rect 121564 281654 121592 282231
rect 121552 281648 121604 281654
rect 121458 281616 121514 281625
rect 121552 281590 121604 281596
rect 121458 281551 121460 281560
rect 121512 281551 121514 281560
rect 121460 281522 121512 281528
rect 121366 280936 121422 280945
rect 121366 280871 121422 280880
rect 120816 272536 120868 272542
rect 120816 272478 120868 272484
rect 120828 238882 120856 272478
rect 121380 268394 121408 280871
rect 121458 280256 121514 280265
rect 121458 280191 121460 280200
rect 121512 280191 121514 280200
rect 121460 280162 121512 280168
rect 121458 278896 121514 278905
rect 121458 278831 121514 278840
rect 121472 278798 121500 278831
rect 121460 278792 121512 278798
rect 121460 278734 121512 278740
rect 121552 278724 121604 278730
rect 121552 278666 121604 278672
rect 121564 277545 121592 278666
rect 121550 277536 121606 277545
rect 121550 277471 121606 277480
rect 121460 277364 121512 277370
rect 121460 277306 121512 277312
rect 121472 276865 121500 277306
rect 121458 276856 121514 276865
rect 121458 276791 121514 276800
rect 121458 276176 121514 276185
rect 121458 276111 121514 276120
rect 121472 276078 121500 276111
rect 121460 276072 121512 276078
rect 121460 276014 121512 276020
rect 121458 275496 121514 275505
rect 121458 275431 121514 275440
rect 121472 274786 121500 275431
rect 121550 274816 121606 274825
rect 121460 274780 121512 274786
rect 121550 274751 121606 274760
rect 121460 274722 121512 274728
rect 121564 274718 121592 274751
rect 121552 274712 121604 274718
rect 121552 274654 121604 274660
rect 121460 274644 121512 274650
rect 121460 274586 121512 274592
rect 121472 274145 121500 274586
rect 121458 274136 121514 274145
rect 121458 274071 121514 274080
rect 121458 273456 121514 273465
rect 121458 273391 121460 273400
rect 121512 273391 121514 273400
rect 121460 273362 121512 273368
rect 121458 272776 121514 272785
rect 121458 272711 121514 272720
rect 121472 272610 121500 272711
rect 121656 272610 121684 287026
rect 121734 286991 121790 287000
rect 121748 286346 121776 286991
rect 121736 286340 121788 286346
rect 121736 286282 121788 286288
rect 121460 272604 121512 272610
rect 121460 272546 121512 272552
rect 121644 272604 121696 272610
rect 121644 272546 121696 272552
rect 121458 271416 121514 271425
rect 121458 271351 121514 271360
rect 121472 270570 121500 271351
rect 121460 270564 121512 270570
rect 121460 270506 121512 270512
rect 121458 270056 121514 270065
rect 121458 269991 121514 270000
rect 121472 269210 121500 269991
rect 121550 269376 121606 269385
rect 121550 269311 121606 269320
rect 121460 269204 121512 269210
rect 121460 269146 121512 269152
rect 121564 269142 121592 269311
rect 121552 269136 121604 269142
rect 121552 269078 121604 269084
rect 121460 269068 121512 269074
rect 121460 269010 121512 269016
rect 121472 268705 121500 269010
rect 121458 268696 121514 268705
rect 121458 268631 121514 268640
rect 121368 268388 121420 268394
rect 121368 268330 121420 268336
rect 121458 268016 121514 268025
rect 121458 267951 121514 267960
rect 121472 267782 121500 267951
rect 121460 267776 121512 267782
rect 121460 267718 121512 267724
rect 122116 266665 122144 367746
rect 122656 362228 122708 362234
rect 122656 362170 122708 362176
rect 122564 291916 122616 291922
rect 122564 291858 122616 291864
rect 122576 287054 122604 291858
rect 122484 287026 122604 287054
rect 122484 285025 122512 287026
rect 122470 285016 122526 285025
rect 122470 284951 122472 284960
rect 122524 284951 122526 284960
rect 122472 284922 122524 284928
rect 122668 279585 122696 362170
rect 122760 291922 122788 384338
rect 122852 303006 122880 405062
rect 126980 399492 127032 399498
rect 126980 399434 127032 399440
rect 125598 387016 125654 387025
rect 125598 386951 125654 386960
rect 125612 386442 125640 386951
rect 125600 386436 125652 386442
rect 125600 386378 125652 386384
rect 125508 369164 125560 369170
rect 125508 369106 125560 369112
rect 122932 337408 122984 337414
rect 122932 337350 122984 337356
rect 122840 303000 122892 303006
rect 122840 302942 122892 302948
rect 122748 291916 122800 291922
rect 122748 291858 122800 291864
rect 122746 285696 122802 285705
rect 122944 285682 122972 337350
rect 124220 313948 124272 313954
rect 124220 313890 124272 313896
rect 123576 295656 123628 295662
rect 123576 295598 123628 295604
rect 122802 285654 122972 285682
rect 122746 285631 122802 285640
rect 122748 284300 122800 284306
rect 122748 284242 122800 284248
rect 122760 282985 122788 284242
rect 122746 282976 122802 282985
rect 122746 282911 122802 282920
rect 122654 279576 122710 279585
rect 122654 279511 122710 279520
rect 122668 279478 122696 279511
rect 122656 279472 122708 279478
rect 122656 279414 122708 279420
rect 122470 278216 122526 278225
rect 122470 278151 122526 278160
rect 122194 272096 122250 272105
rect 122194 272031 122250 272040
rect 122102 266656 122158 266665
rect 122102 266591 122158 266600
rect 121642 265976 121698 265985
rect 121642 265911 121698 265920
rect 121460 265668 121512 265674
rect 121460 265610 121512 265616
rect 121472 265305 121500 265610
rect 121458 265296 121514 265305
rect 121458 265231 121514 265240
rect 121458 263936 121514 263945
rect 121458 263871 121514 263880
rect 121472 263634 121500 263871
rect 121460 263628 121512 263634
rect 121460 263570 121512 263576
rect 121552 263560 121604 263566
rect 121552 263502 121604 263508
rect 121458 263256 121514 263265
rect 121458 263191 121514 263200
rect 121472 262886 121500 263191
rect 121460 262880 121512 262886
rect 121460 262822 121512 262828
rect 121564 262585 121592 263502
rect 121550 262576 121606 262585
rect 121550 262511 121606 262520
rect 121460 262200 121512 262206
rect 121460 262142 121512 262148
rect 120906 261896 120962 261905
rect 120906 261831 120962 261840
rect 120920 249121 120948 261831
rect 121472 261225 121500 262142
rect 121458 261216 121514 261225
rect 121458 261151 121514 261160
rect 121460 260840 121512 260846
rect 121460 260782 121512 260788
rect 121472 260545 121500 260782
rect 121458 260536 121514 260545
rect 121458 260471 121514 260480
rect 121656 260166 121684 265911
rect 121644 260160 121696 260166
rect 121644 260102 121696 260108
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259486 121500 259791
rect 121460 259480 121512 259486
rect 121460 259422 121512 259428
rect 122102 259176 122158 259185
rect 122102 259111 122158 259120
rect 121458 258496 121514 258505
rect 121458 258431 121514 258440
rect 121472 258126 121500 258431
rect 121460 258120 121512 258126
rect 121460 258062 121512 258068
rect 121550 257816 121606 257825
rect 121550 257751 121606 257760
rect 121458 257136 121514 257145
rect 121458 257071 121514 257080
rect 121472 256834 121500 257071
rect 121460 256828 121512 256834
rect 121460 256770 121512 256776
rect 121564 256766 121592 257751
rect 121552 256760 121604 256766
rect 121552 256702 121604 256708
rect 121458 256456 121514 256465
rect 121458 256391 121514 256400
rect 121472 256154 121500 256391
rect 121460 256148 121512 256154
rect 121460 256090 121512 256096
rect 121458 255776 121514 255785
rect 121458 255711 121514 255720
rect 121472 255338 121500 255711
rect 121460 255332 121512 255338
rect 121460 255274 121512 255280
rect 121458 254416 121514 254425
rect 121458 254351 121514 254360
rect 121472 253978 121500 254351
rect 121460 253972 121512 253978
rect 121460 253914 121512 253920
rect 121552 253904 121604 253910
rect 121552 253846 121604 253852
rect 121458 253736 121514 253745
rect 121458 253671 121514 253680
rect 121472 252618 121500 253671
rect 121564 253065 121592 253846
rect 121550 253056 121606 253065
rect 121550 252991 121606 253000
rect 121460 252612 121512 252618
rect 121460 252554 121512 252560
rect 121550 252376 121606 252385
rect 121550 252311 121606 252320
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 251258 121500 251631
rect 121564 251326 121592 252311
rect 121552 251320 121604 251326
rect 121552 251262 121604 251268
rect 121460 251252 121512 251258
rect 121460 251194 121512 251200
rect 121458 250336 121514 250345
rect 121458 250271 121514 250280
rect 121472 249830 121500 250271
rect 121460 249824 121512 249830
rect 121460 249766 121512 249772
rect 121552 249756 121604 249762
rect 121552 249698 121604 249704
rect 121460 249688 121512 249694
rect 121458 249656 121460 249665
rect 121512 249656 121514 249665
rect 121458 249591 121514 249600
rect 120906 249112 120962 249121
rect 120906 249047 120962 249056
rect 121564 248985 121592 249698
rect 121550 248976 121606 248985
rect 121550 248911 121606 248920
rect 121460 248396 121512 248402
rect 121460 248338 121512 248344
rect 121472 247625 121500 248338
rect 121550 248296 121606 248305
rect 121550 248231 121606 248240
rect 121458 247616 121514 247625
rect 121458 247551 121514 247560
rect 121564 247110 121592 248231
rect 121552 247104 121604 247110
rect 121552 247046 121604 247052
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 121458 246256 121514 246265
rect 121458 246191 121514 246200
rect 121472 245750 121500 246191
rect 121564 245818 121592 246871
rect 121552 245812 121604 245818
rect 121552 245754 121604 245760
rect 121460 245744 121512 245750
rect 121460 245686 121512 245692
rect 121460 245608 121512 245614
rect 121460 245550 121512 245556
rect 121550 245576 121606 245585
rect 121472 244905 121500 245550
rect 121550 245511 121606 245520
rect 121458 244896 121514 244905
rect 121458 244831 121514 244840
rect 121564 244322 121592 245511
rect 121552 244316 121604 244322
rect 121552 244258 121604 244264
rect 121644 244248 121696 244254
rect 121458 244216 121514 244225
rect 121644 244190 121696 244196
rect 121458 244151 121460 244160
rect 121512 244151 121514 244160
rect 121460 244122 121512 244128
rect 121656 243545 121684 244190
rect 121642 243536 121698 243545
rect 121642 243471 121698 243480
rect 121460 242888 121512 242894
rect 121458 242856 121460 242865
rect 121512 242856 121514 242865
rect 121458 242791 121514 242800
rect 121552 242820 121604 242826
rect 121552 242762 121604 242768
rect 121564 242185 121592 242762
rect 121550 242176 121606 242185
rect 121550 242111 121606 242120
rect 121458 240816 121514 240825
rect 121458 240751 121514 240760
rect 121472 240174 121500 240751
rect 121460 240168 121512 240174
rect 121460 240110 121512 240116
rect 121642 240136 121698 240145
rect 121642 240071 121698 240080
rect 120816 238876 120868 238882
rect 120816 238818 120868 238824
rect 120724 237176 120776 237182
rect 120724 237118 120776 237124
rect 120172 229764 120224 229770
rect 120172 229706 120224 229712
rect 120080 215280 120132 215286
rect 120080 215222 120132 215228
rect 117964 199504 118016 199510
rect 117964 199446 118016 199452
rect 115846 192672 115902 192681
rect 115846 192607 115902 192616
rect 113086 191176 113142 191185
rect 113086 191111 113142 191120
rect 114468 186380 114520 186386
rect 114468 186322 114520 186328
rect 114374 182200 114430 182209
rect 114374 182135 114430 182144
rect 112628 180872 112680 180878
rect 112628 180814 112680 180820
rect 112640 177585 112668 180814
rect 114388 177585 114416 182135
rect 112626 177576 112682 177585
rect 112626 177511 112682 177520
rect 114374 177576 114430 177585
rect 114374 177511 114430 177520
rect 114480 177313 114508 186322
rect 120736 185706 120764 237118
rect 121656 235929 121684 240071
rect 121642 235920 121698 235929
rect 121642 235855 121698 235864
rect 120724 185700 120776 185706
rect 120724 185642 120776 185648
rect 122116 182170 122144 259111
rect 122208 256086 122236 272031
rect 122286 267336 122342 267345
rect 122286 267271 122342 267280
rect 122196 256080 122248 256086
rect 122196 256022 122248 256028
rect 122194 255096 122250 255105
rect 122194 255031 122250 255040
rect 122208 230489 122236 255031
rect 122194 230480 122250 230489
rect 122194 230415 122250 230424
rect 122300 228478 122328 267271
rect 122484 267034 122512 278151
rect 122760 278050 122788 282911
rect 122748 278044 122800 278050
rect 122748 277986 122800 277992
rect 123484 273420 123536 273426
rect 123484 273362 123536 273368
rect 122472 267028 122524 267034
rect 122472 266970 122524 266976
rect 122470 264616 122526 264625
rect 122470 264551 122526 264560
rect 122484 256018 122512 264551
rect 122472 256012 122524 256018
rect 122472 255954 122524 255960
rect 122288 228472 122340 228478
rect 122288 228414 122340 228420
rect 123496 188562 123524 273362
rect 123588 225690 123616 295598
rect 123668 292936 123720 292942
rect 123668 292878 123720 292884
rect 123680 275330 123708 292878
rect 124232 284306 124260 313890
rect 124864 297016 124916 297022
rect 124864 296958 124916 296964
rect 124310 296848 124366 296857
rect 124310 296783 124366 296792
rect 124324 286346 124352 296783
rect 124312 286340 124364 286346
rect 124312 286282 124364 286288
rect 124220 284300 124272 284306
rect 124220 284242 124272 284248
rect 123668 275324 123720 275330
rect 123668 275266 123720 275272
rect 123668 254040 123720 254046
rect 123668 253982 123720 253988
rect 123680 238610 123708 253982
rect 123668 238604 123720 238610
rect 123668 238546 123720 238552
rect 123576 225684 123628 225690
rect 123576 225626 123628 225632
rect 124876 207874 124904 296958
rect 125140 280832 125192 280838
rect 125140 280774 125192 280780
rect 125048 267096 125100 267102
rect 125048 267038 125100 267044
rect 124956 245812 125008 245818
rect 124956 245754 125008 245760
rect 124864 207868 124916 207874
rect 124864 207810 124916 207816
rect 123484 188556 123536 188562
rect 123484 188498 123536 188504
rect 124968 188494 124996 245754
rect 125060 239018 125088 267038
rect 125048 239012 125100 239018
rect 125048 238954 125100 238960
rect 124956 188488 125008 188494
rect 124956 188430 125008 188436
rect 125060 184278 125088 238954
rect 125152 235822 125180 280774
rect 125520 265674 125548 369106
rect 125612 285666 125640 386378
rect 126244 365016 126296 365022
rect 126244 364958 126296 364964
rect 125600 285660 125652 285666
rect 125600 285602 125652 285608
rect 125508 265668 125560 265674
rect 125508 265610 125560 265616
rect 126256 244186 126284 364958
rect 126428 302932 126480 302938
rect 126428 302874 126480 302880
rect 126336 290488 126388 290494
rect 126336 290430 126388 290436
rect 126244 244180 126296 244186
rect 126244 244122 126296 244128
rect 125140 235816 125192 235822
rect 125140 235758 125192 235764
rect 126348 233034 126376 290430
rect 126440 277438 126468 302874
rect 126428 277432 126480 277438
rect 126428 277374 126480 277380
rect 126888 269000 126940 269006
rect 126888 268942 126940 268948
rect 126900 267782 126928 268942
rect 126888 267776 126940 267782
rect 126888 267718 126940 267724
rect 126336 233028 126388 233034
rect 126336 232970 126388 232976
rect 126244 231124 126296 231130
rect 126244 231066 126296 231072
rect 125784 205624 125836 205630
rect 125782 205592 125784 205601
rect 125836 205592 125838 205601
rect 125782 205527 125838 205536
rect 126256 205086 126284 231066
rect 126900 213314 126928 267718
rect 126888 213308 126940 213314
rect 126888 213250 126940 213256
rect 126888 205624 126940 205630
rect 126888 205566 126940 205572
rect 126244 205080 126296 205086
rect 126244 205022 126296 205028
rect 126900 204338 126928 205566
rect 126888 204332 126940 204338
rect 126888 204274 126940 204280
rect 126992 204270 127020 399434
rect 127544 398818 127572 405062
rect 130396 402286 130424 405076
rect 132512 405062 133630 405090
rect 136652 405062 136850 405090
rect 130384 402280 130436 402286
rect 130384 402222 130436 402228
rect 130396 401674 130424 402222
rect 129648 401668 129700 401674
rect 129648 401610 129700 401616
rect 130384 401668 130436 401674
rect 130384 401610 130436 401616
rect 127532 398812 127584 398818
rect 127532 398754 127584 398760
rect 127544 398206 127572 398754
rect 127532 398200 127584 398206
rect 127532 398142 127584 398148
rect 128360 367056 128412 367062
rect 128360 366998 128412 367004
rect 127072 305652 127124 305658
rect 127072 305594 127124 305600
rect 127084 256154 127112 305594
rect 128372 303074 128400 366998
rect 129004 303884 129056 303890
rect 129004 303826 129056 303832
rect 128360 303068 128412 303074
rect 128360 303010 128412 303016
rect 127164 300144 127216 300150
rect 127164 300086 127216 300092
rect 127176 260846 127204 300086
rect 127164 260840 127216 260846
rect 127164 260782 127216 260788
rect 127440 260840 127492 260846
rect 127440 260782 127492 260788
rect 127452 260234 127480 260782
rect 127440 260228 127492 260234
rect 127440 260170 127492 260176
rect 127072 256148 127124 256154
rect 127072 256090 127124 256096
rect 127084 255406 127112 256090
rect 127072 255400 127124 255406
rect 127072 255342 127124 255348
rect 127624 255400 127676 255406
rect 127624 255342 127676 255348
rect 127636 240786 127664 255342
rect 128360 242956 128412 242962
rect 128360 242898 128412 242904
rect 128372 242826 128400 242898
rect 128360 242820 128412 242826
rect 128360 242762 128412 242768
rect 127624 240780 127676 240786
rect 127624 240722 127676 240728
rect 129016 210458 129044 303826
rect 129188 301504 129240 301510
rect 129188 301446 129240 301452
rect 129096 294092 129148 294098
rect 129096 294034 129148 294040
rect 129108 233034 129136 294034
rect 129200 249694 129228 301446
rect 129188 249688 129240 249694
rect 129188 249630 129240 249636
rect 129188 247104 129240 247110
rect 129188 247046 129240 247052
rect 129096 233028 129148 233034
rect 129096 232970 129148 232976
rect 129004 210452 129056 210458
rect 129004 210394 129056 210400
rect 126980 204264 127032 204270
rect 126980 204206 127032 204212
rect 127440 204264 127492 204270
rect 127440 204206 127492 204212
rect 127452 203590 127480 204206
rect 127440 203584 127492 203590
rect 127440 203526 127492 203532
rect 129200 189922 129228 247046
rect 129660 242962 129688 401610
rect 132408 399560 132460 399566
rect 132408 399502 132460 399508
rect 130382 389872 130438 389881
rect 130382 389807 130438 389816
rect 129740 300280 129792 300286
rect 129740 300222 129792 300228
rect 129752 249762 129780 300222
rect 130396 269006 130424 389807
rect 130568 373312 130620 373318
rect 130568 373254 130620 373260
rect 130476 345704 130528 345710
rect 130476 345646 130528 345652
rect 130384 269000 130436 269006
rect 130384 268942 130436 268948
rect 130384 256080 130436 256086
rect 130384 256022 130436 256028
rect 129740 249756 129792 249762
rect 129740 249698 129792 249704
rect 129752 249082 129780 249698
rect 129740 249076 129792 249082
rect 129740 249018 129792 249024
rect 129648 242956 129700 242962
rect 129648 242898 129700 242904
rect 129188 189916 129240 189922
rect 129188 189858 129240 189864
rect 125048 184272 125100 184278
rect 130396 184249 130424 256022
rect 130488 237046 130516 345646
rect 130580 272542 130608 373254
rect 130660 333328 130712 333334
rect 130660 333270 130712 333276
rect 130672 301646 130700 333270
rect 131856 308440 131908 308446
rect 131856 308382 131908 308388
rect 130660 301640 130712 301646
rect 130660 301582 130712 301588
rect 131764 292868 131816 292874
rect 131764 292810 131816 292816
rect 130568 272536 130620 272542
rect 130568 272478 130620 272484
rect 130568 269204 130620 269210
rect 130568 269146 130620 269152
rect 130476 237040 130528 237046
rect 130476 236982 130528 236988
rect 130580 218822 130608 269146
rect 130660 249144 130712 249150
rect 130660 249086 130712 249092
rect 130568 218816 130620 218822
rect 130568 218758 130620 218764
rect 130672 202434 130700 249086
rect 131776 207806 131804 292810
rect 131868 245682 131896 308382
rect 132420 278730 132448 399502
rect 132512 341562 132540 405062
rect 135904 402280 135956 402286
rect 135904 402222 135956 402228
rect 133880 394052 133932 394058
rect 133880 393994 133932 394000
rect 133144 348424 133196 348430
rect 133144 348366 133196 348372
rect 133156 347818 133184 348366
rect 132592 347812 132644 347818
rect 132592 347754 132644 347760
rect 133144 347812 133196 347818
rect 133144 347754 133196 347760
rect 132500 341556 132552 341562
rect 132500 341498 132552 341504
rect 132500 311160 132552 311166
rect 132500 311102 132552 311108
rect 132408 278724 132460 278730
rect 132408 278666 132460 278672
rect 132420 278118 132448 278666
rect 132408 278112 132460 278118
rect 132408 278054 132460 278060
rect 132512 263566 132540 311102
rect 132500 263560 132552 263566
rect 132500 263502 132552 263508
rect 131948 259480 132000 259486
rect 131948 259422 132000 259428
rect 131856 245676 131908 245682
rect 131856 245618 131908 245624
rect 131868 238746 131896 245618
rect 131856 238740 131908 238746
rect 131856 238682 131908 238688
rect 131960 229838 131988 259422
rect 132604 251190 132632 347754
rect 133144 294228 133196 294234
rect 133144 294170 133196 294176
rect 132592 251184 132644 251190
rect 132592 251126 132644 251132
rect 131948 229832 132000 229838
rect 131948 229774 132000 229780
rect 131764 207800 131816 207806
rect 131764 207742 131816 207748
rect 130660 202428 130712 202434
rect 130660 202370 130712 202376
rect 133156 196722 133184 294170
rect 133892 289746 133920 393994
rect 135916 391406 135944 402222
rect 135904 391400 135956 391406
rect 135904 391342 135956 391348
rect 135904 383104 135956 383110
rect 135904 383046 135956 383052
rect 134616 356176 134668 356182
rect 134616 356118 134668 356124
rect 134524 328500 134576 328506
rect 134524 328442 134576 328448
rect 134536 304434 134564 328442
rect 134524 304428 134576 304434
rect 134524 304370 134576 304376
rect 134524 297084 134576 297090
rect 134524 297026 134576 297032
rect 133880 289740 133932 289746
rect 133880 289682 133932 289688
rect 133328 265736 133380 265742
rect 133328 265678 133380 265684
rect 133236 249824 133288 249830
rect 133236 249766 133288 249772
rect 133248 213382 133276 249766
rect 133340 237114 133368 265678
rect 133788 263560 133840 263566
rect 133788 263502 133840 263508
rect 133800 262857 133828 263502
rect 133786 262848 133842 262857
rect 133786 262783 133842 262792
rect 133328 237108 133380 237114
rect 133328 237050 133380 237056
rect 133236 213376 133288 213382
rect 133236 213318 133288 213324
rect 133144 196716 133196 196722
rect 133144 196658 133196 196664
rect 125048 184214 125100 184220
rect 130382 184240 130438 184249
rect 130382 184175 130438 184184
rect 124128 183592 124180 183598
rect 124128 183534 124180 183540
rect 122104 182164 122156 182170
rect 122104 182106 122156 182112
rect 121184 180940 121236 180946
rect 121184 180882 121236 180888
rect 115848 179648 115900 179654
rect 115848 179590 115900 179596
rect 114466 177304 114522 177313
rect 114466 177239 114522 177248
rect 115860 177177 115888 179590
rect 116952 179580 117004 179586
rect 116952 179522 117004 179528
rect 116964 177177 116992 179522
rect 118424 178288 118476 178294
rect 118424 178230 118476 178236
rect 115846 177168 115902 177177
rect 115846 177103 115902 177112
rect 116950 177168 117006 177177
rect 116950 177103 117006 177112
rect 118436 176769 118464 178230
rect 121196 177585 121224 180882
rect 124140 177585 124168 183534
rect 127808 182232 127860 182238
rect 127808 182174 127860 182180
rect 124956 179716 125008 179722
rect 124956 179658 125008 179664
rect 121182 177576 121238 177585
rect 121182 177511 121238 177520
rect 124126 177576 124182 177585
rect 124126 177511 124182 177520
rect 124968 177177 124996 179658
rect 125784 178084 125836 178090
rect 125784 178026 125836 178032
rect 124954 177168 125010 177177
rect 124954 177103 125010 177112
rect 125796 176769 125824 178026
rect 127820 177585 127848 182174
rect 134536 180169 134564 297026
rect 134628 239494 134656 356118
rect 134708 295520 134760 295526
rect 134708 295462 134760 295468
rect 134616 239488 134668 239494
rect 134616 239430 134668 239436
rect 134720 194138 134748 295462
rect 135168 289740 135220 289746
rect 135168 289682 135220 289688
rect 135180 289105 135208 289682
rect 135166 289096 135222 289105
rect 135166 289031 135222 289040
rect 134800 280220 134852 280226
rect 134800 280162 134852 280168
rect 134708 194132 134760 194138
rect 134708 194074 134760 194080
rect 134812 189854 134840 280162
rect 135916 233170 135944 383046
rect 135994 368656 136050 368665
rect 135994 368591 136050 368600
rect 136008 244254 136036 368591
rect 136088 305108 136140 305114
rect 136088 305050 136140 305056
rect 135996 244248 136048 244254
rect 135996 244190 136048 244196
rect 135904 233164 135956 233170
rect 135904 233106 135956 233112
rect 136100 193866 136128 305050
rect 136180 292732 136232 292738
rect 136180 292674 136232 292680
rect 136088 193860 136140 193866
rect 136088 193802 136140 193808
rect 134800 189848 134852 189854
rect 134800 189790 134852 189796
rect 136192 189786 136220 292674
rect 136652 223514 136680 405062
rect 140056 401713 140084 405076
rect 140594 405039 140650 405048
rect 142172 405062 143290 405090
rect 140042 401704 140098 401713
rect 140042 401639 140098 401648
rect 140608 397390 140636 405039
rect 140596 397384 140648 397390
rect 140596 397326 140648 397332
rect 139308 377460 139360 377466
rect 139308 377402 139360 377408
rect 138020 366376 138072 366382
rect 138020 366318 138072 366324
rect 138032 365838 138060 366318
rect 138020 365832 138072 365838
rect 138020 365774 138072 365780
rect 136732 318096 136784 318102
rect 136732 318038 136784 318044
rect 136744 317490 136772 318038
rect 136732 317484 136784 317490
rect 136732 317426 136784 317432
rect 136744 239426 136772 317426
rect 137284 299668 137336 299674
rect 137284 299610 137336 299616
rect 136732 239420 136784 239426
rect 136732 239362 136784 239368
rect 136640 223508 136692 223514
rect 136640 223450 136692 223456
rect 137100 223508 137152 223514
rect 137100 223450 137152 223456
rect 137112 222970 137140 223450
rect 137100 222964 137152 222970
rect 137100 222906 137152 222912
rect 137296 192710 137324 299610
rect 138032 235890 138060 365774
rect 138664 303816 138716 303822
rect 138664 303758 138716 303764
rect 138020 235884 138072 235890
rect 138020 235826 138072 235832
rect 138676 195362 138704 303758
rect 139320 301578 139348 377402
rect 140044 362296 140096 362302
rect 140044 362238 140096 362244
rect 139308 301572 139360 301578
rect 139308 301514 139360 301520
rect 138756 292664 138808 292670
rect 138756 292606 138808 292612
rect 138664 195356 138716 195362
rect 138664 195298 138716 195304
rect 137284 192704 137336 192710
rect 137284 192646 137336 192652
rect 136180 189780 136232 189786
rect 136180 189722 136232 189728
rect 138768 189689 138796 292606
rect 138848 286408 138900 286414
rect 138848 286350 138900 286356
rect 138860 242894 138888 286350
rect 140056 253910 140084 362238
rect 140136 289944 140188 289950
rect 140136 289886 140188 289892
rect 140044 253904 140096 253910
rect 140044 253846 140096 253852
rect 138848 242888 138900 242894
rect 138848 242830 138900 242836
rect 138754 189680 138810 189689
rect 138754 189615 138810 189624
rect 134616 186448 134668 186454
rect 134616 186390 134668 186396
rect 134522 180160 134578 180169
rect 134522 180095 134578 180104
rect 132040 178424 132092 178430
rect 132040 178366 132092 178372
rect 130752 178152 130804 178158
rect 130752 178094 130804 178100
rect 127806 177576 127862 177585
rect 127806 177511 127862 177520
rect 128176 176860 128228 176866
rect 128176 176802 128228 176808
rect 128188 176769 128216 176802
rect 130764 176769 130792 178094
rect 132052 176769 132080 178366
rect 134628 178022 134656 186390
rect 140148 184346 140176 289886
rect 140608 256698 140636 397326
rect 140688 385688 140740 385694
rect 140688 385630 140740 385636
rect 140596 256692 140648 256698
rect 140596 256634 140648 256640
rect 140608 237250 140636 256634
rect 140596 237244 140648 237250
rect 140596 237186 140648 237192
rect 140608 236706 140636 237186
rect 140596 236700 140648 236706
rect 140596 236642 140648 236648
rect 140700 209710 140728 385630
rect 141516 298308 141568 298314
rect 141516 298250 141568 298256
rect 141424 294296 141476 294302
rect 141424 294238 141476 294244
rect 140688 209704 140740 209710
rect 140688 209646 140740 209652
rect 140700 209166 140728 209646
rect 140688 209160 140740 209166
rect 140688 209102 140740 209108
rect 141436 196790 141464 294238
rect 141528 213450 141556 298250
rect 141608 291848 141660 291854
rect 141608 291790 141660 291796
rect 141620 231198 141648 291790
rect 142172 286414 142200 405062
rect 144920 402348 144972 402354
rect 144920 402290 144972 402296
rect 142804 392012 142856 392018
rect 142804 391954 142856 391960
rect 142816 325694 142844 391954
rect 144184 363044 144236 363050
rect 144184 362986 144236 362992
rect 142816 325666 143028 325694
rect 143000 300937 143028 325666
rect 142986 300928 143042 300937
rect 142986 300863 143042 300872
rect 142804 299600 142856 299606
rect 142804 299542 142856 299548
rect 142160 286408 142212 286414
rect 142160 286350 142212 286356
rect 141608 231192 141660 231198
rect 141608 231134 141660 231140
rect 141516 213444 141568 213450
rect 141516 213386 141568 213392
rect 142816 203794 142844 299542
rect 142896 277432 142948 277438
rect 142896 277374 142948 277380
rect 142908 218006 142936 277374
rect 143000 242350 143028 300863
rect 143080 272604 143132 272610
rect 143080 272546 143132 272552
rect 142988 242344 143040 242350
rect 142988 242286 143040 242292
rect 143092 230382 143120 272546
rect 144196 238814 144224 362986
rect 144276 301572 144328 301578
rect 144276 301514 144328 301520
rect 144184 238808 144236 238814
rect 144184 238750 144236 238756
rect 143080 230376 143132 230382
rect 143080 230318 143132 230324
rect 142896 218000 142948 218006
rect 142896 217942 142948 217948
rect 142804 203788 142856 203794
rect 142804 203730 142856 203736
rect 144288 202366 144316 301514
rect 144368 296948 144420 296954
rect 144368 296890 144420 296896
rect 144380 203930 144408 296890
rect 144460 274780 144512 274786
rect 144460 274722 144512 274728
rect 144472 223446 144500 274722
rect 144460 223440 144512 223446
rect 144460 223382 144512 223388
rect 144932 213926 144960 402290
rect 146496 402082 146524 405076
rect 149072 405062 149730 405090
rect 151832 405062 152950 405090
rect 155972 405062 156170 405090
rect 146484 402076 146536 402082
rect 146484 402018 146536 402024
rect 147680 402076 147732 402082
rect 147680 402018 147732 402024
rect 145564 367192 145616 367198
rect 145564 367134 145616 367140
rect 145576 289814 145604 367134
rect 146944 358896 146996 358902
rect 146944 358838 146996 358844
rect 146298 322960 146354 322969
rect 146298 322895 146300 322904
rect 146352 322895 146354 322904
rect 146300 322866 146352 322872
rect 145656 298376 145708 298382
rect 145656 298318 145708 298324
rect 145564 289808 145616 289814
rect 145564 289750 145616 289756
rect 145564 278792 145616 278798
rect 145564 278734 145616 278740
rect 144920 213920 144972 213926
rect 144920 213862 144972 213868
rect 144368 203924 144420 203930
rect 144368 203866 144420 203872
rect 144276 202360 144328 202366
rect 144276 202302 144328 202308
rect 145576 198218 145604 278734
rect 145668 242282 145696 298318
rect 145656 242276 145708 242282
rect 145656 242218 145708 242224
rect 146956 234530 146984 358838
rect 147588 318096 147640 318102
rect 147588 318038 147640 318044
rect 147600 317490 147628 318038
rect 147588 317484 147640 317490
rect 147588 317426 147640 317432
rect 147036 291236 147088 291242
rect 147036 291178 147088 291184
rect 146944 234524 146996 234530
rect 146944 234466 146996 234472
rect 146208 213920 146260 213926
rect 146208 213862 146260 213868
rect 146220 213518 146248 213862
rect 146208 213512 146260 213518
rect 146208 213454 146260 213460
rect 147048 209302 147076 291178
rect 147494 244352 147550 244361
rect 147494 244287 147496 244296
rect 147548 244287 147550 244296
rect 147496 244258 147548 244264
rect 147036 209296 147088 209302
rect 147036 209238 147088 209244
rect 145564 198212 145616 198218
rect 145564 198154 145616 198160
rect 141424 196784 141476 196790
rect 141424 196726 141476 196732
rect 147508 186998 147536 244258
rect 147600 213246 147628 317426
rect 147692 215286 147720 402018
rect 148324 377596 148376 377602
rect 148324 377538 148376 377544
rect 148336 290494 148364 377538
rect 149072 333266 149100 405062
rect 151084 399492 151136 399498
rect 151084 399434 151136 399440
rect 149060 333260 149112 333266
rect 149060 333202 149112 333208
rect 149796 301028 149848 301034
rect 149796 300970 149848 300976
rect 149704 298444 149756 298450
rect 149704 298386 149756 298392
rect 148508 295384 148560 295390
rect 148508 295326 148560 295332
rect 148324 290488 148376 290494
rect 148324 290430 148376 290436
rect 148324 281648 148376 281654
rect 148324 281590 148376 281596
rect 148336 218890 148364 281590
rect 148416 245744 148468 245750
rect 148416 245686 148468 245692
rect 148324 218884 148376 218890
rect 148324 218826 148376 218832
rect 147680 215280 147732 215286
rect 147680 215222 147732 215228
rect 147692 215150 147720 215222
rect 147680 215144 147732 215150
rect 147680 215086 147732 215092
rect 147588 213240 147640 213246
rect 147588 213182 147640 213188
rect 148428 190058 148456 245686
rect 148520 240106 148548 295326
rect 148508 240100 148560 240106
rect 148508 240042 148560 240048
rect 149716 198150 149744 298386
rect 149704 198144 149756 198150
rect 149704 198086 149756 198092
rect 148416 190052 148468 190058
rect 148416 189994 148468 190000
rect 147496 186992 147548 186998
rect 147496 186934 147548 186940
rect 140136 184340 140188 184346
rect 140136 184282 140188 184288
rect 149808 181665 149836 300970
rect 149980 260228 150032 260234
rect 149980 260170 150032 260176
rect 149888 240168 149940 240174
rect 149888 240110 149940 240116
rect 149900 191214 149928 240110
rect 149992 227730 150020 260170
rect 150072 256828 150124 256834
rect 150072 256770 150124 256776
rect 150084 240922 150112 256770
rect 150072 240916 150124 240922
rect 150072 240858 150124 240864
rect 151096 233238 151124 399434
rect 151832 378894 151860 405062
rect 155868 402280 155920 402286
rect 155868 402222 155920 402228
rect 153200 388544 153252 388550
rect 153200 388486 153252 388492
rect 154120 388544 154172 388550
rect 154120 388486 154172 388492
rect 152556 388476 152608 388482
rect 152556 388418 152608 388424
rect 151820 378888 151872 378894
rect 151820 378830 151872 378836
rect 152464 306400 152516 306406
rect 152464 306342 152516 306348
rect 151176 294160 151228 294166
rect 151176 294102 151228 294108
rect 151084 233232 151136 233238
rect 151084 233174 151136 233180
rect 149980 227724 150032 227730
rect 149980 227666 150032 227672
rect 151188 216034 151216 294102
rect 151360 291304 151412 291310
rect 151360 291246 151412 291252
rect 151268 269136 151320 269142
rect 151268 269078 151320 269084
rect 151176 216028 151228 216034
rect 151176 215970 151228 215976
rect 151280 205154 151308 269078
rect 151372 234054 151400 291246
rect 151360 234048 151412 234054
rect 151360 233990 151412 233996
rect 152476 217977 152504 306342
rect 152568 299538 152596 388418
rect 152924 379500 152976 379506
rect 152924 379442 152976 379448
rect 152936 378894 152964 379442
rect 152924 378888 152976 378894
rect 152924 378830 152976 378836
rect 153108 361684 153160 361690
rect 153108 361626 153160 361632
rect 152556 299532 152608 299538
rect 152556 299474 152608 299480
rect 152568 266354 152596 299474
rect 152648 292800 152700 292806
rect 152648 292742 152700 292748
rect 152660 278186 152688 292742
rect 152648 278180 152700 278186
rect 152648 278122 152700 278128
rect 152740 270564 152792 270570
rect 152740 270506 152792 270512
rect 152556 266348 152608 266354
rect 152556 266290 152608 266296
rect 152648 255332 152700 255338
rect 152648 255274 152700 255280
rect 152660 233170 152688 255274
rect 152648 233164 152700 233170
rect 152648 233106 152700 233112
rect 152462 217968 152518 217977
rect 152462 217903 152518 217912
rect 151268 205148 151320 205154
rect 151268 205090 151320 205096
rect 149888 191208 149940 191214
rect 149888 191150 149940 191156
rect 152752 185774 152780 270506
rect 153120 206990 153148 361626
rect 153212 262886 153240 388486
rect 154132 387938 154160 388486
rect 154120 387932 154172 387938
rect 154120 387874 154172 387880
rect 154488 356244 154540 356250
rect 154488 356186 154540 356192
rect 153844 303748 153896 303754
rect 153844 303690 153896 303696
rect 153200 262880 153252 262886
rect 153200 262822 153252 262828
rect 153856 218754 153884 303690
rect 154394 283520 154450 283529
rect 154394 283455 154450 283464
rect 153936 262880 153988 262886
rect 153936 262822 153988 262828
rect 153948 222154 153976 262822
rect 153936 222148 153988 222154
rect 153936 222090 153988 222096
rect 154408 220114 154436 283455
rect 154396 220108 154448 220114
rect 154396 220050 154448 220056
rect 153844 218748 153896 218754
rect 153844 218690 153896 218696
rect 153108 206984 153160 206990
rect 153108 206926 153160 206932
rect 152740 185768 152792 185774
rect 152740 185710 152792 185716
rect 154500 183054 154528 356186
rect 155776 300824 155828 300830
rect 155776 300766 155828 300772
rect 155224 295452 155276 295458
rect 155224 295394 155276 295400
rect 155236 184385 155264 295394
rect 155316 256012 155368 256018
rect 155316 255954 155368 255960
rect 155328 235822 155356 255954
rect 155788 240854 155816 300766
rect 155776 240848 155828 240854
rect 155776 240790 155828 240796
rect 155316 235816 155368 235822
rect 155316 235758 155368 235764
rect 155880 206922 155908 402222
rect 155972 386306 156000 405062
rect 158732 401674 158760 405076
rect 159364 405068 159416 405074
rect 159364 405010 159416 405016
rect 157984 401668 158036 401674
rect 157984 401610 158036 401616
rect 158720 401668 158772 401674
rect 158720 401610 158772 401616
rect 155960 386300 156012 386306
rect 155960 386242 156012 386248
rect 156420 386300 156472 386306
rect 156420 386242 156472 386248
rect 156432 385694 156460 386242
rect 156420 385688 156472 385694
rect 156420 385630 156472 385636
rect 157996 374134 158024 401610
rect 158628 391264 158680 391270
rect 158628 391206 158680 391212
rect 157984 374128 158036 374134
rect 157984 374070 158036 374076
rect 157248 314696 157300 314702
rect 157248 314638 157300 314644
rect 156602 298208 156658 298217
rect 156602 298143 156658 298152
rect 155868 206916 155920 206922
rect 155868 206858 155920 206864
rect 155880 206446 155908 206858
rect 155868 206440 155920 206446
rect 155868 206382 155920 206388
rect 155222 184376 155278 184385
rect 155222 184311 155278 184320
rect 154488 183048 154540 183054
rect 154488 182990 154540 182996
rect 149794 181656 149850 181665
rect 149794 181591 149850 181600
rect 148232 179512 148284 179518
rect 148232 179454 148284 179460
rect 134616 178016 134668 178022
rect 134616 177958 134668 177964
rect 148244 177177 148272 179454
rect 156616 177313 156644 298143
rect 157156 286408 157208 286414
rect 157156 286350 157208 286356
rect 156696 258120 156748 258126
rect 156696 258062 156748 258068
rect 156708 237250 156736 258062
rect 156696 237244 156748 237250
rect 156696 237186 156748 237192
rect 157168 228410 157196 286350
rect 157260 239465 157288 314638
rect 157996 311234 158024 374070
rect 157984 311228 158036 311234
rect 157984 311170 158036 311176
rect 157984 302320 158036 302326
rect 157984 302262 158036 302268
rect 157246 239456 157302 239465
rect 157246 239391 157302 239400
rect 157156 228404 157208 228410
rect 157156 228346 157208 228352
rect 156696 220244 156748 220250
rect 156696 220186 156748 220192
rect 156708 181490 156736 220186
rect 157996 182986 158024 302262
rect 158168 296744 158220 296750
rect 158168 296686 158220 296692
rect 158076 281580 158128 281586
rect 158076 281522 158128 281528
rect 158088 205222 158116 281522
rect 158180 261526 158208 296686
rect 158640 284306 158668 391206
rect 159376 300830 159404 405010
rect 161952 397322 161980 405076
rect 164252 405062 165186 405090
rect 161940 397316 161992 397322
rect 161940 397258 161992 397264
rect 162768 397316 162820 397322
rect 162768 397258 162820 397264
rect 160744 393372 160796 393378
rect 160744 393314 160796 393320
rect 159456 306536 159508 306542
rect 159456 306478 159508 306484
rect 159364 300824 159416 300830
rect 159364 300766 159416 300772
rect 159364 296880 159416 296886
rect 159364 296822 159416 296828
rect 158628 284300 158680 284306
rect 158628 284242 158680 284248
rect 158640 283529 158668 284242
rect 158626 283520 158682 283529
rect 158626 283455 158682 283464
rect 158720 272536 158772 272542
rect 158720 272478 158772 272484
rect 158732 271930 158760 272478
rect 158720 271924 158772 271930
rect 158720 271866 158772 271872
rect 158168 261520 158220 261526
rect 158168 261462 158220 261468
rect 158628 261520 158680 261526
rect 158628 261462 158680 261468
rect 158168 252612 158220 252618
rect 158168 252554 158220 252560
rect 158180 231130 158208 252554
rect 158258 240136 158314 240145
rect 158258 240071 158314 240080
rect 158272 233238 158300 240071
rect 158640 239494 158668 261462
rect 158628 239488 158680 239494
rect 158628 239430 158680 239436
rect 158260 233232 158312 233238
rect 158260 233174 158312 233180
rect 158168 231124 158220 231130
rect 158168 231066 158220 231072
rect 158168 228540 158220 228546
rect 158168 228482 158220 228488
rect 158076 205216 158128 205222
rect 158076 205158 158128 205164
rect 158180 200025 158208 228482
rect 158166 200016 158222 200025
rect 158166 199951 158222 199960
rect 159376 185745 159404 296822
rect 159468 243574 159496 306478
rect 160100 275324 160152 275330
rect 160100 275266 160152 275272
rect 160112 274786 160140 275266
rect 160100 274780 160152 274786
rect 160100 274722 160152 274728
rect 160008 271924 160060 271930
rect 160008 271866 160060 271872
rect 159548 251320 159600 251326
rect 159548 251262 159600 251268
rect 159456 243568 159508 243574
rect 159456 243510 159508 243516
rect 159560 235754 159588 251262
rect 159548 235748 159600 235754
rect 159548 235690 159600 235696
rect 160020 226302 160048 271866
rect 160756 269074 160784 393314
rect 160836 374672 160888 374678
rect 160836 374614 160888 374620
rect 160848 298246 160876 374614
rect 160928 374128 160980 374134
rect 160928 374070 160980 374076
rect 160940 371958 160968 374070
rect 160928 371952 160980 371958
rect 160928 371894 160980 371900
rect 162780 362982 162808 397258
rect 163504 396840 163556 396846
rect 163504 396782 163556 396788
rect 162308 362976 162360 362982
rect 162308 362918 162360 362924
rect 162768 362976 162820 362982
rect 162768 362918 162820 362924
rect 162124 357740 162176 357746
rect 162124 357682 162176 357688
rect 160928 306468 160980 306474
rect 160928 306410 160980 306416
rect 160836 298240 160888 298246
rect 160836 298182 160888 298188
rect 160848 284374 160876 298182
rect 160836 284368 160888 284374
rect 160836 284310 160888 284316
rect 160836 279472 160888 279478
rect 160836 279414 160888 279420
rect 160744 269068 160796 269074
rect 160744 269010 160796 269016
rect 160008 226296 160060 226302
rect 160008 226238 160060 226244
rect 160848 188426 160876 279414
rect 160940 216578 160968 306410
rect 161296 274780 161348 274786
rect 161296 274722 161348 274728
rect 161308 239426 161336 274722
rect 161388 267776 161440 267782
rect 161388 267718 161440 267724
rect 161296 239420 161348 239426
rect 161296 239362 161348 239368
rect 160928 216572 160980 216578
rect 160928 216514 160980 216520
rect 161400 191282 161428 267718
rect 162136 248402 162164 357682
rect 162216 302252 162268 302258
rect 162216 302194 162268 302200
rect 162124 248396 162176 248402
rect 162124 248338 162176 248344
rect 162124 242956 162176 242962
rect 162124 242898 162176 242904
rect 162136 234462 162164 242898
rect 162124 234456 162176 234462
rect 162124 234398 162176 234404
rect 162228 211954 162256 302194
rect 162320 301510 162348 362918
rect 162308 301504 162360 301510
rect 162308 301446 162360 301452
rect 162768 284368 162820 284374
rect 162768 284310 162820 284316
rect 162308 256760 162360 256766
rect 162308 256702 162360 256708
rect 162216 211948 162268 211954
rect 162216 211890 162268 211896
rect 162320 195430 162348 256702
rect 162780 219366 162808 284310
rect 163516 265742 163544 396782
rect 164252 376718 164280 405062
rect 168288 403776 168340 403782
rect 168288 403718 168340 403724
rect 168196 395344 168248 395350
rect 168196 395286 168248 395292
rect 166816 389836 166868 389842
rect 166816 389778 166868 389784
rect 164240 376712 164292 376718
rect 164240 376654 164292 376660
rect 164884 376712 164936 376718
rect 164884 376654 164936 376660
rect 164896 376106 164924 376654
rect 164884 376100 164936 376106
rect 164884 376042 164936 376048
rect 164148 355496 164200 355502
rect 164148 355438 164200 355444
rect 164160 291174 164188 355438
rect 164896 297401 164924 376042
rect 166632 359576 166684 359582
rect 166632 359518 166684 359524
rect 166264 358828 166316 358834
rect 166264 358770 166316 358776
rect 164976 300960 165028 300966
rect 164976 300902 165028 300908
rect 164882 297392 164938 297401
rect 164882 297327 164938 297336
rect 163688 291168 163740 291174
rect 163688 291110 163740 291116
rect 164148 291168 164200 291174
rect 164148 291110 164200 291116
rect 163700 290494 163728 291110
rect 163688 290488 163740 290494
rect 163688 290430 163740 290436
rect 163596 286340 163648 286346
rect 163596 286282 163648 286288
rect 163504 265736 163556 265742
rect 163504 265678 163556 265684
rect 163608 240825 163636 286282
rect 163700 280838 163728 290430
rect 163688 280832 163740 280838
rect 163688 280774 163740 280780
rect 164884 278112 164936 278118
rect 164884 278054 164936 278060
rect 163688 268388 163740 268394
rect 163688 268330 163740 268336
rect 163594 240816 163650 240825
rect 163594 240751 163650 240760
rect 163700 236774 163728 268330
rect 164148 254040 164200 254046
rect 164148 253982 164200 253988
rect 164056 245676 164108 245682
rect 164056 245618 164108 245624
rect 163688 236768 163740 236774
rect 163688 236710 163740 236716
rect 162768 219360 162820 219366
rect 162768 219302 162820 219308
rect 164068 216646 164096 245618
rect 164056 216640 164108 216646
rect 164056 216582 164108 216588
rect 164160 212430 164188 253982
rect 164148 212424 164200 212430
rect 164148 212366 164200 212372
rect 162308 195424 162360 195430
rect 162308 195366 162360 195372
rect 161388 191276 161440 191282
rect 161388 191218 161440 191224
rect 162124 189984 162176 189990
rect 162124 189926 162176 189932
rect 160836 188420 160888 188426
rect 160836 188362 160888 188368
rect 159362 185736 159418 185745
rect 159362 185671 159418 185680
rect 157984 182980 158036 182986
rect 157984 182922 158036 182928
rect 156696 181484 156748 181490
rect 156696 181426 156748 181432
rect 159272 178356 159324 178362
rect 159272 178298 159324 178304
rect 156602 177304 156658 177313
rect 156602 177239 156658 177248
rect 148230 177168 148286 177177
rect 148230 177103 148286 177112
rect 134432 176928 134484 176934
rect 134432 176870 134484 176876
rect 134444 176769 134472 176870
rect 159284 176769 159312 178298
rect 118422 176760 118478 176769
rect 118422 176695 118478 176704
rect 125782 176760 125838 176769
rect 125782 176695 125838 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 130750 176760 130806 176769
rect 130750 176695 130806 176704
rect 132038 176760 132094 176769
rect 132038 176695 132094 176704
rect 134430 176760 134486 176769
rect 134430 176695 134486 176704
rect 135718 176760 135774 176769
rect 135718 176695 135774 176704
rect 159270 176760 159326 176769
rect 159270 176695 159326 176704
rect 135732 176662 135760 176695
rect 135720 176656 135772 176662
rect 135720 176598 135772 176604
rect 133144 176248 133196 176254
rect 133144 176190 133196 176196
rect 129464 176180 129516 176186
rect 129464 176122 129516 176128
rect 121920 176112 121972 176118
rect 121920 176054 121972 176060
rect 111064 175976 111116 175982
rect 111064 175918 111116 175924
rect 119436 175976 119488 175982
rect 119436 175918 119488 175924
rect 104622 175400 104678 175409
rect 104622 175335 104678 175344
rect 119448 175001 119476 175918
rect 121932 175409 121960 176054
rect 129476 175409 129504 176122
rect 133156 175409 133184 176190
rect 162136 176089 162164 189926
rect 164896 187066 164924 278054
rect 164988 214577 165016 300902
rect 165066 295488 165122 295497
rect 165066 295423 165122 295432
rect 165080 229770 165108 295423
rect 166276 292641 166304 358770
rect 166262 292632 166318 292641
rect 166262 292567 166318 292576
rect 166276 282878 166304 292567
rect 166264 282872 166316 282878
rect 166264 282814 166316 282820
rect 166264 276072 166316 276078
rect 166264 276014 166316 276020
rect 165528 269816 165580 269822
rect 165528 269758 165580 269764
rect 165540 269249 165568 269758
rect 165526 269240 165582 269249
rect 165526 269175 165582 269184
rect 165068 229764 165120 229770
rect 165068 229706 165120 229712
rect 165540 228313 165568 269175
rect 165526 228304 165582 228313
rect 165526 228239 165582 228248
rect 164974 214568 165030 214577
rect 164974 214503 165030 214512
rect 164884 187060 164936 187066
rect 164884 187002 164936 187008
rect 165252 178424 165304 178430
rect 165252 178366 165304 178372
rect 164516 176928 164568 176934
rect 164516 176870 164568 176876
rect 162122 176080 162178 176089
rect 162122 176015 162178 176024
rect 121918 175400 121974 175409
rect 121918 175335 121974 175344
rect 129462 175400 129518 175409
rect 129462 175335 129518 175344
rect 133142 175400 133198 175409
rect 133142 175335 133198 175344
rect 164528 175166 164556 176870
rect 164516 175160 164568 175166
rect 164516 175102 164568 175108
rect 119434 174992 119490 175001
rect 119434 174927 119490 174936
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 65522 128072 65578 128081
rect 65522 128007 65578 128016
rect 65536 127022 65564 128007
rect 65524 127016 65576 127022
rect 65524 126958 65576 126964
rect 66074 122632 66130 122641
rect 66074 122567 66130 122576
rect 66088 121514 66116 122567
rect 66076 121508 66128 121514
rect 66076 121450 66128 121456
rect 66074 102368 66130 102377
rect 66074 102303 66130 102312
rect 66088 89690 66116 102303
rect 66180 93838 66208 129231
rect 67638 126304 67694 126313
rect 67638 126239 67694 126248
rect 67546 125216 67602 125225
rect 67546 125151 67602 125160
rect 67454 123584 67510 123593
rect 67454 123519 67510 123528
rect 67362 120864 67418 120873
rect 67362 120799 67418 120808
rect 67270 100736 67326 100745
rect 67270 100671 67326 100680
rect 66168 93832 66220 93838
rect 66168 93774 66220 93780
rect 67284 91050 67312 100671
rect 67272 91044 67324 91050
rect 67272 90986 67324 90992
rect 67376 89729 67404 120799
rect 67468 90982 67496 123519
rect 67456 90976 67508 90982
rect 67456 90918 67508 90924
rect 67362 89720 67418 89729
rect 66076 89684 66128 89690
rect 67362 89655 67418 89664
rect 66076 89626 66128 89632
rect 67560 85542 67588 125151
rect 67548 85536 67600 85542
rect 67548 85478 67600 85484
rect 64788 82816 64840 82822
rect 64788 82758 64840 82764
rect 63500 76560 63552 76566
rect 63500 76502 63552 76508
rect 62764 59356 62816 59362
rect 62764 59298 62816 59304
rect 63512 16574 63540 76502
rect 67652 74526 67680 126239
rect 165264 173874 165292 178366
rect 166276 178022 166304 276014
rect 166644 255270 166672 359518
rect 166828 358834 166856 389778
rect 166908 381540 166960 381546
rect 166908 381482 166960 381488
rect 166816 358828 166868 358834
rect 166816 358770 166868 358776
rect 166724 278180 166776 278186
rect 166724 278122 166776 278128
rect 166736 277438 166764 278122
rect 166724 277432 166776 277438
rect 166724 277374 166776 277380
rect 166632 255264 166684 255270
rect 166632 255206 166684 255212
rect 166644 254046 166672 255206
rect 166632 254040 166684 254046
rect 166632 253982 166684 253988
rect 166736 235890 166764 277374
rect 166724 235884 166776 235890
rect 166724 235826 166776 235832
rect 166920 231742 166948 381482
rect 168208 356153 168236 395286
rect 168194 356144 168250 356153
rect 168194 356079 168250 356088
rect 167000 355428 167052 355434
rect 167000 355370 167052 355376
rect 167012 354754 167040 355370
rect 167000 354748 167052 354754
rect 167000 354690 167052 354696
rect 167012 245614 167040 354690
rect 167736 304292 167788 304298
rect 167736 304234 167788 304240
rect 167092 299464 167144 299470
rect 167092 299406 167144 299412
rect 167104 298790 167132 299406
rect 167092 298784 167144 298790
rect 167092 298726 167144 298732
rect 167644 289876 167696 289882
rect 167644 289818 167696 289824
rect 167000 245608 167052 245614
rect 167000 245550 167052 245556
rect 166908 231736 166960 231742
rect 166908 231678 166960 231684
rect 166448 179716 166500 179722
rect 166448 179658 166500 179664
rect 166356 178288 166408 178294
rect 166356 178230 166408 178236
rect 166264 178016 166316 178022
rect 166264 177958 166316 177964
rect 165528 176248 165580 176254
rect 165528 176190 165580 176196
rect 165540 175234 165568 176190
rect 166172 176180 166224 176186
rect 166172 176122 166224 176128
rect 165528 175228 165580 175234
rect 165528 175170 165580 175176
rect 165252 173868 165304 173874
rect 165252 173810 165304 173816
rect 166184 172514 166212 176122
rect 166264 176112 166316 176118
rect 166264 176054 166316 176060
rect 166172 172508 166224 172514
rect 166172 172450 166224 172456
rect 166276 168366 166304 176054
rect 166264 168360 166316 168366
rect 166264 168302 166316 168308
rect 166368 167006 166396 178230
rect 166460 169726 166488 179658
rect 167656 177342 167684 289818
rect 167748 231334 167776 304234
rect 168208 299470 168236 356079
rect 168196 299464 168248 299470
rect 168196 299406 168248 299412
rect 168300 294642 168328 403718
rect 168392 398954 168420 405076
rect 171612 404394 171640 405076
rect 171600 404388 171652 404394
rect 171600 404330 171652 404336
rect 169024 403640 169076 403646
rect 169024 403582 169076 403588
rect 168380 398948 168432 398954
rect 168380 398890 168432 398896
rect 168288 294636 168340 294642
rect 168288 294578 168340 294584
rect 168300 294001 168328 294578
rect 168286 293992 168342 294001
rect 168286 293927 168342 293936
rect 169036 267102 169064 403582
rect 172428 402348 172480 402354
rect 172428 402290 172480 402296
rect 169760 398948 169812 398954
rect 169760 398890 169812 398896
rect 169772 398750 169800 398890
rect 169760 398744 169812 398750
rect 169760 398686 169812 398692
rect 169772 398290 169800 398686
rect 169588 398262 169800 398290
rect 169116 357536 169168 357542
rect 169116 357478 169168 357484
rect 169128 296002 169156 357478
rect 169116 295996 169168 296002
rect 169116 295938 169168 295944
rect 169116 284980 169168 284986
rect 169116 284922 169168 284928
rect 169024 267096 169076 267102
rect 169024 267038 169076 267044
rect 167828 260160 167880 260166
rect 167828 260102 167880 260108
rect 167736 231328 167788 231334
rect 167736 231270 167788 231276
rect 167840 226234 167868 260102
rect 167828 226228 167880 226234
rect 167828 226170 167880 226176
rect 168932 220788 168984 220794
rect 168932 220730 168984 220736
rect 168944 220250 168972 220730
rect 168932 220244 168984 220250
rect 168932 220186 168984 220192
rect 167920 182232 167972 182238
rect 167920 182174 167972 182180
rect 167736 180872 167788 180878
rect 167736 180814 167788 180820
rect 167644 177336 167696 177342
rect 167644 177278 167696 177284
rect 167000 176860 167052 176866
rect 167000 176802 167052 176808
rect 167012 172446 167040 176802
rect 167000 172440 167052 172446
rect 167000 172382 167052 172388
rect 166448 169720 166500 169726
rect 166448 169662 166500 169668
rect 166356 167000 166408 167006
rect 166356 166942 166408 166948
rect 167748 164218 167776 180814
rect 167828 179648 167880 179654
rect 167828 179590 167880 179596
rect 167840 165578 167868 179590
rect 167932 171086 167960 182174
rect 169128 180130 169156 284922
rect 169208 278044 169260 278050
rect 169208 277986 169260 277992
rect 169220 224806 169248 277986
rect 169300 267028 169352 267034
rect 169300 266970 169352 266976
rect 169312 233918 169340 266970
rect 169300 233912 169352 233918
rect 169300 233854 169352 233860
rect 169208 224800 169260 224806
rect 169208 224742 169260 224748
rect 169588 220250 169616 398262
rect 171048 392692 171100 392698
rect 171048 392634 171100 392640
rect 170956 359508 171008 359514
rect 170956 359450 171008 359456
rect 170496 357672 170548 357678
rect 170496 357614 170548 357620
rect 169760 333940 169812 333946
rect 169760 333882 169812 333888
rect 169772 333334 169800 333882
rect 169760 333328 169812 333334
rect 169760 333270 169812 333276
rect 170404 310548 170456 310554
rect 170404 310490 170456 310496
rect 169576 220244 169628 220250
rect 169576 220186 169628 220192
rect 170416 202298 170444 310490
rect 170508 274650 170536 357614
rect 170588 356108 170640 356114
rect 170588 356050 170640 356056
rect 170600 298178 170628 356050
rect 170968 333946 170996 359450
rect 170956 333940 171008 333946
rect 170956 333882 171008 333888
rect 171060 312594 171088 392634
rect 172336 373380 172388 373386
rect 172336 373322 172388 373328
rect 171784 370660 171836 370666
rect 171784 370602 171836 370608
rect 171140 356312 171192 356318
rect 171140 356254 171192 356260
rect 171152 353258 171180 356254
rect 171140 353252 171192 353258
rect 171140 353194 171192 353200
rect 170680 312588 170732 312594
rect 170680 312530 170732 312536
rect 171048 312588 171100 312594
rect 171048 312530 171100 312536
rect 170692 300218 170720 312530
rect 170680 300212 170732 300218
rect 170680 300154 170732 300160
rect 170588 298172 170640 298178
rect 170588 298114 170640 298120
rect 170600 288318 170628 298114
rect 170588 288312 170640 288318
rect 170588 288254 170640 288260
rect 170588 274712 170640 274718
rect 170588 274654 170640 274660
rect 170496 274644 170548 274650
rect 170496 274586 170548 274592
rect 170496 242208 170548 242214
rect 170496 242150 170548 242156
rect 170404 202292 170456 202298
rect 170404 202234 170456 202240
rect 170404 184952 170456 184958
rect 170404 184894 170456 184900
rect 169208 183592 169260 183598
rect 169208 183534 169260 183540
rect 169116 180124 169168 180130
rect 169116 180066 169168 180072
rect 169024 176792 169076 176798
rect 169024 176734 169076 176740
rect 168010 171592 168066 171601
rect 168010 171527 168066 171536
rect 168024 171154 168052 171527
rect 168012 171148 168064 171154
rect 168012 171090 168064 171096
rect 167920 171080 167972 171086
rect 167920 171022 167972 171028
rect 167828 165572 167880 165578
rect 167828 165514 167880 165520
rect 167736 164212 167788 164218
rect 167736 164154 167788 164160
rect 169036 161430 169064 176734
rect 169220 169658 169248 183534
rect 169300 180940 169352 180946
rect 169300 180882 169352 180888
rect 169208 169652 169260 169658
rect 169208 169594 169260 169600
rect 169312 168298 169340 180882
rect 169300 168292 169352 168298
rect 169300 168234 169352 168240
rect 169024 161424 169076 161430
rect 169024 161366 169076 161372
rect 170416 157350 170444 184894
rect 170508 180033 170536 242150
rect 170600 223038 170628 274654
rect 171152 262206 171180 353194
rect 171796 349858 171824 370602
rect 171784 349852 171836 349858
rect 171784 349794 171836 349800
rect 172348 306134 172376 373322
rect 172336 306128 172388 306134
rect 172336 306070 172388 306076
rect 172348 305726 172376 306070
rect 172336 305720 172388 305726
rect 172336 305662 172388 305668
rect 172336 296948 172388 296954
rect 172336 296890 172388 296896
rect 172348 296818 172376 296890
rect 172336 296812 172388 296818
rect 172336 296754 172388 296760
rect 171876 263628 171928 263634
rect 171876 263570 171928 263576
rect 171140 262200 171192 262206
rect 171140 262142 171192 262148
rect 170680 251252 170732 251258
rect 170680 251194 170732 251200
rect 170692 239601 170720 251194
rect 171784 243568 171836 243574
rect 171784 243510 171836 243516
rect 170678 239592 170734 239601
rect 170678 239527 170734 239536
rect 170588 223032 170640 223038
rect 170588 222974 170640 222980
rect 170680 222964 170732 222970
rect 170680 222906 170732 222912
rect 170692 211818 170720 222906
rect 170680 211812 170732 211818
rect 170680 211754 170732 211760
rect 171796 209234 171824 243510
rect 171888 229906 171916 263570
rect 172348 237386 172376 296754
rect 172336 237380 172388 237386
rect 172336 237322 172388 237328
rect 171876 229900 171928 229906
rect 171876 229842 171928 229848
rect 172440 227594 172468 402290
rect 174832 399498 174860 405076
rect 178052 404462 178080 405076
rect 181286 405062 181484 405090
rect 178040 404456 178092 404462
rect 178040 404398 178092 404404
rect 174820 399492 174872 399498
rect 174820 399434 174872 399440
rect 173164 395412 173216 395418
rect 173164 395354 173216 395360
rect 173176 283626 173204 395354
rect 178052 394398 178080 404398
rect 181456 402966 181484 405062
rect 183572 405062 184506 405090
rect 181444 402960 181496 402966
rect 181444 402902 181496 402908
rect 178040 394392 178092 394398
rect 178040 394334 178092 394340
rect 178684 394392 178736 394398
rect 178684 394334 178736 394340
rect 178696 393378 178724 394334
rect 179328 394052 179380 394058
rect 179328 393994 179380 394000
rect 178684 393372 178736 393378
rect 178684 393314 178736 393320
rect 178696 383042 178724 393314
rect 178684 383036 178736 383042
rect 178684 382978 178736 382984
rect 176568 381608 176620 381614
rect 176568 381550 176620 381556
rect 176382 373280 176438 373289
rect 176382 373215 176438 373224
rect 176290 371920 176346 371929
rect 176290 371855 176346 371864
rect 173716 365084 173768 365090
rect 173716 365026 173768 365032
rect 173728 345710 173756 365026
rect 175186 362264 175242 362273
rect 175186 362199 175242 362208
rect 175096 361616 175148 361622
rect 175096 361558 175148 361564
rect 173808 355428 173860 355434
rect 173808 355370 173860 355376
rect 173716 345704 173768 345710
rect 173716 345646 173768 345652
rect 173256 325712 173308 325718
rect 173256 325654 173308 325660
rect 173268 318102 173296 325654
rect 173256 318096 173308 318102
rect 173256 318038 173308 318044
rect 173820 310282 173848 355370
rect 174544 354816 174596 354822
rect 174544 354758 174596 354764
rect 173348 310276 173400 310282
rect 173348 310218 173400 310224
rect 173808 310276 173860 310282
rect 173808 310218 173860 310224
rect 173256 304428 173308 304434
rect 173256 304370 173308 304376
rect 173164 283620 173216 283626
rect 173164 283562 173216 283568
rect 173164 253972 173216 253978
rect 173164 253914 173216 253920
rect 172428 227588 172480 227594
rect 172428 227530 172480 227536
rect 172440 227050 172468 227530
rect 172428 227044 172480 227050
rect 172428 226986 172480 226992
rect 171784 209228 171836 209234
rect 171784 209170 171836 209176
rect 171508 187128 171560 187134
rect 171508 187070 171560 187076
rect 171520 182889 171548 187070
rect 173176 183122 173204 253914
rect 173268 220318 173296 304370
rect 173360 304366 173388 310218
rect 173348 304360 173400 304366
rect 173348 304302 173400 304308
rect 173348 294024 173400 294030
rect 173348 293966 173400 293972
rect 173360 286414 173388 293966
rect 174556 288386 174584 354758
rect 175108 345014 175136 361558
rect 175016 344986 175136 345014
rect 175016 340882 175044 344986
rect 175004 340876 175056 340882
rect 175004 340818 175056 340824
rect 175016 337414 175044 340818
rect 175096 338156 175148 338162
rect 175096 338098 175148 338104
rect 175004 337408 175056 337414
rect 175004 337350 175056 337356
rect 174544 288380 174596 288386
rect 174544 288322 174596 288328
rect 173348 286408 173400 286414
rect 173348 286350 173400 286356
rect 174636 284368 174688 284374
rect 174636 284310 174688 284316
rect 173348 283620 173400 283626
rect 173348 283562 173400 283568
rect 173360 238882 173388 283562
rect 174648 280158 174676 284310
rect 174636 280152 174688 280158
rect 174636 280094 174688 280100
rect 174544 265668 174596 265674
rect 174544 265610 174596 265616
rect 173348 238876 173400 238882
rect 173348 238818 173400 238824
rect 173256 220312 173308 220318
rect 173256 220254 173308 220260
rect 173164 183116 173216 183122
rect 173164 183058 173216 183064
rect 171506 182880 171562 182889
rect 171506 182815 171562 182824
rect 170494 180024 170550 180033
rect 170494 179959 170550 179968
rect 173164 179580 173216 179586
rect 173164 179522 173216 179528
rect 171784 178220 171836 178226
rect 171784 178162 171836 178168
rect 170496 176044 170548 176050
rect 170496 175986 170548 175992
rect 170508 160070 170536 175986
rect 170588 175976 170640 175982
rect 170588 175918 170640 175924
rect 170600 166938 170628 175918
rect 170588 166932 170640 166938
rect 170588 166874 170640 166880
rect 170496 160064 170548 160070
rect 170496 160006 170548 160012
rect 170404 157344 170456 157350
rect 170404 157286 170456 157292
rect 171796 155922 171824 178162
rect 171876 176724 171928 176730
rect 171876 176666 171928 176672
rect 171888 159390 171916 176666
rect 173176 166870 173204 179522
rect 173164 166864 173216 166870
rect 173164 166806 173216 166812
rect 171876 159384 171928 159390
rect 171876 159326 171928 159332
rect 171784 155916 171836 155922
rect 171784 155858 171836 155864
rect 171784 145036 171836 145042
rect 171784 144978 171836 144984
rect 166264 144968 166316 144974
rect 166264 144910 166316 144916
rect 164884 98048 164936 98054
rect 164884 97990 164936 97996
rect 151726 94888 151782 94897
rect 151726 94823 151782 94832
rect 94962 94752 95018 94761
rect 94962 94687 95018 94696
rect 113178 94752 113234 94761
rect 113178 94687 113234 94696
rect 115846 94752 115902 94761
rect 115846 94687 115902 94696
rect 126518 94752 126574 94761
rect 126518 94687 126574 94696
rect 94976 93906 95004 94687
rect 113192 94042 113220 94687
rect 115860 94110 115888 94687
rect 115848 94104 115900 94110
rect 115848 94046 115900 94052
rect 113180 94036 113232 94042
rect 113180 93978 113232 93984
rect 126532 93974 126560 94687
rect 126520 93968 126572 93974
rect 126520 93910 126572 93916
rect 94964 93900 95016 93906
rect 94964 93842 95016 93848
rect 130750 93664 130806 93673
rect 130750 93599 130806 93608
rect 97262 93528 97318 93537
rect 97262 93463 97318 93472
rect 113822 93528 113878 93537
rect 113822 93463 113878 93472
rect 97276 93226 97304 93463
rect 113836 93294 113864 93463
rect 130764 93430 130792 93599
rect 130752 93424 130804 93430
rect 130752 93366 130804 93372
rect 151740 93362 151768 94823
rect 151728 93356 151780 93362
rect 151728 93298 151780 93304
rect 113824 93288 113876 93294
rect 110142 93256 110198 93265
rect 97264 93220 97316 93226
rect 113824 93230 113876 93236
rect 110142 93191 110198 93200
rect 97264 93162 97316 93168
rect 98184 92472 98236 92478
rect 87142 92440 87198 92449
rect 87142 92375 87198 92384
rect 98182 92440 98184 92449
rect 98236 92440 98238 92449
rect 98182 92375 98238 92384
rect 98642 92440 98698 92449
rect 98642 92375 98698 92384
rect 107382 92440 107438 92449
rect 107382 92375 107438 92384
rect 75366 91216 75422 91225
rect 75366 91151 75422 91160
rect 85486 91216 85542 91225
rect 85486 91151 85542 91160
rect 86406 91216 86462 91225
rect 86406 91151 86462 91160
rect 86866 91216 86922 91225
rect 86866 91151 86922 91160
rect 75380 88330 75408 91151
rect 75368 88324 75420 88330
rect 75368 88266 75420 88272
rect 75920 76628 75972 76634
rect 75920 76570 75972 76576
rect 67640 74520 67692 74526
rect 67640 74462 67692 74468
rect 69020 71052 69072 71058
rect 69020 70994 69072 71000
rect 64880 69692 64932 69698
rect 64880 69634 64932 69640
rect 64892 16574 64920 69634
rect 67640 50380 67692 50386
rect 67640 50322 67692 50328
rect 66260 31136 66312 31142
rect 66260 31078 66312 31084
rect 66272 16574 66300 31078
rect 60752 16546 61608 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 60832 6180 60884 6186
rect 60832 6122 60884 6128
rect 60844 480 60872 6122
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 50322
rect 69032 16574 69060 70994
rect 74540 69760 74592 69766
rect 74540 69702 74592 69708
rect 70400 62892 70452 62898
rect 70400 62834 70452 62840
rect 70412 16574 70440 62834
rect 71780 61396 71832 61402
rect 71780 61338 71832 61344
rect 71792 16574 71820 61338
rect 73160 53168 73212 53174
rect 73160 53110 73212 53116
rect 73172 16574 73200 53110
rect 74552 16574 74580 69702
rect 69032 16546 69152 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69124 480 69152 16546
rect 69848 15904 69900 15910
rect 69848 15846 69900 15852
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 15846
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 76570
rect 85500 75886 85528 91151
rect 86420 88262 86448 91151
rect 86408 88256 86460 88262
rect 86408 88198 86460 88204
rect 86880 78606 86908 91151
rect 87156 91118 87184 92375
rect 89626 91216 89682 91225
rect 89626 91151 89682 91160
rect 90638 91216 90694 91225
rect 90638 91151 90694 91160
rect 92386 91216 92442 91225
rect 92386 91151 92442 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97906 91216 97962 91225
rect 98656 91186 98684 92375
rect 99746 91760 99802 91769
rect 99746 91695 99802 91704
rect 99286 91216 99342 91225
rect 97906 91151 97962 91160
rect 98644 91180 98696 91186
rect 87144 91112 87196 91118
rect 87144 91054 87196 91060
rect 89640 79830 89668 91151
rect 90652 85474 90680 91151
rect 90640 85468 90692 85474
rect 90640 85410 90692 85416
rect 92400 80034 92428 91151
rect 93780 81394 93808 91151
rect 95160 83978 95188 91151
rect 96540 84046 96568 91151
rect 96528 84040 96580 84046
rect 96528 83982 96580 83988
rect 95148 83972 95200 83978
rect 95148 83914 95200 83920
rect 97920 82550 97948 91151
rect 99286 91151 99342 91160
rect 98644 91122 98696 91128
rect 97908 82544 97960 82550
rect 97908 82486 97960 82492
rect 93768 81388 93820 81394
rect 93768 81330 93820 81336
rect 92388 80028 92440 80034
rect 92388 79970 92440 79976
rect 89628 79824 89680 79830
rect 89628 79766 89680 79772
rect 99300 78674 99328 91151
rect 99760 89554 99788 91695
rect 101954 91352 102010 91361
rect 101954 91287 102010 91296
rect 104806 91352 104862 91361
rect 104806 91287 104862 91296
rect 100666 91216 100722 91225
rect 100666 91151 100722 91160
rect 101678 91216 101734 91225
rect 101678 91151 101734 91160
rect 99748 89548 99800 89554
rect 99748 89490 99800 89496
rect 100680 81190 100708 91151
rect 101692 85513 101720 91151
rect 101678 85504 101734 85513
rect 101678 85439 101734 85448
rect 101968 84114 101996 91287
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 102966 91216 103022 91225
rect 102966 91151 103022 91160
rect 103334 91216 103390 91225
rect 103334 91151 103390 91160
rect 104714 91216 104770 91225
rect 104714 91151 104770 91160
rect 101956 84108 102008 84114
rect 101956 84050 102008 84056
rect 100668 81184 100720 81190
rect 100668 81126 100720 81132
rect 102060 80073 102088 91151
rect 102980 86698 103008 91151
rect 103348 86834 103376 91151
rect 103336 86828 103388 86834
rect 103336 86770 103388 86776
rect 102968 86692 103020 86698
rect 102968 86634 103020 86640
rect 104728 84182 104756 91151
rect 104716 84176 104768 84182
rect 104716 84118 104768 84124
rect 102046 80064 102102 80073
rect 102046 79999 102102 80008
rect 99288 78668 99340 78674
rect 99288 78610 99340 78616
rect 86868 78600 86920 78606
rect 86868 78542 86920 78548
rect 85488 75880 85540 75886
rect 85488 75822 85540 75828
rect 104820 73166 104848 91287
rect 107396 91254 107424 92375
rect 108946 91352 109002 91361
rect 108946 91287 109002 91296
rect 107384 91248 107436 91254
rect 105726 91216 105782 91225
rect 107384 91190 107436 91196
rect 107474 91216 107530 91225
rect 105726 91151 105782 91160
rect 107474 91151 107530 91160
rect 108854 91216 108910 91225
rect 108854 91151 108910 91160
rect 105740 88194 105768 91151
rect 105728 88188 105780 88194
rect 105728 88130 105780 88136
rect 107488 81122 107516 91151
rect 108868 82754 108896 91151
rect 108856 82748 108908 82754
rect 108856 82690 108908 82696
rect 108960 82618 108988 91287
rect 109774 91216 109830 91225
rect 109774 91151 109830 91160
rect 109788 88233 109816 91151
rect 110156 90846 110184 93191
rect 121460 93152 121512 93158
rect 121460 93094 121512 93100
rect 121472 92478 121500 93094
rect 121460 92472 121512 92478
rect 116766 92440 116822 92449
rect 116766 92375 116822 92384
rect 120354 92440 120410 92449
rect 125784 92472 125836 92478
rect 121460 92414 121512 92420
rect 124034 92440 124090 92449
rect 120354 92375 120356 92384
rect 116780 92342 116808 92375
rect 120408 92375 120410 92384
rect 124034 92375 124090 92384
rect 125782 92440 125784 92449
rect 125836 92440 125838 92449
rect 125782 92375 125838 92384
rect 129462 92440 129518 92449
rect 129462 92375 129518 92384
rect 133142 92440 133198 92449
rect 133142 92375 133198 92384
rect 135718 92440 135774 92449
rect 135718 92375 135774 92384
rect 151542 92440 151598 92449
rect 151542 92375 151598 92384
rect 152094 92440 152150 92449
rect 152094 92375 152150 92384
rect 120356 92346 120408 92352
rect 116768 92336 116820 92342
rect 116768 92278 116820 92284
rect 117134 91760 117190 91769
rect 117134 91695 117190 91704
rect 110326 91624 110382 91633
rect 110326 91559 110382 91568
rect 110144 90840 110196 90846
rect 110144 90782 110196 90788
rect 110340 89486 110368 91559
rect 112442 91352 112498 91361
rect 112442 91287 112498 91296
rect 111062 91216 111118 91225
rect 111062 91151 111118 91160
rect 111706 91216 111762 91225
rect 111706 91151 111762 91160
rect 110328 89480 110380 89486
rect 110328 89422 110380 89428
rect 109774 88224 109830 88233
rect 109774 88159 109830 88168
rect 111076 85406 111104 91151
rect 111064 85400 111116 85406
rect 111064 85342 111116 85348
rect 108948 82612 109000 82618
rect 108948 82554 109000 82560
rect 111720 81258 111748 91151
rect 112456 86902 112484 91287
rect 113086 91216 113142 91225
rect 113086 91151 113142 91160
rect 115294 91216 115350 91225
rect 115294 91151 115350 91160
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 116584 91180 116636 91186
rect 112444 86896 112496 86902
rect 112444 86838 112496 86844
rect 111708 81252 111760 81258
rect 111708 81194 111760 81200
rect 107476 81116 107528 81122
rect 107476 81058 107528 81064
rect 113100 77178 113128 91151
rect 115308 85270 115336 91151
rect 115296 85264 115348 85270
rect 115296 85206 115348 85212
rect 115860 79966 115888 91151
rect 116584 91122 116636 91128
rect 115848 79960 115900 79966
rect 115848 79902 115900 79908
rect 116596 77246 116624 91122
rect 117148 89622 117176 91695
rect 122838 91488 122894 91497
rect 122838 91423 122894 91432
rect 119344 91248 119396 91254
rect 118054 91216 118110 91225
rect 118054 91151 118110 91160
rect 118606 91216 118662 91225
rect 119344 91190 119396 91196
rect 119894 91216 119950 91225
rect 118606 91151 118662 91160
rect 117136 89616 117188 89622
rect 117136 89558 117188 89564
rect 118068 86766 118096 91151
rect 118056 86760 118108 86766
rect 118056 86702 118108 86708
rect 118620 83910 118648 91151
rect 118608 83904 118660 83910
rect 118608 83846 118660 83852
rect 116584 77240 116636 77246
rect 116584 77182 116636 77188
rect 113088 77172 113140 77178
rect 113088 77114 113140 77120
rect 119356 75818 119384 91190
rect 119894 91151 119950 91160
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 121918 91216 121974 91225
rect 121918 91151 121974 91160
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 119908 88058 119936 91151
rect 119896 88052 119948 88058
rect 119896 87994 119948 88000
rect 121380 87990 121408 91151
rect 121368 87984 121420 87990
rect 121368 87926 121420 87932
rect 121932 85338 121960 91151
rect 121920 85332 121972 85338
rect 121920 85274 121972 85280
rect 122760 79898 122788 91151
rect 122852 86630 122880 91423
rect 124048 90778 124076 92375
rect 125414 91352 125470 91361
rect 125414 91287 125470 91296
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 124036 90772 124088 90778
rect 124036 90714 124088 90720
rect 122840 86624 122892 86630
rect 122840 86566 122892 86572
rect 122748 79892 122800 79898
rect 122748 79834 122800 79840
rect 124140 78538 124168 91151
rect 125428 83842 125456 91287
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 126886 91216 126942 91225
rect 126886 91151 126942 91160
rect 125416 83836 125468 83842
rect 125416 83778 125468 83784
rect 125520 82686 125548 91151
rect 125508 82680 125560 82686
rect 125508 82622 125560 82628
rect 126900 81326 126928 91151
rect 129476 90914 129504 92375
rect 133156 92206 133184 92375
rect 133144 92200 133196 92206
rect 133144 92142 133196 92148
rect 135732 92138 135760 92375
rect 135720 92132 135772 92138
rect 135720 92074 135772 92080
rect 132222 91624 132278 91633
rect 132222 91559 132278 91568
rect 151358 91624 151414 91633
rect 151358 91559 151414 91568
rect 129464 90908 129516 90914
rect 129464 90850 129516 90856
rect 132236 89350 132264 91559
rect 134798 91216 134854 91225
rect 134798 91151 134854 91160
rect 134524 91112 134576 91118
rect 134524 91054 134576 91060
rect 132224 89344 132276 89350
rect 132224 89286 132276 89292
rect 126888 81320 126940 81326
rect 126888 81262 126940 81268
rect 124128 78532 124180 78538
rect 124128 78474 124180 78480
rect 134536 78470 134564 91054
rect 134812 88126 134840 91151
rect 151372 89418 151400 91559
rect 151556 90710 151584 92375
rect 152108 92274 152136 92375
rect 152096 92268 152148 92274
rect 152096 92210 152148 92216
rect 151544 90704 151596 90710
rect 151544 90646 151596 90652
rect 151360 89412 151412 89418
rect 151360 89354 151412 89360
rect 164896 88262 164924 97990
rect 166276 89350 166304 144910
rect 170404 133952 170456 133958
rect 170404 133894 170456 133900
rect 167644 124228 167696 124234
rect 167644 124170 167696 124176
rect 166356 122868 166408 122874
rect 166356 122810 166408 122816
rect 166264 89344 166316 89350
rect 166264 89286 166316 89292
rect 164884 88256 164936 88262
rect 164884 88198 164936 88204
rect 134800 88120 134852 88126
rect 134800 88062 134852 88068
rect 166368 87990 166396 122810
rect 166448 107704 166500 107710
rect 166448 107646 166500 107652
rect 166356 87984 166408 87990
rect 166356 87926 166408 87932
rect 166460 83978 166488 107646
rect 166540 101448 166592 101454
rect 166540 101390 166592 101396
rect 166552 92138 166580 101390
rect 166540 92132 166592 92138
rect 166540 92074 166592 92080
rect 167656 86630 167684 124170
rect 169024 121508 169076 121514
rect 169024 121450 169076 121456
rect 167736 118720 167788 118726
rect 167736 118662 167788 118668
rect 167644 86624 167696 86630
rect 167644 86566 167696 86572
rect 167748 85270 167776 118662
rect 168288 111784 168340 111790
rect 168286 111752 168288 111761
rect 168340 111752 168342 111761
rect 168286 111687 168342 111696
rect 167828 110424 167880 110430
rect 167828 110366 167880 110372
rect 167840 110129 167868 110366
rect 167826 110120 167882 110129
rect 167826 110055 167882 110064
rect 168104 108996 168156 109002
rect 168104 108938 168156 108944
rect 168116 108769 168144 108938
rect 168102 108760 168158 108769
rect 168102 108695 168158 108704
rect 167920 102808 167972 102814
rect 167920 102750 167972 102756
rect 167828 99408 167880 99414
rect 167828 99350 167880 99356
rect 167736 85264 167788 85270
rect 167736 85206 167788 85212
rect 166448 83972 166500 83978
rect 166448 83914 166500 83920
rect 167840 79830 167868 99350
rect 167932 92206 167960 102750
rect 167920 92200 167972 92206
rect 167920 92142 167972 92148
rect 169036 88058 169064 121450
rect 169300 120148 169352 120154
rect 169300 120090 169352 120096
rect 169208 117360 169260 117366
rect 169208 117302 169260 117308
rect 169116 111852 169168 111858
rect 169116 111794 169168 111800
rect 169024 88052 169076 88058
rect 169024 87994 169076 88000
rect 169128 81190 169156 111794
rect 169220 90846 169248 117302
rect 169312 94110 169340 120090
rect 169300 94104 169352 94110
rect 169300 94046 169352 94052
rect 169208 90840 169260 90846
rect 169208 90782 169260 90788
rect 170416 88233 170444 133894
rect 170496 127016 170548 127022
rect 170496 126958 170548 126964
rect 170402 88224 170458 88233
rect 170402 88159 170458 88168
rect 170508 82550 170536 126958
rect 170588 109064 170640 109070
rect 170588 109006 170640 109012
rect 170600 84046 170628 109006
rect 170680 107772 170732 107778
rect 170680 107714 170732 107720
rect 170692 93906 170720 107714
rect 170680 93900 170732 93906
rect 170680 93842 170732 93848
rect 171796 93430 171824 144978
rect 171876 136672 171928 136678
rect 171876 136614 171928 136620
rect 171784 93424 171836 93430
rect 171784 93366 171836 93372
rect 171888 92342 171916 136614
rect 173164 132524 173216 132530
rect 173164 132466 173216 132472
rect 171968 124296 172020 124302
rect 171968 124238 172020 124244
rect 171876 92336 171928 92342
rect 171876 92278 171928 92284
rect 171980 90778 172008 124238
rect 172060 98116 172112 98122
rect 172060 98058 172112 98064
rect 171968 90772 172020 90778
rect 171968 90714 172020 90720
rect 170588 84040 170640 84046
rect 170588 83982 170640 83988
rect 170496 82544 170548 82550
rect 170496 82486 170548 82492
rect 169116 81184 169168 81190
rect 169116 81126 169168 81132
rect 167828 79824 167880 79830
rect 167828 79766 167880 79772
rect 172072 78606 172100 98058
rect 173176 81122 173204 132466
rect 173348 118788 173400 118794
rect 173348 118730 173400 118736
rect 173256 113212 173308 113218
rect 173256 113154 173308 113160
rect 173268 86698 173296 113154
rect 173360 93294 173388 118730
rect 173440 110492 173492 110498
rect 173440 110434 173492 110440
rect 173348 93288 173400 93294
rect 173348 93230 173400 93236
rect 173452 89554 173480 110434
rect 174556 96626 174584 265610
rect 175004 242344 175056 242350
rect 175004 242286 175056 242292
rect 175016 241534 175044 242286
rect 175004 241528 175056 241534
rect 175004 241470 175056 241476
rect 175016 237153 175044 241470
rect 175002 237144 175058 237153
rect 175002 237079 175058 237088
rect 175108 224262 175136 338098
rect 175200 334626 175228 362199
rect 175924 357808 175976 357814
rect 175924 357750 175976 357756
rect 175936 340202 175964 357750
rect 175924 340196 175976 340202
rect 175924 340138 175976 340144
rect 175188 334620 175240 334626
rect 175188 334562 175240 334568
rect 175200 331906 175228 334562
rect 175188 331900 175240 331906
rect 175188 331842 175240 331848
rect 175188 321632 175240 321638
rect 175188 321574 175240 321580
rect 175096 224256 175148 224262
rect 175096 224198 175148 224204
rect 174636 134020 174688 134026
rect 174636 133962 174688 133968
rect 174544 96620 174596 96626
rect 174544 96562 174596 96568
rect 173440 89548 173492 89554
rect 173440 89490 173492 89496
rect 173256 86692 173308 86698
rect 173256 86634 173308 86640
rect 174648 85406 174676 133962
rect 174728 109132 174780 109138
rect 174728 109074 174780 109080
rect 174740 93226 174768 109074
rect 174728 93220 174780 93226
rect 174728 93162 174780 93168
rect 174636 85400 174688 85406
rect 174636 85342 174688 85348
rect 173164 81116 173216 81122
rect 173164 81058 173216 81064
rect 172060 78600 172112 78606
rect 172060 78542 172112 78548
rect 134524 78464 134576 78470
rect 134524 78406 134576 78412
rect 119344 75812 119396 75818
rect 119344 75754 119396 75760
rect 139400 75268 139452 75274
rect 139400 75210 139452 75216
rect 104808 73160 104860 73166
rect 104808 73102 104860 73108
rect 124220 72548 124272 72554
rect 124220 72490 124272 72496
rect 88340 71120 88392 71126
rect 88340 71062 88392 71068
rect 80060 65544 80112 65550
rect 80060 65486 80112 65492
rect 77300 49088 77352 49094
rect 77300 49030 77352 49036
rect 77312 16574 77340 49030
rect 78680 26920 78732 26926
rect 78680 26862 78732 26868
rect 78692 16574 78720 26862
rect 80072 16574 80100 65486
rect 85580 58676 85632 58682
rect 85580 58618 85632 58624
rect 81440 43512 81492 43518
rect 81440 43454 81492 43460
rect 81452 16574 81480 43454
rect 82820 25628 82872 25634
rect 82820 25570 82872 25576
rect 82832 16574 82860 25570
rect 77312 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77392 4956 77444 4962
rect 77392 4898 77444 4904
rect 77404 480 77432 4898
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 84200 14476 84252 14482
rect 84200 14418 84252 14424
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 14418
rect 85592 3602 85620 58618
rect 85672 40792 85724 40798
rect 85672 40734 85724 40740
rect 85580 3596 85632 3602
rect 85580 3538 85632 3544
rect 85684 480 85712 40734
rect 86960 28348 87012 28354
rect 86960 28290 87012 28296
rect 86972 16574 87000 28290
rect 88352 16574 88380 71062
rect 89720 68332 89772 68338
rect 89720 68274 89772 68280
rect 89732 16574 89760 68274
rect 100760 66972 100812 66978
rect 100760 66914 100812 66920
rect 95240 61464 95292 61470
rect 95240 61406 95292 61412
rect 92480 47660 92532 47666
rect 92480 47602 92532 47608
rect 91100 32428 91152 32434
rect 91100 32370 91152 32376
rect 91112 16574 91140 32370
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 86500 3596 86552 3602
rect 86500 3538 86552 3544
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3538
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 47602
rect 93860 28280 93912 28286
rect 93860 28222 93912 28228
rect 93872 6914 93900 28222
rect 93952 18624 94004 18630
rect 93952 18566 94004 18572
rect 93964 16574 93992 18566
rect 95252 16574 95280 61406
rect 99380 60104 99432 60110
rect 99380 60046 99432 60052
rect 98000 29640 98052 29646
rect 98000 29582 98052 29588
rect 96620 17332 96672 17338
rect 96620 17274 96672 17280
rect 96632 16574 96660 17274
rect 98012 16574 98040 29582
rect 99392 16574 99420 60046
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 66914
rect 110420 65612 110472 65618
rect 110420 65554 110472 65560
rect 106280 58744 106332 58750
rect 106280 58686 106332 58692
rect 103520 57316 103572 57322
rect 103520 57258 103572 57264
rect 102140 20052 102192 20058
rect 102140 19994 102192 20000
rect 102152 16574 102180 19994
rect 103532 16574 103560 57258
rect 104900 17264 104952 17270
rect 104900 17206 104952 17212
rect 104912 16574 104940 17206
rect 106292 16574 106320 58686
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 102244 480 102272 16546
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103348 480 103376 3538
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108120 14544 108172 14550
rect 108120 14486 108172 14492
rect 108132 480 108160 14486
rect 109040 13116 109092 13122
rect 109040 13058 109092 13064
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 13058
rect 110432 3398 110460 65554
rect 110512 55956 110564 55962
rect 110512 55898 110564 55904
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 55898
rect 118700 42152 118752 42158
rect 118700 42094 118752 42100
rect 117320 26988 117372 26994
rect 117320 26930 117372 26936
rect 113180 24132 113232 24138
rect 113180 24074 113232 24080
rect 111800 21412 111852 21418
rect 111800 21354 111852 21360
rect 111812 16574 111840 21354
rect 113192 16574 113220 24074
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 115204 7676 115256 7682
rect 115204 7618 115256 7624
rect 115216 480 115244 7618
rect 116400 6248 116452 6254
rect 116400 6190 116452 6196
rect 116412 480 116440 6190
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 26930
rect 118712 16574 118740 42094
rect 121460 39500 121512 39506
rect 121460 39442 121512 39448
rect 121472 16574 121500 39442
rect 124232 16574 124260 72490
rect 128360 38004 128412 38010
rect 128360 37946 128412 37952
rect 128372 16574 128400 37946
rect 139412 16574 139440 75210
rect 143540 33924 143592 33930
rect 143540 33866 143592 33872
rect 118712 16546 118832 16574
rect 121472 16546 122328 16574
rect 124232 16546 124720 16574
rect 128372 16546 128952 16574
rect 139412 16546 139624 16574
rect 118804 480 118832 16546
rect 120632 10328 120684 10334
rect 120632 10270 120684 10276
rect 119896 9036 119948 9042
rect 119896 8978 119948 8984
rect 119908 480 119936 8978
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 10270
rect 122300 480 122328 16546
rect 123484 9104 123536 9110
rect 123484 9046 123536 9052
rect 123496 480 123524 9046
rect 124692 480 124720 16546
rect 125874 3360 125930 3369
rect 125874 3295 125930 3304
rect 125888 480 125916 3295
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 135258 13016 135314 13025
rect 135258 12951 135314 12960
rect 132960 3664 133012 3670
rect 132960 3606 133012 3612
rect 132972 480 133000 3606
rect 135272 3398 135300 12951
rect 135260 3392 135312 3398
rect 135260 3334 135312 3340
rect 136456 3392 136508 3398
rect 136456 3334 136508 3340
rect 136468 480 136496 3334
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 143552 480 143580 33866
rect 175200 6322 175228 321574
rect 176304 271862 176332 371855
rect 176292 271856 176344 271862
rect 176292 271798 176344 271804
rect 176396 263945 176424 373215
rect 176580 336705 176608 381550
rect 177948 380248 178000 380254
rect 177948 380190 178000 380196
rect 177764 370592 177816 370598
rect 177764 370534 177816 370540
rect 176658 348120 176714 348129
rect 176658 348055 176714 348064
rect 176672 347818 176700 348055
rect 176660 347812 176712 347818
rect 176660 347754 176712 347760
rect 176660 345704 176712 345710
rect 176660 345646 176712 345652
rect 176672 345545 176700 345646
rect 176658 345536 176714 345545
rect 176658 345471 176714 345480
rect 177670 342272 177726 342281
rect 177670 342207 177726 342216
rect 176658 341320 176714 341329
rect 176658 341255 176714 341264
rect 176672 340882 176700 341255
rect 176660 340876 176712 340882
rect 176660 340818 176712 340824
rect 176658 339280 176714 339289
rect 176658 339215 176714 339224
rect 176672 338162 176700 339215
rect 176660 338156 176712 338162
rect 176660 338098 176712 338104
rect 176566 336696 176622 336705
rect 176566 336631 176622 336640
rect 176658 334656 176714 334665
rect 176658 334591 176660 334600
rect 176712 334591 176714 334600
rect 176660 334562 176712 334568
rect 176660 333940 176712 333946
rect 176660 333882 176712 333888
rect 176672 332625 176700 333882
rect 176658 332616 176714 332625
rect 176658 332551 176714 332560
rect 176566 327720 176622 327729
rect 176566 327655 176622 327664
rect 176474 301200 176530 301209
rect 176474 301135 176530 301144
rect 176382 263936 176438 263945
rect 176382 263871 176438 263880
rect 176382 250880 176438 250889
rect 176382 250815 176438 250824
rect 175924 249076 175976 249082
rect 175924 249018 175976 249024
rect 175936 95169 175964 249018
rect 176396 240281 176424 250815
rect 176382 240272 176438 240281
rect 176382 240207 176438 240216
rect 175922 95160 175978 95169
rect 175922 95095 175978 95104
rect 176488 19310 176516 301135
rect 176580 23458 176608 327655
rect 176658 325816 176714 325825
rect 176658 325751 176714 325760
rect 176672 325718 176700 325751
rect 176660 325712 176712 325718
rect 176660 325654 176712 325660
rect 177580 321632 177632 321638
rect 177578 321600 177580 321609
rect 177632 321600 177634 321609
rect 177578 321535 177634 321544
rect 176658 312760 176714 312769
rect 176658 312695 176714 312704
rect 176672 312594 176700 312695
rect 176660 312588 176712 312594
rect 176660 312530 176712 312536
rect 176660 310276 176712 310282
rect 176660 310218 176712 310224
rect 176672 310185 176700 310218
rect 176658 310176 176714 310185
rect 176658 310111 176714 310120
rect 176660 306128 176712 306134
rect 176658 306096 176660 306105
rect 176712 306096 176714 306105
rect 176658 306031 176714 306040
rect 176660 299464 176712 299470
rect 176660 299406 176712 299412
rect 176672 299305 176700 299406
rect 176658 299296 176714 299305
rect 176658 299231 176714 299240
rect 176658 297120 176714 297129
rect 176658 297055 176714 297064
rect 176672 296954 176700 297055
rect 176660 296948 176712 296954
rect 176660 296890 176712 296896
rect 176658 295080 176714 295089
rect 176658 295015 176714 295024
rect 176672 294030 176700 295015
rect 176660 294024 176712 294030
rect 176660 293966 176712 293972
rect 176660 290488 176712 290494
rect 176658 290456 176660 290465
rect 176712 290456 176714 290465
rect 176658 290391 176714 290400
rect 176660 288312 176712 288318
rect 176658 288280 176660 288289
rect 176712 288280 176714 288289
rect 176658 288215 176714 288224
rect 177302 286240 177358 286249
rect 177302 286175 177358 286184
rect 176660 284300 176712 284306
rect 176660 284242 176712 284248
rect 176672 283665 176700 284242
rect 176658 283656 176714 283665
rect 176658 283591 176714 283600
rect 176660 282872 176712 282878
rect 176660 282814 176712 282820
rect 176672 281625 176700 282814
rect 176658 281616 176714 281625
rect 176658 281551 176714 281560
rect 176660 280152 176712 280158
rect 176660 280094 176712 280100
rect 176672 279585 176700 280094
rect 176658 279576 176714 279585
rect 176658 279511 176714 279520
rect 176658 277536 176714 277545
rect 176658 277471 176714 277480
rect 176672 277438 176700 277471
rect 176660 277432 176712 277438
rect 176660 277374 176712 277380
rect 176658 274816 176714 274825
rect 176658 274751 176660 274760
rect 176712 274751 176714 274760
rect 176660 274722 176712 274728
rect 176658 272640 176714 272649
rect 176658 272575 176714 272584
rect 176672 271930 176700 272575
rect 176660 271924 176712 271930
rect 176660 271866 176712 271872
rect 177316 269822 177344 286175
rect 177304 269816 177356 269822
rect 177304 269758 177356 269764
rect 176658 268560 176714 268569
rect 176658 268495 176714 268504
rect 176672 267782 176700 268495
rect 176660 267776 176712 267782
rect 176660 267718 176712 267724
rect 176660 266348 176712 266354
rect 176660 266290 176712 266296
rect 176672 265985 176700 266290
rect 176658 265976 176714 265985
rect 176658 265911 176714 265920
rect 176658 261760 176714 261769
rect 176658 261695 176714 261704
rect 176672 261526 176700 261695
rect 176660 261520 176712 261526
rect 176660 261462 176712 261468
rect 176658 257000 176714 257009
rect 176658 256935 176714 256944
rect 176672 256766 176700 256935
rect 176660 256760 176712 256766
rect 176660 256702 176712 256708
rect 176660 255264 176712 255270
rect 176660 255206 176712 255212
rect 176672 255105 176700 255206
rect 176658 255096 176714 255105
rect 176658 255031 176714 255040
rect 176658 246120 176714 246129
rect 176658 246055 176714 246064
rect 176672 245682 176700 246055
rect 176660 245676 176712 245682
rect 176660 245618 176712 245624
rect 176658 242040 176714 242049
rect 176658 241975 176714 241984
rect 176672 241534 176700 241975
rect 176660 241528 176712 241534
rect 176660 241470 176712 241476
rect 177684 193934 177712 342207
rect 177776 321638 177804 370534
rect 177856 359644 177908 359650
rect 177856 359586 177908 359592
rect 177868 343505 177896 359586
rect 177854 343496 177910 343505
rect 177854 343431 177910 343440
rect 177868 342281 177896 343431
rect 177854 342272 177910 342281
rect 177854 342207 177910 342216
rect 177854 330440 177910 330449
rect 177854 330375 177910 330384
rect 177764 321632 177816 321638
rect 177764 321574 177816 321580
rect 177762 259720 177818 259729
rect 177762 259655 177818 259664
rect 177672 193928 177724 193934
rect 177672 193870 177724 193876
rect 177776 73982 177804 259655
rect 177764 73976 177816 73982
rect 177764 73918 177816 73924
rect 177868 42226 177896 330375
rect 177960 317422 177988 380190
rect 179236 365152 179288 365158
rect 179236 365094 179288 365100
rect 179142 355328 179198 355337
rect 179142 355263 179198 355272
rect 178682 354920 178738 354929
rect 178682 354855 178738 354864
rect 178696 345030 178724 354855
rect 178684 345024 178736 345030
rect 178684 344966 178736 344972
rect 179156 319025 179184 355263
rect 179248 354385 179276 365094
rect 179234 354376 179290 354385
rect 179234 354311 179290 354320
rect 179248 347070 179276 354311
rect 179236 347064 179288 347070
rect 179236 347006 179288 347012
rect 179142 319016 179198 319025
rect 179142 318951 179198 318960
rect 177948 317416 178000 317422
rect 177948 317358 178000 317364
rect 179144 317416 179196 317422
rect 179144 317358 179196 317364
rect 179156 316849 179184 317358
rect 179142 316840 179198 316849
rect 179142 316775 179198 316784
rect 177946 303920 178002 303929
rect 177946 303855 178002 303864
rect 177856 42220 177908 42226
rect 177856 42162 177908 42168
rect 176568 23452 176620 23458
rect 176568 23394 176620 23400
rect 176476 19304 176528 19310
rect 176476 19246 176528 19252
rect 177960 13190 177988 303855
rect 178684 292596 178736 292602
rect 178684 292538 178736 292544
rect 178696 238746 178724 292538
rect 178684 238740 178736 238746
rect 178684 238682 178736 238688
rect 179156 204950 179184 316775
rect 179340 314854 179368 393994
rect 181456 387190 181484 402902
rect 182180 387864 182232 387870
rect 182180 387806 182232 387812
rect 181444 387184 181496 387190
rect 181444 387126 181496 387132
rect 179880 384464 179932 384470
rect 179880 384406 179932 384412
rect 179420 354884 179472 354890
rect 179420 354826 179472 354832
rect 179432 354006 179460 354826
rect 179420 354000 179472 354006
rect 179420 353942 179472 353948
rect 179892 350033 179920 384406
rect 180798 368520 180854 368529
rect 180798 368455 180854 368464
rect 180812 364334 180840 368455
rect 182192 364334 182220 387806
rect 183572 383110 183600 405062
rect 187712 402354 187740 405076
rect 187700 402348 187752 402354
rect 187700 402290 187752 402296
rect 190932 402286 190960 405076
rect 194152 403646 194180 405076
rect 194140 403640 194192 403646
rect 194140 403582 194192 403588
rect 190920 402280 190972 402286
rect 190920 402222 190972 402228
rect 191748 402280 191800 402286
rect 191748 402222 191800 402228
rect 189724 394120 189776 394126
rect 189724 394062 189776 394068
rect 183560 383104 183612 383110
rect 183560 383046 183612 383052
rect 186964 376032 187016 376038
rect 186964 375974 187016 375980
rect 180812 364306 180932 364334
rect 182192 364306 182864 364334
rect 180904 355042 180932 364306
rect 182836 355042 182864 364306
rect 184938 357504 184994 357513
rect 184938 357439 184994 357448
rect 184952 355042 184980 357439
rect 186780 356244 186832 356250
rect 186780 356186 186832 356192
rect 186792 355042 186820 356186
rect 186976 355337 187004 375974
rect 189080 365900 189132 365906
rect 189080 365842 189132 365848
rect 189092 364334 189120 365842
rect 189092 364306 189304 364334
rect 186962 355328 187018 355337
rect 186962 355263 187018 355272
rect 189276 355042 189304 364306
rect 189736 355434 189764 394062
rect 191760 378894 191788 402222
rect 195244 396772 195296 396778
rect 195244 396714 195296 396720
rect 191104 378888 191156 378894
rect 191104 378830 191156 378836
rect 191748 378888 191800 378894
rect 191748 378830 191800 378836
rect 191116 355502 191144 378830
rect 191746 360224 191802 360233
rect 191746 360159 191802 360168
rect 191104 355496 191156 355502
rect 191104 355438 191156 355444
rect 189724 355428 189776 355434
rect 189724 355370 189776 355376
rect 191760 355042 191788 360159
rect 193404 358964 193456 358970
rect 193404 358906 193456 358912
rect 193416 356250 193444 358906
rect 195256 357814 195284 396714
rect 197372 395350 197400 405076
rect 200592 404258 200620 405076
rect 202892 405062 203826 405090
rect 201408 404456 201460 404462
rect 201408 404398 201460 404404
rect 201420 404258 201448 404398
rect 200580 404252 200632 404258
rect 200580 404194 200632 404200
rect 201408 404252 201460 404258
rect 201408 404194 201460 404200
rect 200592 402974 200620 404194
rect 200592 402946 200804 402974
rect 197360 395344 197412 395350
rect 197360 395286 197412 395292
rect 197360 391332 197412 391338
rect 197360 391274 197412 391280
rect 197372 364334 197400 391274
rect 200776 377670 200804 402946
rect 202144 385688 202196 385694
rect 202144 385630 202196 385636
rect 200764 377664 200816 377670
rect 200764 377606 200816 377612
rect 197372 364306 197676 364334
rect 195244 357808 195296 357814
rect 195244 357750 195296 357756
rect 193404 356244 193456 356250
rect 193404 356186 193456 356192
rect 180904 355014 181332 355042
rect 182836 355014 183264 355042
rect 184952 355014 185196 355042
rect 186792 355014 187128 355042
rect 189276 355014 189704 355042
rect 191636 355014 191788 355042
rect 193416 354906 193444 356186
rect 195256 355042 195284 357750
rect 197648 355042 197676 364306
rect 202156 361690 202184 385630
rect 201592 361684 201644 361690
rect 201592 361626 201644 361632
rect 202144 361684 202196 361690
rect 202144 361626 202196 361632
rect 199660 356312 199712 356318
rect 199660 356254 199712 356260
rect 199672 355042 199700 356254
rect 201604 355042 201632 361626
rect 202892 357542 202920 405062
rect 206388 396846 206416 405076
rect 208412 405062 209622 405090
rect 212552 405062 212842 405090
rect 215312 405062 216062 405090
rect 219282 405062 219388 405090
rect 206376 396840 206428 396846
rect 206376 396782 206428 396788
rect 205640 391400 205692 391406
rect 205640 391342 205692 391348
rect 202972 387932 203024 387938
rect 202972 387874 203024 387880
rect 202984 364334 203012 387874
rect 205652 364334 205680 391342
rect 208412 367878 208440 405062
rect 209780 379568 209832 379574
rect 209780 379510 209832 379516
rect 208492 370728 208544 370734
rect 208492 370670 208544 370676
rect 208400 367872 208452 367878
rect 208400 367814 208452 367820
rect 208504 367198 208532 370670
rect 208492 367192 208544 367198
rect 208492 367134 208544 367140
rect 202984 364306 203472 364334
rect 205652 364306 206048 364334
rect 202880 357536 202932 357542
rect 202880 357478 202932 357484
rect 203444 355042 203472 364306
rect 206020 355042 206048 364306
rect 208504 355042 208532 367134
rect 209792 364334 209820 379510
rect 209792 364306 209912 364334
rect 195256 355014 195500 355042
rect 197648 355014 198076 355042
rect 199672 355014 200160 355042
rect 201604 355014 201940 355042
rect 203444 355014 203872 355042
rect 206020 355014 206448 355042
rect 208380 355014 208532 355042
rect 209884 355042 209912 364306
rect 212552 363050 212580 405062
rect 214564 395344 214616 395350
rect 214564 395286 214616 395292
rect 212540 363044 212592 363050
rect 212540 362986 212592 362992
rect 212552 362370 212580 362986
rect 212540 362364 212592 362370
rect 212540 362306 212592 362312
rect 214576 357814 214604 395286
rect 215312 375358 215340 405062
rect 219360 402966 219388 405062
rect 219348 402960 219400 402966
rect 219348 402902 219400 402908
rect 219360 387938 219388 402902
rect 222488 402898 222516 405076
rect 222476 402892 222528 402898
rect 222476 402834 222528 402840
rect 225708 402257 225736 405076
rect 227732 405062 228942 405090
rect 225694 402248 225750 402257
rect 225694 402183 225750 402192
rect 227628 396840 227680 396846
rect 227628 396782 227680 396788
rect 218704 387932 218756 387938
rect 218704 387874 218756 387880
rect 219348 387932 219400 387938
rect 219348 387874 219400 387880
rect 218716 380186 218744 387874
rect 219440 381676 219492 381682
rect 219440 381618 219492 381624
rect 218704 380180 218756 380186
rect 218704 380122 218756 380128
rect 215300 375352 215352 375358
rect 215300 375294 215352 375300
rect 218060 367260 218112 367266
rect 218060 367202 218112 367208
rect 216680 366376 216732 366382
rect 216680 366318 216732 366324
rect 212356 357808 212408 357814
rect 212356 357750 212408 357756
rect 214564 357808 214616 357814
rect 214564 357750 214616 357756
rect 212368 356794 212396 357750
rect 212448 357604 212500 357610
rect 212448 357546 212500 357552
rect 212460 357406 212488 357546
rect 212448 357400 212500 357406
rect 212448 357342 212500 357348
rect 212356 356788 212408 356794
rect 212356 356730 212408 356736
rect 212460 355042 212488 357342
rect 209884 355014 210312 355042
rect 212244 355014 212488 355042
rect 214576 355042 214604 357750
rect 216692 355314 216720 366318
rect 218072 364334 218100 367202
rect 218072 364306 218284 364334
rect 216692 355286 216766 355314
rect 214576 355014 214820 355042
rect 216738 355028 216766 355286
rect 218256 355042 218284 364306
rect 218256 355014 218684 355042
rect 193416 354878 193568 354906
rect 200132 354793 200160 355014
rect 200118 354784 200174 354793
rect 209884 354754 209912 355014
rect 219452 354890 219480 381618
rect 222200 379636 222252 379642
rect 222200 379578 222252 379584
rect 222212 364334 222240 379578
rect 224960 369232 225012 369238
rect 224960 369174 225012 369180
rect 222212 364306 222792 364334
rect 222764 355042 222792 364306
rect 224972 355042 225000 369174
rect 227640 361690 227668 396782
rect 227732 386374 227760 405062
rect 232148 403714 232176 405076
rect 234632 405062 235382 405090
rect 238602 405062 238708 405090
rect 232504 403844 232556 403850
rect 232504 403786 232556 403792
rect 232136 403708 232188 403714
rect 232136 403650 232188 403656
rect 227720 386368 227772 386374
rect 227720 386310 227772 386316
rect 228364 386368 228416 386374
rect 228364 386310 228416 386316
rect 228376 366353 228404 386310
rect 231124 383104 231176 383110
rect 231124 383046 231176 383052
rect 228362 366344 228418 366353
rect 228362 366279 228418 366288
rect 228824 363724 228876 363730
rect 228824 363666 228876 363672
rect 227352 361684 227404 361690
rect 227352 361626 227404 361632
rect 227628 361684 227680 361690
rect 227628 361626 227680 361632
rect 227364 355042 227392 361626
rect 222764 355014 223192 355042
rect 224972 355014 225124 355042
rect 227056 355014 227392 355042
rect 220464 354890 220616 354906
rect 219440 354884 219492 354890
rect 219440 354826 219492 354832
rect 220452 354884 220616 354890
rect 220504 354878 220616 354884
rect 220452 354826 220504 354832
rect 228836 354770 228864 363666
rect 231136 357610 231164 383046
rect 232516 370530 232544 403786
rect 234632 383110 234660 405062
rect 238680 402830 238708 405062
rect 241808 404326 241836 405076
rect 241796 404320 241848 404326
rect 241796 404262 241848 404268
rect 241808 404122 241836 404262
rect 241796 404116 241848 404122
rect 241796 404058 241848 404064
rect 242808 404116 242860 404122
rect 242808 404058 242860 404064
rect 238668 402824 238720 402830
rect 238668 402766 238720 402772
rect 238680 389201 238708 402766
rect 242820 398954 242848 404058
rect 242808 398948 242860 398954
rect 242808 398890 242860 398896
rect 238760 392080 238812 392086
rect 238760 392022 238812 392028
rect 238022 389192 238078 389201
rect 238022 389127 238078 389136
rect 238666 389192 238722 389201
rect 238666 389127 238722 389136
rect 234712 385076 234764 385082
rect 234712 385018 234764 385024
rect 234620 383104 234672 383110
rect 234620 383046 234672 383052
rect 234724 377534 234752 385018
rect 238036 377602 238064 389127
rect 238024 377596 238076 377602
rect 238024 377538 238076 377544
rect 234712 377528 234764 377534
rect 234712 377470 234764 377476
rect 234724 373994 234752 377470
rect 237380 376168 237432 376174
rect 237380 376110 237432 376116
rect 234632 373966 234752 373994
rect 232504 370524 232556 370530
rect 232504 370466 232556 370472
rect 234632 364334 234660 373966
rect 237392 371890 237420 376110
rect 237380 371884 237432 371890
rect 237380 371826 237432 371832
rect 234632 364306 235028 364334
rect 233790 358864 233846 358873
rect 233790 358799 233846 358808
rect 231124 357604 231176 357610
rect 231124 357546 231176 357552
rect 231136 355042 231164 357546
rect 233804 355042 233832 358799
rect 231136 355014 231564 355042
rect 233496 355014 233832 355042
rect 235000 355042 235028 364306
rect 237392 355314 237420 371826
rect 238772 364334 238800 392022
rect 241520 387184 241572 387190
rect 241520 387126 241572 387132
rect 238772 364306 239536 364334
rect 237346 355286 237420 355314
rect 235000 355014 235428 355042
rect 237346 355028 237374 355286
rect 239508 355042 239536 364306
rect 241532 355042 241560 387126
rect 242820 370666 242848 398890
rect 242912 392630 242940 567166
rect 242992 532772 243044 532778
rect 242992 532714 243044 532720
rect 242900 392624 242952 392630
rect 242900 392566 242952 392572
rect 242808 370660 242860 370666
rect 242808 370602 242860 370608
rect 243004 362234 243032 532714
rect 243096 373998 243124 586570
rect 244188 580984 244240 580990
rect 244188 580926 244240 580932
rect 243544 580576 243596 580582
rect 243544 580518 243596 580524
rect 243556 568546 243584 580518
rect 244200 579873 244228 580926
rect 244186 579864 244242 579873
rect 244186 579799 244242 579808
rect 244200 579698 244228 579799
rect 244188 579692 244240 579698
rect 244188 579634 244240 579640
rect 243544 568540 243596 568546
rect 243544 568482 243596 568488
rect 244936 562358 244964 586774
rect 245108 586764 245160 586770
rect 245108 586706 245160 586712
rect 245014 586664 245070 586673
rect 245014 586599 245070 586608
rect 244924 562352 244976 562358
rect 244924 562294 244976 562300
rect 244924 561672 244976 561678
rect 244924 561614 244976 561620
rect 244278 543144 244334 543153
rect 244278 543079 244334 543088
rect 244188 534064 244240 534070
rect 244188 534006 244240 534012
rect 244200 532953 244228 534006
rect 244186 532944 244242 532953
rect 244186 532879 244242 532888
rect 244200 532778 244228 532879
rect 244188 532772 244240 532778
rect 244188 532714 244240 532720
rect 244186 398712 244242 398721
rect 244186 398647 244242 398656
rect 243084 373992 243136 373998
rect 243084 373934 243136 373940
rect 243096 373386 243124 373934
rect 243084 373380 243136 373386
rect 243084 373322 243136 373328
rect 244200 367810 244228 398647
rect 244292 384402 244320 543079
rect 244370 418704 244426 418713
rect 244370 418639 244426 418648
rect 244384 395350 244412 418639
rect 244372 395344 244424 395350
rect 244372 395286 244424 395292
rect 244280 384396 244332 384402
rect 244280 384338 244332 384344
rect 244936 381682 244964 561614
rect 245028 558249 245056 586599
rect 245120 578950 245148 586706
rect 245108 578944 245160 578950
rect 245108 578886 245160 578892
rect 245672 576570 245700 702714
rect 251088 702568 251140 702574
rect 267660 702545 267688 703520
rect 251088 702510 251140 702516
rect 267646 702536 267702 702545
rect 247040 700324 247092 700330
rect 247040 700266 247092 700272
rect 245844 614780 245896 614786
rect 245844 614722 245896 614728
rect 245750 583264 245806 583273
rect 245750 583199 245806 583208
rect 245764 582418 245792 583199
rect 245752 582412 245804 582418
rect 245752 582354 245804 582360
rect 245752 582276 245804 582282
rect 245752 582218 245804 582224
rect 245660 576564 245712 576570
rect 245660 576506 245712 576512
rect 245658 576464 245714 576473
rect 245658 576399 245714 576408
rect 245672 575550 245700 576399
rect 245660 575544 245712 575550
rect 245660 575486 245712 575492
rect 245658 573064 245714 573073
rect 245658 572999 245714 573008
rect 245672 572014 245700 572999
rect 245660 572008 245712 572014
rect 245660 571950 245712 571956
rect 245658 569664 245714 569673
rect 245658 569599 245714 569608
rect 245672 569226 245700 569599
rect 245660 569220 245712 569226
rect 245660 569162 245712 569168
rect 245566 562864 245622 562873
rect 245566 562799 245622 562808
rect 245580 561678 245608 562799
rect 245568 561672 245620 561678
rect 245568 561614 245620 561620
rect 245014 558240 245070 558249
rect 245014 558175 245070 558184
rect 245658 556744 245714 556753
rect 245658 556679 245714 556688
rect 245672 551342 245700 556679
rect 245660 551336 245712 551342
rect 245660 551278 245712 551284
rect 245292 543720 245344 543726
rect 245292 543662 245344 543668
rect 245304 543153 245332 543662
rect 245290 543144 245346 543153
rect 245290 543079 245346 543088
rect 245764 516066 245792 582218
rect 245856 536353 245884 614722
rect 245936 584588 245988 584594
rect 245936 584530 245988 584536
rect 245948 582282 245976 584530
rect 245936 582276 245988 582282
rect 245936 582218 245988 582224
rect 245936 576564 245988 576570
rect 245936 576506 245988 576512
rect 245948 569226 245976 576506
rect 245936 569220 245988 569226
rect 245936 569162 245988 569168
rect 245934 566264 245990 566273
rect 245934 566199 245990 566208
rect 245948 565894 245976 566199
rect 245936 565888 245988 565894
rect 245936 565830 245988 565836
rect 245934 560144 245990 560153
rect 245934 560079 245990 560088
rect 245948 558958 245976 560079
rect 245936 558952 245988 558958
rect 245936 558894 245988 558900
rect 245934 553344 245990 553353
rect 245934 553279 245990 553288
rect 245948 552090 245976 553279
rect 245936 552084 245988 552090
rect 245936 552026 245988 552032
rect 245934 549944 245990 549953
rect 245934 549879 245990 549888
rect 245948 549302 245976 549879
rect 245936 549296 245988 549302
rect 245936 549238 245988 549244
rect 245934 546544 245990 546553
rect 245934 546479 245936 546488
rect 245988 546479 245990 546488
rect 245936 546450 245988 546456
rect 246946 540288 247002 540297
rect 246946 540223 247002 540232
rect 245842 536344 245898 536353
rect 245842 536279 245898 536288
rect 245856 536110 245884 536279
rect 245844 536104 245896 536110
rect 245844 536046 245896 536052
rect 246854 529544 246910 529553
rect 246854 529479 246910 529488
rect 246868 528562 246896 529479
rect 246960 529242 246988 540223
rect 246948 529236 247000 529242
rect 246948 529178 247000 529184
rect 246856 528556 246908 528562
rect 246856 528498 246908 528504
rect 246868 527202 246896 528498
rect 246304 527196 246356 527202
rect 246304 527138 246356 527144
rect 246856 527196 246908 527202
rect 246856 527138 246908 527144
rect 245842 526144 245898 526153
rect 245842 526079 245898 526088
rect 245856 525065 245884 526079
rect 245842 525056 245898 525065
rect 245842 524991 245898 525000
rect 245842 522744 245898 522753
rect 245842 522679 245898 522688
rect 245856 521694 245884 522679
rect 245844 521688 245896 521694
rect 245844 521630 245896 521636
rect 245842 519344 245898 519353
rect 245842 519279 245898 519288
rect 245856 518974 245884 519279
rect 245844 518968 245896 518974
rect 245844 518910 245896 518916
rect 245764 516038 245976 516066
rect 245842 515944 245898 515953
rect 245842 515879 245898 515888
rect 245660 513324 245712 513330
rect 245660 513266 245712 513272
rect 245672 512553 245700 513266
rect 245658 512544 245714 512553
rect 245658 512479 245714 512488
rect 245856 512394 245884 515879
rect 245672 512366 245884 512394
rect 245014 492824 245070 492833
rect 245014 492759 245070 492768
rect 245028 389230 245056 492759
rect 245672 392018 245700 512366
rect 245844 509924 245896 509930
rect 245844 509866 245896 509872
rect 245856 509833 245884 509866
rect 245842 509824 245898 509833
rect 245842 509759 245898 509768
rect 245948 509234 245976 516038
rect 245764 509206 245976 509234
rect 245764 482633 245792 509206
rect 245842 506424 245898 506433
rect 245842 506359 245898 506368
rect 245856 505782 245884 506359
rect 245844 505776 245896 505782
rect 245844 505718 245896 505724
rect 245844 500540 245896 500546
rect 245844 500482 245896 500488
rect 245856 499633 245884 500482
rect 245842 499624 245898 499633
rect 245842 499559 245898 499568
rect 245842 496224 245898 496233
rect 245842 496159 245898 496168
rect 245856 495514 245884 496159
rect 245844 495508 245896 495514
rect 245844 495450 245896 495456
rect 245842 486024 245898 486033
rect 245842 485959 245898 485968
rect 245856 485858 245884 485959
rect 245844 485852 245896 485858
rect 245844 485794 245896 485800
rect 245750 482624 245806 482633
rect 245750 482559 245806 482568
rect 245764 482322 245792 482559
rect 245752 482316 245804 482322
rect 245752 482258 245804 482264
rect 245750 475824 245806 475833
rect 245750 475759 245806 475768
rect 245764 474774 245792 475759
rect 245752 474768 245804 474774
rect 245752 474710 245804 474716
rect 245842 472424 245898 472433
rect 245842 472359 245898 472368
rect 245856 472054 245884 472359
rect 245844 472048 245896 472054
rect 245844 471990 245896 471996
rect 245844 469192 245896 469198
rect 245844 469134 245896 469140
rect 245856 469033 245884 469134
rect 245842 469024 245898 469033
rect 245842 468959 245898 468968
rect 245842 465624 245898 465633
rect 245842 465559 245898 465568
rect 245856 465118 245884 465559
rect 245844 465112 245896 465118
rect 245844 465054 245896 465060
rect 245842 462224 245898 462233
rect 245842 462159 245898 462168
rect 245856 461650 245884 462159
rect 245844 461644 245896 461650
rect 245844 461586 245896 461592
rect 245842 459504 245898 459513
rect 245842 459439 245898 459448
rect 245856 458250 245884 459439
rect 245844 458244 245896 458250
rect 245844 458186 245896 458192
rect 245842 456104 245898 456113
rect 245842 456039 245898 456048
rect 245856 455462 245884 456039
rect 245844 455456 245896 455462
rect 245844 455398 245896 455404
rect 245844 454096 245896 454102
rect 245844 454038 245896 454044
rect 245856 452713 245884 454038
rect 245842 452704 245898 452713
rect 245842 452639 245898 452648
rect 245842 445904 245898 445913
rect 245842 445839 245898 445848
rect 245856 445806 245884 445839
rect 245844 445800 245896 445806
rect 245844 445742 245896 445748
rect 245842 439104 245898 439113
rect 245842 439039 245898 439048
rect 245856 438938 245884 439039
rect 245844 438932 245896 438938
rect 245844 438874 245896 438880
rect 245750 435704 245806 435713
rect 245750 435639 245806 435648
rect 245764 434790 245792 435639
rect 245752 434784 245804 434790
rect 245752 434726 245804 434732
rect 245844 432608 245896 432614
rect 245844 432550 245896 432556
rect 245856 432313 245884 432550
rect 245842 432304 245898 432313
rect 245842 432239 245898 432248
rect 245750 428904 245806 428913
rect 245750 428839 245806 428848
rect 245764 427854 245792 428839
rect 245752 427848 245804 427854
rect 245752 427790 245804 427796
rect 245842 425504 245898 425513
rect 245842 425439 245898 425448
rect 245856 425134 245884 425439
rect 245844 425128 245896 425134
rect 245844 425070 245896 425076
rect 245750 422104 245806 422113
rect 245750 422039 245806 422048
rect 245764 420986 245792 422039
rect 245752 420980 245804 420986
rect 245752 420922 245804 420928
rect 245844 415404 245896 415410
rect 245844 415346 245896 415352
rect 245856 415313 245884 415346
rect 245842 415304 245898 415313
rect 245842 415239 245898 415248
rect 245842 411904 245898 411913
rect 245842 411839 245898 411848
rect 245856 411330 245884 411839
rect 245844 411324 245896 411330
rect 245844 411266 245896 411272
rect 245842 409184 245898 409193
rect 245842 409119 245844 409128
rect 245896 409119 245898 409128
rect 245844 409090 245896 409096
rect 245844 406428 245896 406434
rect 245844 406370 245896 406376
rect 245856 405793 245884 406370
rect 245842 405784 245898 405793
rect 245842 405719 245898 405728
rect 245856 393314 245884 405719
rect 246316 399566 246344 527138
rect 246946 503024 247002 503033
rect 246946 502959 247002 502968
rect 246960 501634 246988 502959
rect 246948 501628 247000 501634
rect 246948 501570 247000 501576
rect 246394 442504 246450 442513
rect 246394 442439 246450 442448
rect 246304 399560 246356 399566
rect 246304 399502 246356 399508
rect 246408 394670 246436 442439
rect 247052 402966 247080 700266
rect 249800 610088 249852 610094
rect 249800 610030 249852 610036
rect 248512 588124 248564 588130
rect 248512 588066 248564 588072
rect 247776 585404 247828 585410
rect 247776 585346 247828 585352
rect 247684 585336 247736 585342
rect 247684 585278 247736 585284
rect 247696 484362 247724 585278
rect 247788 487830 247816 585346
rect 248418 557424 248474 557433
rect 248418 557359 248474 557368
rect 247776 487824 247828 487830
rect 247776 487766 247828 487772
rect 247684 484356 247736 484362
rect 247684 484298 247736 484304
rect 247684 482316 247736 482322
rect 247684 482258 247736 482264
rect 247040 402960 247092 402966
rect 247040 402902 247092 402908
rect 246578 399936 246634 399945
rect 246578 399871 246634 399880
rect 246396 394664 246448 394670
rect 246396 394606 246448 394612
rect 245764 393286 245884 393314
rect 245660 392012 245712 392018
rect 245660 391954 245712 391960
rect 245016 389224 245068 389230
rect 245016 389166 245068 389172
rect 244924 381676 244976 381682
rect 244924 381618 244976 381624
rect 245028 370734 245056 389166
rect 245660 371952 245712 371958
rect 245660 371894 245712 371900
rect 245016 370728 245068 370734
rect 245016 370670 245068 370676
rect 245672 368558 245700 371894
rect 245660 368552 245712 368558
rect 245660 368494 245712 368500
rect 244188 367804 244240 367810
rect 244188 367746 244240 367752
rect 242992 362228 243044 362234
rect 242992 362170 243044 362176
rect 243912 359712 243964 359718
rect 243912 359654 243964 359660
rect 243924 357474 243952 359654
rect 243912 357468 243964 357474
rect 243912 357410 243964 357416
rect 239508 355014 239936 355042
rect 241532 355014 241868 355042
rect 243924 354906 243952 357410
rect 245672 355314 245700 368494
rect 245764 365022 245792 393286
rect 246592 369170 246620 399871
rect 246948 394664 247000 394670
rect 246948 394606 247000 394612
rect 246580 369164 246632 369170
rect 246580 369106 246632 369112
rect 245752 365016 245804 365022
rect 245752 364958 245804 364964
rect 246960 363050 246988 394606
rect 245752 363044 245804 363050
rect 245752 362986 245804 362992
rect 246948 363044 247000 363050
rect 246948 362986 247000 362992
rect 245764 362302 245792 362986
rect 245752 362296 245804 362302
rect 245752 362238 245804 362244
rect 247696 357746 247724 482258
rect 247776 436144 247828 436150
rect 247776 436086 247828 436092
rect 247788 380254 247816 436086
rect 247776 380248 247828 380254
rect 247776 380190 247828 380196
rect 248432 359582 248460 557359
rect 248524 402286 248552 588066
rect 249706 557424 249762 557433
rect 249706 557359 249762 557368
rect 249720 556850 249748 557359
rect 249708 556844 249760 556850
rect 249708 556786 249760 556792
rect 249064 527876 249116 527882
rect 249064 527818 249116 527824
rect 249076 500546 249104 527818
rect 249064 500540 249116 500546
rect 249064 500482 249116 500488
rect 249064 489932 249116 489938
rect 249064 489874 249116 489880
rect 249076 404462 249104 489874
rect 249064 404456 249116 404462
rect 249064 404398 249116 404404
rect 249812 403850 249840 610030
rect 250444 560312 250496 560318
rect 250444 560254 250496 560260
rect 249800 403844 249852 403850
rect 249800 403786 249852 403792
rect 248512 402280 248564 402286
rect 248512 402222 248564 402228
rect 250456 370598 250484 560254
rect 250536 514820 250588 514826
rect 250536 514762 250588 514768
rect 250548 396846 250576 514762
rect 251100 509930 251128 702510
rect 267646 702471 267702 702480
rect 283852 702434 283880 703520
rect 300136 702642 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 702636 300176 702642
rect 300124 702578 300176 702584
rect 282932 702406 283880 702434
rect 269120 700392 269172 700398
rect 269120 700334 269172 700340
rect 261484 699712 261536 699718
rect 261484 699654 261536 699660
rect 260104 615528 260156 615534
rect 260104 615470 260156 615476
rect 253940 608728 253992 608734
rect 253940 608670 253992 608676
rect 252560 608660 252612 608666
rect 252560 608602 252612 608608
rect 251180 603288 251232 603294
rect 251180 603230 251232 603236
rect 251088 509924 251140 509930
rect 251088 509866 251140 509872
rect 251088 420232 251140 420238
rect 251088 420174 251140 420180
rect 250536 396840 250588 396846
rect 250536 396782 250588 396788
rect 250444 370592 250496 370598
rect 250444 370534 250496 370540
rect 251100 360398 251128 420174
rect 251192 400994 251220 603230
rect 252468 603220 252520 603226
rect 252468 603162 252520 603168
rect 251824 589484 251876 589490
rect 251824 589426 251876 589432
rect 251836 502994 251864 589426
rect 251824 502988 251876 502994
rect 251824 502930 251876 502936
rect 251916 425128 251968 425134
rect 251916 425070 251968 425076
rect 251824 422340 251876 422346
rect 251824 422282 251876 422288
rect 251180 400988 251232 400994
rect 251180 400930 251232 400936
rect 251836 373318 251864 422282
rect 251928 394602 251956 425070
rect 252480 403034 252508 603162
rect 252468 403028 252520 403034
rect 252468 402970 252520 402976
rect 252480 402898 252508 402970
rect 252468 402892 252520 402898
rect 252468 402834 252520 402840
rect 251916 394596 251968 394602
rect 251916 394538 251968 394544
rect 252468 394596 252520 394602
rect 252468 394538 252520 394544
rect 252480 393378 252508 394538
rect 252468 393372 252520 393378
rect 252468 393314 252520 393320
rect 252480 392698 252508 393314
rect 252468 392692 252520 392698
rect 252468 392634 252520 392640
rect 252572 378826 252600 608602
rect 253204 600500 253256 600506
rect 253204 600442 253256 600448
rect 253216 402830 253244 600442
rect 253296 588056 253348 588062
rect 253296 587998 253348 588004
rect 253308 485110 253336 587998
rect 253296 485104 253348 485110
rect 253296 485046 253348 485052
rect 253296 431996 253348 432002
rect 253296 431938 253348 431944
rect 253308 415410 253336 431938
rect 253296 415404 253348 415410
rect 253296 415346 253348 415352
rect 253952 403782 253980 608670
rect 256608 596216 256660 596222
rect 256608 596158 256660 596164
rect 255320 585200 255372 585206
rect 255320 585142 255372 585148
rect 255228 549296 255280 549302
rect 255228 549238 255280 549244
rect 255240 507414 255268 549238
rect 255228 507408 255280 507414
rect 255228 507350 255280 507356
rect 255332 505782 255360 585142
rect 255320 505776 255372 505782
rect 255320 505718 255372 505724
rect 255332 504422 255360 505718
rect 255320 504416 255372 504422
rect 255320 504358 255372 504364
rect 255320 465112 255372 465118
rect 255320 465054 255372 465060
rect 254584 449948 254636 449954
rect 254584 449890 254636 449896
rect 253940 403776 253992 403782
rect 253940 403718 253992 403724
rect 253204 402824 253256 402830
rect 253204 402766 253256 402772
rect 252560 378820 252612 378826
rect 252560 378762 252612 378768
rect 251824 373312 251876 373318
rect 251824 373254 251876 373260
rect 250536 360392 250588 360398
rect 250536 360334 250588 360340
rect 251088 360392 251140 360398
rect 251088 360334 251140 360340
rect 248420 359576 248472 359582
rect 248420 359518 248472 359524
rect 247684 357740 247736 357746
rect 247684 357682 247736 357688
rect 248144 357740 248196 357746
rect 248144 357682 248196 357688
rect 245672 355286 245746 355314
rect 245718 355028 245746 355286
rect 243800 354878 243952 354906
rect 248156 354770 248184 357682
rect 250548 355042 250576 360334
rect 254596 359650 254624 449890
rect 255332 386238 255360 465054
rect 256516 426488 256568 426494
rect 256516 426430 256568 426436
rect 255320 386232 255372 386238
rect 255320 386174 255372 386180
rect 255332 385694 255360 386174
rect 255320 385688 255372 385694
rect 255320 385630 255372 385636
rect 256528 369918 256556 426430
rect 255320 369912 255372 369918
rect 255320 369854 255372 369860
rect 256516 369912 256568 369918
rect 256516 369854 256568 369860
rect 255332 369238 255360 369854
rect 255320 369232 255372 369238
rect 255320 369174 255372 369180
rect 256620 367198 256648 596158
rect 257344 589416 257396 589422
rect 257344 589358 257396 589364
rect 257252 552696 257304 552702
rect 257252 552638 257304 552644
rect 257264 552090 257292 552638
rect 256700 552084 256752 552090
rect 256700 552026 256752 552032
rect 257252 552084 257304 552090
rect 257252 552026 257304 552032
rect 256712 377466 256740 552026
rect 256792 487824 256844 487830
rect 256792 487766 256844 487772
rect 256804 487218 256832 487766
rect 256792 487212 256844 487218
rect 256792 487154 256844 487160
rect 256804 396778 256832 487154
rect 257356 415410 257384 589358
rect 259460 509924 259512 509930
rect 259460 509866 259512 509872
rect 258080 507408 258132 507414
rect 258080 507350 258132 507356
rect 257344 415404 257396 415410
rect 257344 415346 257396 415352
rect 256792 396772 256844 396778
rect 256792 396714 256844 396720
rect 258092 391270 258120 507350
rect 259472 395418 259500 509866
rect 259460 395412 259512 395418
rect 259460 395354 259512 395360
rect 258080 391264 258132 391270
rect 258080 391206 258132 391212
rect 260116 384470 260144 615470
rect 260196 585268 260248 585274
rect 260196 585210 260248 585216
rect 260208 505782 260236 585210
rect 260196 505776 260248 505782
rect 260196 505718 260248 505724
rect 260748 395820 260800 395826
rect 260748 395762 260800 395768
rect 260760 395418 260788 395762
rect 260748 395412 260800 395418
rect 260748 395354 260800 395360
rect 260104 384464 260156 384470
rect 260104 384406 260156 384412
rect 256700 377460 256752 377466
rect 256700 377402 256752 377408
rect 259460 376780 259512 376786
rect 259460 376722 259512 376728
rect 255964 367192 256016 367198
rect 255964 367134 256016 367140
rect 256608 367192 256660 367198
rect 256608 367134 256660 367140
rect 254584 359644 254636 359650
rect 254584 359586 254636 359592
rect 255976 359514 256004 367134
rect 259472 364334 259500 376722
rect 261496 367878 261524 699654
rect 265624 698964 265676 698970
rect 265624 698906 265676 698912
rect 264244 614168 264296 614174
rect 264244 614110 264296 614116
rect 262220 569220 262272 569226
rect 262220 569162 262272 569168
rect 262232 568614 262260 569162
rect 262220 568608 262272 568614
rect 262220 568550 262272 568556
rect 261576 445800 261628 445806
rect 261576 445742 261628 445748
rect 260748 367872 260800 367878
rect 260748 367814 260800 367820
rect 261484 367872 261536 367878
rect 261484 367814 261536 367820
rect 259472 364306 260144 364334
rect 256700 362364 256752 362370
rect 256700 362306 256752 362312
rect 255964 359508 256016 359514
rect 255964 359450 256016 359456
rect 252466 357504 252522 357513
rect 251088 357468 251140 357474
rect 256712 357474 256740 362306
rect 258908 362228 258960 362234
rect 258908 362170 258960 362176
rect 252466 357439 252522 357448
rect 253940 357468 253992 357474
rect 251088 357410 251140 357416
rect 251100 356726 251128 357410
rect 251088 356720 251140 356726
rect 251088 356662 251140 356668
rect 252480 355042 252508 357439
rect 253940 357410 253992 357416
rect 256700 357468 256752 357474
rect 256700 357410 256752 357416
rect 250240 355014 250576 355042
rect 252172 355014 252508 355042
rect 253952 355042 253980 357410
rect 254400 355428 254452 355434
rect 254400 355370 254452 355376
rect 254412 355042 254440 355370
rect 256712 355314 256740 357410
rect 253952 355014 254440 355042
rect 256666 355286 256740 355314
rect 256666 355028 256694 355286
rect 258920 355042 258948 362170
rect 258612 355014 258948 355042
rect 260116 355042 260144 364306
rect 260760 360913 260788 367814
rect 260746 360904 260802 360913
rect 260746 360839 260802 360848
rect 261588 357406 261616 445742
rect 262232 394126 262260 568550
rect 262220 394120 262272 394126
rect 262220 394062 262272 394068
rect 262864 370660 262916 370666
rect 262864 370602 262916 370608
rect 262876 364334 262904 370602
rect 263600 367328 263652 367334
rect 263600 367270 263652 367276
rect 263612 366382 263640 367270
rect 263600 366376 263652 366382
rect 263600 366318 263652 366324
rect 264256 365158 264284 614110
rect 264336 546508 264388 546514
rect 264336 546450 264388 546456
rect 264348 532030 264376 546450
rect 264336 532024 264388 532030
rect 264336 531966 264388 531972
rect 264336 525836 264388 525842
rect 264336 525778 264388 525784
rect 264348 513330 264376 525778
rect 264336 513324 264388 513330
rect 264336 513266 264388 513272
rect 265532 456068 265584 456074
rect 265532 456010 265584 456016
rect 265544 455462 265572 456010
rect 264980 455456 265032 455462
rect 264980 455398 265032 455404
rect 265532 455456 265584 455462
rect 265532 455398 265584 455404
rect 264888 425128 264940 425134
rect 264888 425070 264940 425076
rect 264900 367334 264928 425070
rect 264992 374678 265020 455398
rect 265636 445806 265664 698906
rect 266360 587920 266412 587926
rect 266360 587862 266412 587868
rect 265716 495508 265768 495514
rect 265716 495450 265768 495456
rect 265624 445800 265676 445806
rect 265624 445742 265676 445748
rect 265728 397254 265756 495450
rect 265716 397248 265768 397254
rect 265716 397190 265768 397196
rect 265624 377664 265676 377670
rect 265624 377606 265676 377612
rect 264980 374672 265032 374678
rect 264980 374614 265032 374620
rect 264888 367328 264940 367334
rect 264888 367270 264940 367276
rect 264244 365152 264296 365158
rect 264244 365094 264296 365100
rect 262784 364306 262904 364334
rect 261576 357400 261628 357406
rect 261576 357342 261628 357348
rect 262128 357400 262180 357406
rect 262128 357342 262180 357348
rect 262140 356794 262168 357342
rect 262128 356788 262180 356794
rect 262128 356730 262180 356736
rect 262784 356318 262812 364306
rect 265636 357746 265664 377606
rect 262864 357740 262916 357746
rect 262864 357682 262916 357688
rect 265348 357740 265400 357746
rect 265348 357682 265400 357688
rect 265624 357740 265676 357746
rect 265624 357682 265676 357688
rect 262876 356726 262904 357682
rect 262864 356720 262916 356726
rect 262864 356662 262916 356668
rect 262772 356312 262824 356318
rect 262772 356254 262824 356260
rect 262784 355042 262812 356254
rect 265360 355042 265388 357682
rect 266372 356182 266400 587862
rect 269028 559564 269080 559570
rect 269028 559506 269080 559512
rect 269040 558958 269068 559506
rect 267740 558952 267792 558958
rect 267740 558894 267792 558900
rect 269028 558952 269080 558958
rect 269028 558894 269080 558900
rect 267752 389842 267780 558894
rect 269132 409154 269160 700334
rect 282932 620294 282960 702406
rect 300136 699718 300164 702578
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 282920 620288 282972 620294
rect 282920 620230 282972 620236
rect 289728 618316 289780 618322
rect 289728 618258 289780 618264
rect 288348 614236 288400 614242
rect 288348 614178 288400 614184
rect 275284 611516 275336 611522
rect 275284 611458 275336 611464
rect 273904 608796 273956 608802
rect 273904 608738 273956 608744
rect 271142 586392 271198 586401
rect 271142 586327 271198 586336
rect 269764 551336 269816 551342
rect 269764 551278 269816 551284
rect 269776 527134 269804 551278
rect 269764 527128 269816 527134
rect 269764 527070 269816 527076
rect 270500 518968 270552 518974
rect 270500 518910 270552 518916
rect 269764 491360 269816 491366
rect 269764 491302 269816 491308
rect 269212 472048 269264 472054
rect 269212 471990 269264 471996
rect 269224 468518 269252 471990
rect 269776 469198 269804 491302
rect 269764 469192 269816 469198
rect 269764 469134 269816 469140
rect 269212 468512 269264 468518
rect 269212 468454 269264 468460
rect 269120 409148 269172 409154
rect 269120 409090 269172 409096
rect 269764 409148 269816 409154
rect 269764 409090 269816 409096
rect 267740 389836 267792 389842
rect 267740 389778 267792 389784
rect 269776 380186 269804 409090
rect 270512 388482 270540 518910
rect 271156 409902 271184 586327
rect 271144 409896 271196 409902
rect 271144 409838 271196 409844
rect 271156 405074 271184 409838
rect 271144 405068 271196 405074
rect 271144 405010 271196 405016
rect 270500 388476 270552 388482
rect 270500 388418 270552 388424
rect 270500 387932 270552 387938
rect 270500 387874 270552 387880
rect 269764 380180 269816 380186
rect 269764 380122 269816 380128
rect 267740 374128 267792 374134
rect 267740 374070 267792 374076
rect 267752 364334 267780 374070
rect 267752 364306 268516 364334
rect 266360 356176 266412 356182
rect 266360 356118 266412 356124
rect 266820 356176 266872 356182
rect 266820 356118 266872 356124
rect 260116 355014 260544 355042
rect 262476 355014 262812 355042
rect 265052 355014 265388 355042
rect 266832 354770 266860 356118
rect 268488 355042 268516 364306
rect 270408 356176 270460 356182
rect 270408 356118 270460 356124
rect 270420 356046 270448 356118
rect 270408 356040 270460 356046
rect 270408 355982 270460 355988
rect 270512 355042 270540 387874
rect 273916 379642 273944 608738
rect 273996 590708 274048 590714
rect 273996 590650 274048 590656
rect 274008 396778 274036 590650
rect 273996 396772 274048 396778
rect 273996 396714 274048 396720
rect 273996 386436 274048 386442
rect 273996 386378 274048 386384
rect 273904 379636 273956 379642
rect 273904 379578 273956 379584
rect 273916 363866 273944 379578
rect 274008 365702 274036 386378
rect 275296 381614 275324 611458
rect 287704 604716 287756 604722
rect 287704 604658 287756 604664
rect 283564 602064 283616 602070
rect 283564 602006 283616 602012
rect 279424 597644 279476 597650
rect 279424 597586 279476 597592
rect 277400 586696 277452 586702
rect 277400 586638 277452 586644
rect 276020 578944 276072 578950
rect 276020 578886 276072 578892
rect 276032 578270 276060 578886
rect 276020 578264 276072 578270
rect 276020 578206 276072 578212
rect 276664 578264 276716 578270
rect 276664 578206 276716 578212
rect 275284 381608 275336 381614
rect 275284 381550 275336 381556
rect 274640 369980 274692 369986
rect 274640 369922 274692 369928
rect 273996 365696 274048 365702
rect 273996 365638 274048 365644
rect 274548 365696 274600 365702
rect 274548 365638 274600 365644
rect 273904 363860 273956 363866
rect 273904 363802 273956 363808
rect 274560 357406 274588 365638
rect 274652 364334 274680 369922
rect 274652 364306 274956 364334
rect 273720 357400 273772 357406
rect 273720 357342 273772 357348
rect 274548 357400 274600 357406
rect 274548 357342 274600 357348
rect 273732 356182 273760 357342
rect 273720 356176 273772 356182
rect 273720 356118 273772 356124
rect 273732 355042 273760 356118
rect 268488 355014 268916 355042
rect 270512 355014 271184 355042
rect 273424 355014 273760 355042
rect 274928 355042 274956 364306
rect 276676 358902 276704 578206
rect 276848 369844 276900 369850
rect 276848 369786 276900 369792
rect 276860 368558 276888 369786
rect 276848 368552 276900 368558
rect 276848 368494 276900 368500
rect 277308 368552 277360 368558
rect 277308 368494 277360 368500
rect 277320 363798 277348 368494
rect 277308 363792 277360 363798
rect 277308 363734 277360 363740
rect 277412 359718 277440 586638
rect 278044 496868 278096 496874
rect 278044 496810 278096 496816
rect 278056 369850 278084 496810
rect 279436 375358 279464 597586
rect 280804 474768 280856 474774
rect 280804 474710 280856 474716
rect 280068 458856 280120 458862
rect 280068 458798 280120 458804
rect 280080 458250 280108 458798
rect 279516 458244 279568 458250
rect 279516 458186 279568 458192
rect 280068 458244 280120 458250
rect 280068 458186 280120 458192
rect 279424 375352 279476 375358
rect 279424 375294 279476 375300
rect 278044 369844 278096 369850
rect 278044 369786 278096 369792
rect 277400 359712 277452 359718
rect 277400 359654 277452 359660
rect 279436 358902 279464 375294
rect 279528 365022 279556 458186
rect 280816 398313 280844 474710
rect 282828 429208 282880 429214
rect 282828 429150 282880 429156
rect 280802 398304 280858 398313
rect 280802 398239 280858 398248
rect 281446 398304 281502 398313
rect 281446 398239 281502 398248
rect 281460 370598 281488 398239
rect 281448 370592 281500 370598
rect 281448 370534 281500 370540
rect 279516 365016 279568 365022
rect 279516 364958 279568 364964
rect 276664 358896 276716 358902
rect 276664 358838 276716 358844
rect 277124 358896 277176 358902
rect 277124 358838 277176 358844
rect 279424 358896 279476 358902
rect 279424 358838 279476 358844
rect 274928 355014 275356 355042
rect 200118 354719 200174 354728
rect 209872 354748 209924 354754
rect 228836 354742 228988 354770
rect 248156 354742 248308 354770
rect 266832 354742 266984 354770
rect 271156 354754 271184 355014
rect 277136 354770 277164 358838
rect 279436 355042 279464 358838
rect 282840 358737 282868 429150
rect 283576 397322 283604 602006
rect 283656 438932 283708 438938
rect 283656 438874 283708 438880
rect 283564 397316 283616 397322
rect 283564 397258 283616 397264
rect 283668 365974 283696 438874
rect 286968 389836 287020 389842
rect 286968 389778 287020 389784
rect 283656 365968 283708 365974
rect 283656 365910 283708 365916
rect 282090 358728 282146 358737
rect 282090 358663 282146 358672
rect 282826 358728 282882 358737
rect 282826 358663 282882 358672
rect 282104 357649 282132 358663
rect 283668 357678 283696 365910
rect 286980 357814 287008 389778
rect 287716 379506 287744 604658
rect 288360 387258 288388 614178
rect 289084 612876 289136 612882
rect 289084 612818 289136 612824
rect 289096 433294 289124 612818
rect 289176 485852 289228 485858
rect 289176 485794 289228 485800
rect 288624 433288 288676 433294
rect 288624 433230 288676 433236
rect 289084 433288 289136 433294
rect 289084 433230 289136 433236
rect 288636 432614 288664 433230
rect 288624 432608 288676 432614
rect 288624 432550 288676 432556
rect 288636 431390 288664 432550
rect 288624 431384 288676 431390
rect 288624 431326 288676 431332
rect 288348 387252 288400 387258
rect 288348 387194 288400 387200
rect 287704 379500 287756 379506
rect 287704 379442 287756 379448
rect 287716 360874 287744 379442
rect 287704 360868 287756 360874
rect 287704 360810 287756 360816
rect 285956 357808 286008 357814
rect 285956 357750 286008 357756
rect 286968 357808 287020 357814
rect 286968 357750 287020 357756
rect 283656 357672 283708 357678
rect 282090 357640 282146 357649
rect 283656 357614 283708 357620
rect 282090 357575 282146 357584
rect 282104 355042 282132 357575
rect 285968 355042 285996 357750
rect 287336 357672 287388 357678
rect 287336 357614 287388 357620
rect 279068 355014 279464 355042
rect 281796 355014 282132 355042
rect 285660 355014 285996 355042
rect 287348 355042 287376 357614
rect 289188 355366 289216 485794
rect 289740 362234 289768 618258
rect 331232 616146 331260 702986
rect 332416 700324 332468 700330
rect 332416 700266 332468 700272
rect 331220 616140 331272 616146
rect 331220 616082 331272 616088
rect 300216 612808 300268 612814
rect 300216 612750 300268 612756
rect 292396 610156 292448 610162
rect 292396 610098 292448 610104
rect 290464 541000 290516 541006
rect 290464 540942 290516 540948
rect 290476 381546 290504 540942
rect 292408 393314 292436 610098
rect 295984 607300 296036 607306
rect 295984 607242 296036 607248
rect 293866 594960 293922 594969
rect 293866 594895 293922 594904
rect 292488 583772 292540 583778
rect 292488 583714 292540 583720
rect 292316 393286 292436 393314
rect 292028 392624 292080 392630
rect 292028 392566 292080 392572
rect 292040 392086 292068 392566
rect 292028 392080 292080 392086
rect 292028 392022 292080 392028
rect 292040 383654 292068 392022
rect 292316 392018 292344 393286
rect 292304 392012 292356 392018
rect 292304 391954 292356 391960
rect 292316 391338 292344 391954
rect 292304 391332 292356 391338
rect 292304 391274 292356 391280
rect 292040 383626 292344 383654
rect 290464 381540 290516 381546
rect 290464 381482 290516 381488
rect 291108 377460 291160 377466
rect 291108 377402 291160 377408
rect 291120 376786 291148 377402
rect 291108 376780 291160 376786
rect 291108 376722 291160 376728
rect 289728 362228 289780 362234
rect 289728 362170 289780 362176
rect 290464 358148 290516 358154
rect 290464 358090 290516 358096
rect 289176 355360 289228 355366
rect 289176 355302 289228 355308
rect 290476 355042 290504 358090
rect 291120 356017 291148 376722
rect 291200 360256 291252 360262
rect 291200 360198 291252 360204
rect 291106 356008 291162 356017
rect 291106 355943 291162 355952
rect 287348 355014 287592 355042
rect 290168 355014 290504 355042
rect 279068 354822 279096 355014
rect 279056 354816 279108 354822
rect 271144 354748 271196 354754
rect 209872 354690 209924 354696
rect 277136 354742 277288 354770
rect 284024 354816 284076 354822
rect 279056 354758 279108 354764
rect 283728 354764 284024 354770
rect 283728 354758 284076 354764
rect 283728 354742 284064 354758
rect 271144 354690 271196 354696
rect 291212 354657 291240 360198
rect 291842 355056 291898 355065
rect 291842 354991 291898 355000
rect 291856 354793 291884 354991
rect 292316 354958 292344 383626
rect 292304 354952 292356 354958
rect 292304 354894 292356 354900
rect 291842 354784 291898 354793
rect 291842 354719 291898 354728
rect 291198 354648 291254 354657
rect 292500 354634 292528 583714
rect 293880 464409 293908 594895
rect 295340 585132 295392 585138
rect 295340 585074 295392 585080
rect 295352 584662 295380 585074
rect 295996 584662 296024 607242
rect 298008 601996 298060 602002
rect 298008 601938 298060 601944
rect 295340 584656 295392 584662
rect 295340 584598 295392 584604
rect 295984 584656 296036 584662
rect 295984 584598 296036 584604
rect 293960 572008 294012 572014
rect 293960 571950 294012 571956
rect 293972 571334 294000 571950
rect 293960 571328 294012 571334
rect 293960 571270 294012 571276
rect 295248 571328 295300 571334
rect 295248 571270 295300 571276
rect 293866 464400 293922 464409
rect 293866 464335 293922 464344
rect 293960 462392 294012 462398
rect 293960 462334 294012 462340
rect 293972 461650 294000 462334
rect 293960 461644 294012 461650
rect 293960 461586 294012 461592
rect 293040 431384 293092 431390
rect 293040 431326 293092 431332
rect 292580 383036 292632 383042
rect 292580 382978 292632 382984
rect 292592 382226 292620 382978
rect 292580 382220 292632 382226
rect 292580 382162 292632 382168
rect 292580 354952 292632 354958
rect 292580 354894 292632 354900
rect 292592 354657 292620 354894
rect 292100 354606 292528 354634
rect 291198 354583 291254 354592
rect 292500 354550 292528 354606
rect 292578 354648 292634 354657
rect 292578 354583 292634 354592
rect 292488 354544 292540 354550
rect 292488 354486 292540 354492
rect 179878 350024 179934 350033
rect 179878 349959 179934 349968
rect 179510 314868 179566 314877
rect 179340 314826 179510 314854
rect 179340 314702 179368 314826
rect 179510 314803 179566 314812
rect 179328 314696 179380 314702
rect 179328 314638 179380 314644
rect 179510 308068 179566 308077
rect 179510 308003 179566 308012
rect 179234 292360 179290 292369
rect 179234 292295 179290 292304
rect 179144 204944 179196 204950
rect 179144 204886 179196 204892
rect 179248 87650 179276 292295
rect 179418 270600 179474 270609
rect 179418 270535 179474 270544
rect 179326 252920 179382 252929
rect 179326 252855 179382 252864
rect 179236 87644 179288 87650
rect 179236 87586 179288 87592
rect 179340 25702 179368 252855
rect 179432 35358 179460 270535
rect 179524 243545 179552 308003
rect 293052 277001 293080 431326
rect 293316 384328 293368 384334
rect 293316 384270 293368 384276
rect 293328 383042 293356 384270
rect 293316 383036 293368 383042
rect 293316 382978 293368 382984
rect 293132 382220 293184 382226
rect 293132 382162 293184 382168
rect 293144 331945 293172 382162
rect 293224 357604 293276 357610
rect 293224 357546 293276 357552
rect 293236 351218 293264 357546
rect 293316 354544 293368 354550
rect 293314 354512 293316 354521
rect 293368 354512 293370 354521
rect 293314 354447 293370 354456
rect 293224 351212 293276 351218
rect 293224 351154 293276 351160
rect 293130 331936 293186 331945
rect 293130 331871 293186 331880
rect 293866 331936 293922 331945
rect 293866 331871 293922 331880
rect 293880 331294 293908 331871
rect 293868 331288 293920 331294
rect 293868 331230 293920 331236
rect 293132 327072 293184 327078
rect 293132 327014 293184 327020
rect 293144 325825 293172 327014
rect 293130 325816 293186 325825
rect 293130 325751 293186 325760
rect 293038 276992 293094 277001
rect 293038 276927 293094 276936
rect 293052 276690 293080 276927
rect 293040 276684 293092 276690
rect 293040 276626 293092 276632
rect 179696 271856 179748 271862
rect 179696 271798 179748 271804
rect 179708 270677 179736 271798
rect 179694 270668 179750 270677
rect 179694 270603 179750 270612
rect 293038 258904 293094 258913
rect 293038 258839 293094 258848
rect 179510 243536 179566 243545
rect 179510 243471 179566 243480
rect 179880 242276 179932 242282
rect 179880 242218 179932 242224
rect 179512 240780 179564 240786
rect 179512 240722 179564 240728
rect 179524 238814 179552 240722
rect 179512 238808 179564 238814
rect 179512 238750 179564 238756
rect 179892 237182 179920 242218
rect 271142 240680 271198 240689
rect 184204 240644 184256 240650
rect 271198 240638 271828 240666
rect 271142 240615 271198 240624
rect 184204 240586 184256 240592
rect 182822 240272 182878 240281
rect 182822 240207 182878 240216
rect 180030 239850 180058 240108
rect 179984 239822 180058 239850
rect 180812 240094 181976 240122
rect 179880 237176 179932 237182
rect 179880 237118 179932 237124
rect 179984 219434 180012 239822
rect 179524 219406 180012 219434
rect 179420 35352 179472 35358
rect 179420 35294 179472 35300
rect 179328 25696 179380 25702
rect 179328 25638 179380 25644
rect 179524 16046 179552 219406
rect 180812 214441 180840 240094
rect 180798 214432 180854 214441
rect 180798 214367 180854 214376
rect 182086 214432 182142 214441
rect 182086 214367 182142 214376
rect 182100 214033 182128 214367
rect 182086 214024 182142 214033
rect 182086 213959 182142 213968
rect 182100 151094 182128 213959
rect 182088 151088 182140 151094
rect 182088 151030 182140 151036
rect 181444 135312 181496 135318
rect 181444 135254 181496 135260
rect 181456 94042 181484 135254
rect 181536 116000 181588 116006
rect 181536 115942 181588 115948
rect 181444 94036 181496 94042
rect 181444 93978 181496 93984
rect 181548 89486 181576 115942
rect 182836 105602 182864 240207
rect 183572 240094 183908 240122
rect 182916 139460 182968 139466
rect 182916 139402 182968 139408
rect 182824 105596 182876 105602
rect 182824 105538 182876 105544
rect 182928 92410 182956 139402
rect 183008 122936 183060 122942
rect 183008 122878 183060 122884
rect 182916 92404 182968 92410
rect 182916 92346 182968 92352
rect 181536 89480 181588 89486
rect 181536 89422 181588 89428
rect 183020 85338 183048 122878
rect 183008 85332 183060 85338
rect 183008 85274 183060 85280
rect 179512 16040 179564 16046
rect 179512 15982 179564 15988
rect 177948 13184 178000 13190
rect 177948 13126 178000 13132
rect 183572 11014 183600 240094
rect 184216 230314 184244 240586
rect 191944 240514 192280 240530
rect 191932 240508 192280 240514
rect 191984 240502 192280 240508
rect 191932 240450 191984 240456
rect 190196 240366 190348 240394
rect 184952 240094 185840 240122
rect 184204 230308 184256 230314
rect 184204 230250 184256 230256
rect 184204 129804 184256 129810
rect 184204 129746 184256 129752
rect 184216 86834 184244 129746
rect 184296 114572 184348 114578
rect 184296 114514 184348 114520
rect 184308 88194 184336 114514
rect 184296 88188 184348 88194
rect 184296 88130 184348 88136
rect 184204 86828 184256 86834
rect 184204 86770 184256 86776
rect 184952 67046 184980 240094
rect 187758 239850 187786 240108
rect 187712 239822 187786 239850
rect 185582 239592 185638 239601
rect 185582 239527 185638 239536
rect 185596 227594 185624 239527
rect 185584 227588 185636 227594
rect 185584 227530 185636 227536
rect 187712 222193 187740 239822
rect 190196 239154 190224 240366
rect 193232 240094 194212 240122
rect 196144 240094 196480 240122
rect 189080 239148 189132 239154
rect 189080 239090 189132 239096
rect 190184 239148 190236 239154
rect 190184 239090 190236 239096
rect 189092 238814 189120 239090
rect 189080 238808 189132 238814
rect 189080 238750 189132 238756
rect 189724 229900 189776 229906
rect 189724 229842 189776 229848
rect 187698 222184 187754 222193
rect 187698 222119 187754 222128
rect 188986 222184 189042 222193
rect 188986 222119 189042 222128
rect 185582 221504 185638 221513
rect 185582 221439 185638 221448
rect 185596 179382 185624 221439
rect 189000 220969 189028 222119
rect 188986 220960 189042 220969
rect 188986 220895 189042 220904
rect 185584 179376 185636 179382
rect 185584 179318 185636 179324
rect 185584 153264 185636 153270
rect 185584 153206 185636 153212
rect 185596 90710 185624 153206
rect 188344 146328 188396 146334
rect 188344 146270 188396 146276
rect 186964 128376 187016 128382
rect 186964 128318 187016 128324
rect 185676 116068 185728 116074
rect 185676 116010 185728 116016
rect 185584 90704 185636 90710
rect 185584 90646 185636 90652
rect 185688 82618 185716 116010
rect 185676 82612 185728 82618
rect 185676 82554 185728 82560
rect 185584 80708 185636 80714
rect 185584 80650 185636 80656
rect 184940 67040 184992 67046
rect 184940 66982 184992 66988
rect 183560 11008 183612 11014
rect 183560 10950 183612 10956
rect 175188 6316 175240 6322
rect 175188 6258 175240 6264
rect 185596 3466 185624 80650
rect 186976 78674 187004 128318
rect 188356 88126 188384 146270
rect 188436 117428 188488 117434
rect 188436 117370 188488 117376
rect 188344 88120 188396 88126
rect 188344 88062 188396 88068
rect 188448 81258 188476 117370
rect 188436 81252 188488 81258
rect 188436 81194 188488 81200
rect 186964 78668 187016 78674
rect 186964 78610 187016 78616
rect 189000 18698 189028 220895
rect 189736 185842 189764 229842
rect 193232 223514 193260 240094
rect 196452 238746 196480 240094
rect 198706 239850 198734 240108
rect 200132 240094 200652 240122
rect 201512 240094 202584 240122
rect 204516 240094 204852 240122
rect 198706 239822 198780 239850
rect 196440 238740 196492 238746
rect 196440 238682 196492 238688
rect 196452 238406 196480 238682
rect 196440 238400 196492 238406
rect 196440 238342 196492 238348
rect 193956 236768 194008 236774
rect 193956 236710 194008 236716
rect 193220 223508 193272 223514
rect 193220 223450 193272 223456
rect 193864 204332 193916 204338
rect 193864 204274 193916 204280
rect 192484 202360 192536 202366
rect 192484 202302 192536 202308
rect 189908 189100 189960 189106
rect 189908 189042 189960 189048
rect 189816 187740 189868 187746
rect 189816 187682 189868 187688
rect 189724 185836 189776 185842
rect 189724 185778 189776 185784
rect 189828 160002 189856 187682
rect 189920 161362 189948 189042
rect 189908 161356 189960 161362
rect 189908 161298 189960 161304
rect 189816 159996 189868 160002
rect 189816 159938 189868 159944
rect 191104 151904 191156 151910
rect 191104 151846 191156 151852
rect 189816 151836 189868 151842
rect 189816 151778 189868 151784
rect 189724 142180 189776 142186
rect 189724 142122 189776 142128
rect 189736 92478 189764 142122
rect 189828 109002 189856 151778
rect 189908 121576 189960 121582
rect 189908 121518 189960 121524
rect 189816 108996 189868 109002
rect 189816 108938 189868 108944
rect 189816 102196 189868 102202
rect 189816 102138 189868 102144
rect 189724 92472 189776 92478
rect 189724 92414 189776 92420
rect 189828 86970 189856 102138
rect 189816 86964 189868 86970
rect 189816 86906 189868 86912
rect 189920 83910 189948 121518
rect 191116 92274 191144 151846
rect 191196 103556 191248 103562
rect 191196 103498 191248 103504
rect 191104 92268 191156 92274
rect 191104 92210 191156 92216
rect 191208 85542 191236 103498
rect 192496 92478 192524 202302
rect 192576 143608 192628 143614
rect 192576 143550 192628 143556
rect 192484 92472 192536 92478
rect 192484 92414 192536 92420
rect 192588 90914 192616 143550
rect 192668 99476 192720 99482
rect 192668 99418 192720 99424
rect 192576 90908 192628 90914
rect 192576 90850 192628 90856
rect 192484 90364 192536 90370
rect 192484 90306 192536 90312
rect 191196 85536 191248 85542
rect 191196 85478 191248 85484
rect 189908 83904 189960 83910
rect 189908 83846 189960 83852
rect 188988 18692 189040 18698
rect 188988 18634 189040 18640
rect 192496 3534 192524 90306
rect 192680 78470 192708 99418
rect 193876 95198 193904 204274
rect 193968 202366 193996 236710
rect 198752 231742 198780 239822
rect 198740 231736 198792 231742
rect 198740 231678 198792 231684
rect 199384 231736 199436 231742
rect 199384 231678 199436 231684
rect 194508 223508 194560 223514
rect 194508 223450 194560 223456
rect 194520 223378 194548 223450
rect 194508 223372 194560 223378
rect 194508 223314 194560 223320
rect 193956 202360 194008 202366
rect 193956 202302 194008 202308
rect 194048 150476 194100 150482
rect 194048 150418 194100 150424
rect 193956 138032 194008 138038
rect 193956 137974 194008 137980
rect 193864 95192 193916 95198
rect 193864 95134 193916 95140
rect 193968 86766 193996 137974
rect 194060 110430 194088 150418
rect 194520 140078 194548 223314
rect 196624 223032 196676 223038
rect 196624 222974 196676 222980
rect 196636 201006 196664 222974
rect 196624 201000 196676 201006
rect 196624 200942 196676 200948
rect 198004 191276 198056 191282
rect 198004 191218 198056 191224
rect 196624 186380 196676 186386
rect 196624 186322 196676 186328
rect 196636 164150 196664 186322
rect 196624 164144 196676 164150
rect 196624 164086 196676 164092
rect 195244 153332 195296 153338
rect 195244 153274 195296 153280
rect 194508 140072 194560 140078
rect 194508 140014 194560 140020
rect 194048 110424 194100 110430
rect 194048 110366 194100 110372
rect 194048 106344 194100 106350
rect 194048 106286 194100 106292
rect 193956 86760 194008 86766
rect 193956 86702 194008 86708
rect 194060 80034 194088 106286
rect 195256 93362 195284 153274
rect 196716 150544 196768 150550
rect 196716 150486 196768 150492
rect 196624 140820 196676 140826
rect 196624 140762 196676 140768
rect 195336 103624 195388 103630
rect 195336 103566 195388 103572
rect 195244 93356 195296 93362
rect 195244 93298 195296 93304
rect 194048 80028 194100 80034
rect 194048 79970 194100 79976
rect 192668 78464 192720 78470
rect 192668 78406 192720 78412
rect 195348 74526 195376 103566
rect 196636 83842 196664 140762
rect 196728 111790 196756 150486
rect 196716 111784 196768 111790
rect 196716 111726 196768 111732
rect 196808 104916 196860 104922
rect 196808 104858 196860 104864
rect 196716 100768 196768 100774
rect 196716 100710 196768 100716
rect 196624 83836 196676 83842
rect 196624 83778 196676 83784
rect 196728 75886 196756 100710
rect 196820 95062 196848 104858
rect 196808 95056 196860 95062
rect 196808 94998 196860 95004
rect 196716 75880 196768 75886
rect 196716 75822 196768 75828
rect 195336 74520 195388 74526
rect 195336 74462 195388 74468
rect 198016 61538 198044 191218
rect 198096 113280 198148 113286
rect 198096 113222 198148 113228
rect 198108 73166 198136 113222
rect 198188 104984 198240 104990
rect 198188 104926 198240 104932
rect 198200 93838 198228 104926
rect 198188 93832 198240 93838
rect 198188 93774 198240 93780
rect 199396 83502 199424 231678
rect 199384 83496 199436 83502
rect 199384 83438 199436 83444
rect 198096 73160 198148 73166
rect 198096 73102 198148 73108
rect 198004 61532 198056 61538
rect 198004 61474 198056 61480
rect 200132 27606 200160 240094
rect 200764 125656 200816 125662
rect 200764 125598 200816 125604
rect 200776 93974 200804 125598
rect 200764 93968 200816 93974
rect 200764 93910 200816 93916
rect 201512 31210 201540 240094
rect 204824 238746 204852 240094
rect 207078 239850 207106 240108
rect 207032 239822 207106 239850
rect 208412 240094 209024 240122
rect 210620 240094 210956 240122
rect 212552 240094 212888 240122
rect 215312 240094 215464 240122
rect 216692 240094 217396 240122
rect 204812 238740 204864 238746
rect 204812 238682 204864 238688
rect 204824 237182 204852 238682
rect 204812 237176 204864 237182
rect 204812 237118 204864 237124
rect 203524 229832 203576 229838
rect 203524 229774 203576 229780
rect 202144 213512 202196 213518
rect 202144 213454 202196 213460
rect 202156 95130 202184 213454
rect 203536 189990 203564 229774
rect 203524 189984 203576 189990
rect 203524 189926 203576 189932
rect 203524 187128 203576 187134
rect 203524 187070 203576 187076
rect 202236 135380 202288 135386
rect 202236 135322 202288 135328
rect 202144 95124 202196 95130
rect 202144 95066 202196 95072
rect 202248 77178 202276 135322
rect 202328 111920 202380 111926
rect 202328 111862 202380 111868
rect 202340 84114 202368 111862
rect 202328 84108 202380 84114
rect 202328 84050 202380 84056
rect 202236 77172 202288 77178
rect 202236 77114 202288 77120
rect 201500 31204 201552 31210
rect 201500 31146 201552 31152
rect 200120 27600 200172 27606
rect 200120 27542 200172 27548
rect 203536 3670 203564 187070
rect 206376 178356 206428 178362
rect 206376 178298 206428 178304
rect 204904 151972 204956 151978
rect 204904 151914 204956 151920
rect 203616 125724 203668 125730
rect 203616 125666 203668 125672
rect 203628 82686 203656 125666
rect 203708 114640 203760 114646
rect 203708 114582 203760 114588
rect 203616 82680 203668 82686
rect 203616 82622 203668 82628
rect 203720 75818 203748 114582
rect 204916 89418 204944 151914
rect 206284 151088 206336 151094
rect 206284 151030 206336 151036
rect 204996 106412 205048 106418
rect 204996 106354 205048 106360
rect 204904 89412 204956 89418
rect 204904 89354 204956 89360
rect 205008 81394 205036 106354
rect 204996 81388 205048 81394
rect 204996 81330 205048 81336
rect 203708 75812 203760 75818
rect 203708 75754 203760 75760
rect 203524 3664 203576 3670
rect 203524 3606 203576 3612
rect 192484 3528 192536 3534
rect 192484 3470 192536 3476
rect 206296 3466 206324 151030
rect 206388 149054 206416 178298
rect 206376 149048 206428 149054
rect 206376 148990 206428 148996
rect 206376 140888 206428 140894
rect 206376 140830 206428 140836
rect 206388 78538 206416 140830
rect 206468 120216 206520 120222
rect 206468 120158 206520 120164
rect 206480 89622 206508 120158
rect 206468 89616 206520 89622
rect 206468 89558 206520 89564
rect 206376 78532 206428 78538
rect 206376 78474 206428 78480
rect 207032 35290 207060 239822
rect 208412 220833 208440 240094
rect 210516 238944 210568 238950
rect 210516 238886 210568 238892
rect 208492 238060 208544 238066
rect 208492 238002 208544 238008
rect 208504 237454 208532 238002
rect 208492 237448 208544 237454
rect 208492 237390 208544 237396
rect 209688 237448 209740 237454
rect 209688 237390 209740 237396
rect 209700 223514 209728 237390
rect 210424 233980 210476 233986
rect 210424 233922 210476 233928
rect 209688 223508 209740 223514
rect 209688 223450 209740 223456
rect 208398 220824 208454 220833
rect 208398 220759 208454 220768
rect 209686 220824 209742 220833
rect 209686 220759 209742 220768
rect 207756 135448 207808 135454
rect 207756 135390 207808 135396
rect 207664 132592 207716 132598
rect 207664 132534 207716 132540
rect 207676 82754 207704 132534
rect 207768 92313 207796 135390
rect 209044 102264 209096 102270
rect 209044 102206 209096 102212
rect 207754 92304 207810 92313
rect 207754 92239 207810 92248
rect 209056 90982 209084 102206
rect 209136 96688 209188 96694
rect 209136 96630 209188 96636
rect 209044 90976 209096 90982
rect 209044 90918 209096 90924
rect 209148 89690 209176 96630
rect 209136 89684 209188 89690
rect 209136 89626 209188 89632
rect 207664 82748 207716 82754
rect 207664 82690 207716 82696
rect 209700 38622 209728 220759
rect 210436 211138 210464 233922
rect 210528 226166 210556 238886
rect 210620 237454 210648 240094
rect 210608 237448 210660 237454
rect 210608 237390 210660 237396
rect 211802 227080 211858 227089
rect 211802 227015 211858 227024
rect 210516 226160 210568 226166
rect 210516 226102 210568 226108
rect 210516 218884 210568 218890
rect 210516 218826 210568 218832
rect 210424 211132 210476 211138
rect 210424 211074 210476 211080
rect 210422 199336 210478 199345
rect 210422 199271 210478 199280
rect 209688 38616 209740 38622
rect 209688 38558 209740 38564
rect 207020 35284 207072 35290
rect 207020 35226 207072 35232
rect 210436 17406 210464 199271
rect 210528 180198 210556 218826
rect 211816 184249 211844 227015
rect 211896 211880 211948 211886
rect 211896 211822 211948 211828
rect 211802 184240 211858 184249
rect 211802 184175 211858 184184
rect 211908 183190 211936 211822
rect 212552 191826 212580 240094
rect 214562 239456 214618 239465
rect 214562 239391 214618 239400
rect 214576 231742 214604 239391
rect 215312 238882 215340 240094
rect 215300 238876 215352 238882
rect 215300 238818 215352 238824
rect 215944 234048 215996 234054
rect 215944 233990 215996 233996
rect 214564 231736 214616 231742
rect 214564 231678 214616 231684
rect 214564 225616 214616 225622
rect 214564 225558 214616 225564
rect 212540 191820 212592 191826
rect 212540 191762 212592 191768
rect 214576 188698 214604 225558
rect 214564 188692 214616 188698
rect 214564 188634 214616 188640
rect 214564 186448 214616 186454
rect 214564 186390 214616 186396
rect 211896 183184 211948 183190
rect 211896 183126 211948 183132
rect 210516 180192 210568 180198
rect 210516 180134 210568 180140
rect 211896 179444 211948 179450
rect 211896 179386 211948 179392
rect 211804 171148 211856 171154
rect 211804 171090 211856 171096
rect 211816 150414 211844 171090
rect 211908 162858 211936 179386
rect 214104 178152 214156 178158
rect 214104 178094 214156 178100
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 214012 175228 214064 175234
rect 214012 175170 214064 175176
rect 213920 175160 213972 175166
rect 213920 175102 213972 175108
rect 213932 175001 213960 175102
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175170
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173641 213960 173810
rect 213918 173632 213974 173641
rect 213918 173567 213974 173576
rect 214116 172961 214144 178094
rect 214102 172952 214158 172961
rect 214102 172887 214158 172896
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172281 213960 172450
rect 214012 172440 214064 172446
rect 214012 172382 214064 172388
rect 213918 172272 213974 172281
rect 213918 172207 213974 172216
rect 214024 171601 214052 172382
rect 214010 171592 214066 171601
rect 214010 171527 214066 171536
rect 213920 171080 213972 171086
rect 213918 171048 213920 171057
rect 213972 171048 213974 171057
rect 213918 170983 213974 170992
rect 213920 169720 213972 169726
rect 213918 169688 213920 169697
rect 213972 169688 213974 169697
rect 213918 169623 213974 169632
rect 214012 169652 214064 169658
rect 214012 169594 214064 169600
rect 214024 169017 214052 169594
rect 214010 169008 214066 169017
rect 214010 168943 214066 168952
rect 213920 168360 213972 168366
rect 213918 168328 213920 168337
rect 213972 168328 213974 168337
rect 213918 168263 213974 168272
rect 214012 168292 214064 168298
rect 214012 168234 214064 168240
rect 214024 167657 214052 168234
rect 214010 167648 214066 167657
rect 214010 167583 214066 167592
rect 214104 167000 214156 167006
rect 213918 166968 213974 166977
rect 214104 166942 214156 166948
rect 213918 166903 213920 166912
rect 213972 166903 213974 166912
rect 213920 166874 213972 166880
rect 214012 166864 214064 166870
rect 214012 166806 214064 166812
rect 214024 165753 214052 166806
rect 214116 166433 214144 166942
rect 214102 166424 214158 166433
rect 214102 166359 214158 166368
rect 214010 165744 214066 165753
rect 214010 165679 214066 165688
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165073 213960 165514
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214012 164212 214064 164218
rect 214012 164154 214064 164160
rect 213920 164144 213972 164150
rect 213920 164086 213972 164092
rect 213932 163713 213960 164086
rect 213918 163704 213974 163713
rect 213918 163639 213974 163648
rect 214024 163033 214052 164154
rect 214010 163024 214066 163033
rect 214010 162959 214066 162968
rect 211896 162852 211948 162858
rect 211896 162794 211948 162800
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 161809 213960 162794
rect 213918 161800 213974 161809
rect 213918 161735 213974 161744
rect 213920 161424 213972 161430
rect 213920 161366 213972 161372
rect 213932 161129 213960 161366
rect 214012 161356 214064 161362
rect 214012 161298 214064 161304
rect 213918 161120 213974 161129
rect 213918 161055 213974 161064
rect 214024 160449 214052 161298
rect 214010 160440 214066 160449
rect 214010 160375 214066 160384
rect 214012 160064 214064 160070
rect 214012 160006 214064 160012
rect 213920 159996 213972 160002
rect 213920 159938 213972 159944
rect 213932 159769 213960 159938
rect 213918 159760 213974 159769
rect 213918 159695 213974 159704
rect 214024 159089 214052 160006
rect 214104 159384 214156 159390
rect 214104 159326 214156 159332
rect 214010 159080 214066 159089
rect 214010 159015 214066 159024
rect 213458 157856 213514 157865
rect 213458 157791 213514 157800
rect 213472 157457 213500 157791
rect 213458 157448 213514 157457
rect 213458 157383 213514 157392
rect 213920 157344 213972 157350
rect 213920 157286 213972 157292
rect 213932 156505 213960 157286
rect 214116 157185 214144 159326
rect 214102 157176 214158 157185
rect 214102 157111 214158 157120
rect 213918 156496 213974 156505
rect 213918 156431 213974 156440
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155825 213960 155858
rect 213918 155816 213974 155825
rect 213918 155751 213974 155760
rect 214576 155145 214604 186390
rect 215956 180266 215984 233990
rect 215944 180260 215996 180266
rect 215944 180202 215996 180208
rect 214656 179512 214708 179518
rect 214656 179454 214708 179460
rect 214562 155136 214618 155145
rect 214562 155071 214618 155080
rect 214010 154456 214066 154465
rect 214010 154391 214066 154400
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 213932 153270 213960 153711
rect 214024 153338 214052 154391
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 213918 153096 213974 153105
rect 213918 153031 213974 153040
rect 213932 151978 213960 153031
rect 214010 152552 214066 152561
rect 214010 152487 214066 152496
rect 213920 151972 213972 151978
rect 213920 151914 213972 151920
rect 214024 151910 214052 152487
rect 214012 151904 214064 151910
rect 213918 151872 213974 151881
rect 214012 151846 214064 151852
rect 213918 151807 213920 151816
rect 213972 151807 213974 151816
rect 213920 151778 213972 151784
rect 214010 151192 214066 151201
rect 214010 151127 214066 151136
rect 213920 150544 213972 150550
rect 213918 150512 213920 150521
rect 213972 150512 213974 150521
rect 214024 150482 214052 151127
rect 213918 150447 213974 150456
rect 214012 150476 214064 150482
rect 214012 150418 214064 150424
rect 211804 150408 211856 150414
rect 211804 150350 211856 150356
rect 213920 150408 213972 150414
rect 213920 150350 213972 150356
rect 213932 149161 213960 150350
rect 214668 149841 214696 179454
rect 216588 178764 216640 178770
rect 216588 178706 216640 178712
rect 214932 178084 214984 178090
rect 214932 178026 214984 178032
rect 214944 170377 214972 178026
rect 214930 170368 214986 170377
rect 214930 170303 214986 170312
rect 214654 149832 214710 149841
rect 214654 149767 214710 149776
rect 213918 149152 213974 149161
rect 213918 149087 213974 149096
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148481 213960 148990
rect 213918 148472 213974 148481
rect 213918 148407 213974 148416
rect 214562 147928 214618 147937
rect 214562 147863 214618 147872
rect 213918 147248 213974 147257
rect 213918 147183 213974 147192
rect 213932 146334 213960 147183
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 214010 145888 214066 145897
rect 214010 145823 214066 145832
rect 213918 145208 213974 145217
rect 213918 145143 213974 145152
rect 213932 145042 213960 145143
rect 213920 145036 213972 145042
rect 213920 144978 213972 144984
rect 214024 144974 214052 145823
rect 214012 144968 214064 144974
rect 214012 144910 214064 144916
rect 213918 144528 213974 144537
rect 213918 144463 213974 144472
rect 213932 143614 213960 144463
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 213918 143304 213974 143313
rect 213918 143239 213974 143248
rect 213932 142730 213960 143239
rect 211804 142724 211856 142730
rect 211804 142666 211856 142672
rect 213920 142724 213972 142730
rect 213920 142666 213972 142672
rect 210516 136740 210568 136746
rect 210516 136682 210568 136688
rect 210528 79966 210556 136682
rect 211160 95260 211212 95266
rect 211160 95202 211212 95208
rect 211172 88330 211200 95202
rect 211160 88324 211212 88330
rect 211160 88266 211212 88272
rect 211816 81326 211844 142666
rect 213918 142624 213974 142633
rect 213918 142559 213974 142568
rect 213932 142186 213960 142559
rect 213920 142180 213972 142186
rect 213920 142122 213972 142128
rect 214010 141944 214066 141953
rect 214010 141879 214066 141888
rect 213918 141264 213974 141273
rect 213918 141199 213974 141208
rect 213932 140894 213960 141199
rect 213920 140888 213972 140894
rect 213920 140830 213972 140836
rect 214024 140826 214052 141879
rect 214012 140820 214064 140826
rect 214012 140762 214064 140768
rect 213182 140584 213238 140593
rect 213182 140519 213238 140528
rect 211896 118856 211948 118862
rect 211896 118798 211948 118804
rect 211908 86902 211936 118798
rect 211988 105052 212040 105058
rect 211988 104994 212040 105000
rect 211896 86896 211948 86902
rect 211896 86838 211948 86844
rect 212000 85474 212028 104994
rect 211988 85468 212040 85474
rect 211988 85410 212040 85416
rect 211804 81320 211856 81326
rect 211804 81262 211856 81268
rect 210516 79960 210568 79966
rect 210516 79902 210568 79908
rect 213196 79898 213224 140519
rect 213918 139904 213974 139913
rect 213918 139839 213974 139848
rect 213932 139466 213960 139839
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 213918 138680 213974 138689
rect 213918 138615 213974 138624
rect 213932 138038 213960 138615
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 214102 138000 214158 138009
rect 214102 137935 214158 137944
rect 213918 137320 213974 137329
rect 213918 137255 213974 137264
rect 213932 136746 213960 137255
rect 213920 136740 213972 136746
rect 213920 136682 213972 136688
rect 214116 136678 214144 137935
rect 214104 136672 214156 136678
rect 214010 136640 214066 136649
rect 214104 136614 214156 136620
rect 214010 136575 214066 136584
rect 214024 135454 214052 136575
rect 214102 135960 214158 135969
rect 214102 135895 214158 135904
rect 214012 135448 214064 135454
rect 214012 135390 214064 135396
rect 213920 135380 213972 135386
rect 213920 135322 213972 135328
rect 213932 135289 213960 135322
rect 214116 135318 214144 135895
rect 214104 135312 214156 135318
rect 213918 135280 213974 135289
rect 214104 135254 214156 135260
rect 213918 135215 213974 135224
rect 214010 134600 214066 134609
rect 214010 134535 214066 134544
rect 214024 134026 214052 134535
rect 214012 134020 214064 134026
rect 214012 133962 214064 133968
rect 213920 133952 213972 133958
rect 213918 133920 213920 133929
rect 213972 133920 213974 133929
rect 213918 133855 213974 133864
rect 214010 133376 214066 133385
rect 214010 133311 214066 133320
rect 213918 132696 213974 132705
rect 213918 132631 213974 132640
rect 213932 132530 213960 132631
rect 214024 132598 214052 133311
rect 214012 132592 214064 132598
rect 214012 132534 214064 132540
rect 213920 132524 213972 132530
rect 213920 132466 213972 132472
rect 213274 131336 213330 131345
rect 213274 131271 213330 131280
rect 213288 84182 213316 131271
rect 213918 130656 213974 130665
rect 213918 130591 213974 130600
rect 213932 129810 213960 130591
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 213918 128752 213974 128761
rect 213918 128687 213974 128696
rect 213932 128382 213960 128687
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 213918 127392 213974 127401
rect 213918 127327 213974 127336
rect 213932 127022 213960 127327
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 214010 126712 214066 126721
rect 214010 126647 214066 126656
rect 213918 126032 213974 126041
rect 213918 125967 213974 125976
rect 213932 125730 213960 125967
rect 213920 125724 213972 125730
rect 213920 125666 213972 125672
rect 214024 125662 214052 126647
rect 214012 125656 214064 125662
rect 214012 125598 214064 125604
rect 214010 125352 214066 125361
rect 214010 125287 214066 125296
rect 213918 124672 213974 124681
rect 213918 124607 213974 124616
rect 213932 124234 213960 124607
rect 214024 124302 214052 125287
rect 214012 124296 214064 124302
rect 214012 124238 214064 124244
rect 213920 124228 213972 124234
rect 213920 124170 213972 124176
rect 214010 124128 214066 124137
rect 214010 124063 214066 124072
rect 213918 123448 213974 123457
rect 213918 123383 213974 123392
rect 213932 122874 213960 123383
rect 214024 122942 214052 124063
rect 214012 122936 214064 122942
rect 214012 122878 214064 122884
rect 213920 122868 213972 122874
rect 213920 122810 213972 122816
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121582 213960 122023
rect 213920 121576 213972 121582
rect 213920 121518 213972 121524
rect 214024 121514 214052 122703
rect 214012 121508 214064 121514
rect 214012 121450 214064 121456
rect 214010 121408 214066 121417
rect 214010 121343 214066 121352
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120154 213960 120663
rect 214024 120222 214052 121343
rect 214012 120216 214064 120222
rect 214012 120158 214064 120164
rect 213920 120148 213972 120154
rect 213920 120090 213972 120096
rect 214010 120048 214066 120057
rect 214010 119983 214066 119992
rect 213918 119504 213974 119513
rect 213918 119439 213974 119448
rect 213932 118794 213960 119439
rect 213920 118788 213972 118794
rect 213920 118730 213972 118736
rect 214024 118726 214052 119983
rect 214104 118856 214156 118862
rect 214102 118824 214104 118833
rect 214156 118824 214158 118833
rect 214102 118759 214158 118768
rect 214012 118720 214064 118726
rect 214012 118662 214064 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 214024 117434 214052 118079
rect 213918 117399 213974 117408
rect 214012 117428 214064 117434
rect 213932 117366 213960 117399
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213920 117302 213972 117308
rect 214010 116784 214066 116793
rect 214010 116719 214066 116728
rect 213918 116104 213974 116113
rect 213918 116039 213920 116048
rect 213972 116039 213974 116048
rect 213920 116010 213972 116016
rect 214024 116006 214052 116719
rect 214012 116000 214064 116006
rect 214012 115942 214064 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114578 213960 114815
rect 214024 114646 214052 115359
rect 214012 114640 214064 114646
rect 214012 114582 214064 114588
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 214010 114200 214066 114209
rect 214010 114135 214066 114144
rect 213918 113520 213974 113529
rect 213918 113455 213974 113464
rect 213932 113218 213960 113455
rect 214024 113286 214052 114135
rect 214012 113280 214064 113286
rect 214012 113222 214064 113228
rect 213920 113212 213972 113218
rect 213920 113154 213972 113160
rect 214010 112840 214066 112849
rect 214010 112775 214066 112784
rect 213918 112160 213974 112169
rect 213918 112095 213974 112104
rect 213932 111858 213960 112095
rect 214024 111926 214052 112775
rect 214012 111920 214064 111926
rect 214012 111862 214064 111868
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 213918 111480 213974 111489
rect 213918 111415 213974 111424
rect 213932 110498 213960 111415
rect 213920 110492 213972 110498
rect 213920 110434 213972 110440
rect 214010 110256 214066 110265
rect 214010 110191 214066 110200
rect 213918 109576 213974 109585
rect 213918 109511 213974 109520
rect 213932 109070 213960 109511
rect 214024 109138 214052 110191
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107710 213960 108151
rect 214024 107778 214052 108831
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 107536 214066 107545
rect 214010 107471 214066 107480
rect 213918 106856 213974 106865
rect 213918 106791 213974 106800
rect 213932 106350 213960 106791
rect 214024 106418 214052 107471
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 213918 106176 213974 106185
rect 213918 106111 213974 106120
rect 213932 105058 213960 106111
rect 214010 105632 214066 105641
rect 214010 105567 214066 105576
rect 213920 105052 213972 105058
rect 213920 104994 213972 105000
rect 214024 104990 214052 105567
rect 214012 104984 214064 104990
rect 213918 104952 213974 104961
rect 214012 104926 214064 104932
rect 213918 104887 213920 104896
rect 213972 104887 213974 104896
rect 213920 104858 213972 104864
rect 214010 104272 214066 104281
rect 214010 104207 214066 104216
rect 214024 103630 214052 104207
rect 214012 103624 214064 103630
rect 213918 103592 213974 103601
rect 214012 103566 214064 103572
rect 213918 103527 213920 103536
rect 213972 103527 213974 103536
rect 213920 103498 213972 103504
rect 214010 102912 214066 102921
rect 214010 102847 214066 102856
rect 214024 102270 214052 102847
rect 214012 102264 214064 102270
rect 213918 102232 213974 102241
rect 214012 102206 214064 102212
rect 213918 102167 213920 102176
rect 213972 102167 213974 102176
rect 213920 102138 213972 102144
rect 214576 101454 214604 147863
rect 214654 146568 214710 146577
rect 214654 146503 214710 146512
rect 214668 102814 214696 146503
rect 215944 140072 215996 140078
rect 215944 140014 215996 140020
rect 214838 128072 214894 128081
rect 214838 128007 214894 128016
rect 214852 113174 214880 128007
rect 214852 113146 214972 113174
rect 214746 110800 214802 110809
rect 214746 110735 214802 110744
rect 214656 102808 214708 102814
rect 214656 102750 214708 102756
rect 214564 101448 214616 101454
rect 214564 101390 214616 101396
rect 213918 101008 213974 101017
rect 213918 100943 213974 100952
rect 213932 100774 213960 100943
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214010 100328 214066 100337
rect 214010 100263 214066 100272
rect 213918 99648 213974 99657
rect 213918 99583 213974 99592
rect 213932 99482 213960 99583
rect 213920 99476 213972 99482
rect 213920 99418 213972 99424
rect 214024 99414 214052 100263
rect 214012 99408 214064 99414
rect 214012 99350 214064 99356
rect 214010 98968 214066 98977
rect 214010 98903 214066 98912
rect 213918 98288 213974 98297
rect 213918 98223 213974 98232
rect 213932 98054 213960 98223
rect 214024 98122 214052 98903
rect 214012 98116 214064 98122
rect 214012 98058 214064 98064
rect 213920 98048 213972 98054
rect 213920 97990 213972 97996
rect 213918 97608 213974 97617
rect 213918 97543 213974 97552
rect 213932 96694 213960 97543
rect 214562 96928 214618 96937
rect 214562 96863 214618 96872
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 213918 96384 213974 96393
rect 213918 96319 213974 96328
rect 213932 95266 213960 96319
rect 213920 95260 213972 95266
rect 213920 95202 213972 95208
rect 214576 91050 214604 96863
rect 214564 91044 214616 91050
rect 214564 90986 214616 90992
rect 214562 89040 214618 89049
rect 214562 88975 214618 88984
rect 213276 84176 213328 84182
rect 213276 84118 213328 84124
rect 213184 79892 213236 79898
rect 213184 79834 213236 79840
rect 210424 17400 210476 17406
rect 210424 17342 210476 17348
rect 214576 3602 214604 88975
rect 214760 77246 214788 110735
rect 214944 93158 214972 113146
rect 215022 101552 215078 101561
rect 215022 101487 215078 101496
rect 214932 93152 214984 93158
rect 214932 93094 214984 93100
rect 215036 89729 215064 101487
rect 215022 89720 215078 89729
rect 215022 89655 215078 89664
rect 214748 77240 214800 77246
rect 214748 77182 214800 77188
rect 215956 4146 215984 140014
rect 216036 105596 216088 105602
rect 216036 105538 216088 105544
rect 216048 47734 216076 105538
rect 216600 90438 216628 178706
rect 216588 90432 216640 90438
rect 216588 90374 216640 90380
rect 216036 47728 216088 47734
rect 216036 47670 216088 47676
rect 216692 38010 216720 240094
rect 219314 239850 219342 240108
rect 221260 240094 221596 240122
rect 219314 239822 219388 239850
rect 219360 238610 219388 239822
rect 220176 239488 220228 239494
rect 220176 239430 220228 239436
rect 219440 238944 219492 238950
rect 219440 238886 219492 238892
rect 219348 238604 219400 238610
rect 219348 238546 219400 238552
rect 219452 238406 219480 238886
rect 219440 238400 219492 238406
rect 219440 238342 219492 238348
rect 220188 231130 220216 239430
rect 221568 233986 221596 240094
rect 223822 239850 223850 240108
rect 223776 239822 223850 239850
rect 224972 240094 225768 240122
rect 223776 238814 223804 239822
rect 223764 238808 223816 238814
rect 223764 238750 223816 238756
rect 221556 233980 221608 233986
rect 221556 233922 221608 233928
rect 223776 233034 223804 238750
rect 223764 233028 223816 233034
rect 223764 232970 223816 232976
rect 220084 231124 220136 231130
rect 220084 231066 220136 231072
rect 220176 231124 220228 231130
rect 220176 231066 220228 231072
rect 220096 178702 220124 231066
rect 221464 218816 221516 218822
rect 221464 218758 221516 218764
rect 221476 184414 221504 218758
rect 222844 200864 222896 200870
rect 222844 200806 222896 200812
rect 221464 184408 221516 184414
rect 221464 184350 221516 184356
rect 222856 181558 222884 200806
rect 222844 181552 222896 181558
rect 222844 181494 222896 181500
rect 224972 178770 225000 240094
rect 227686 239850 227714 240108
rect 229112 240094 229632 240122
rect 231872 240094 232208 240122
rect 227686 239822 227760 239850
rect 227732 206922 227760 239822
rect 229112 218822 229140 240094
rect 231872 227798 231900 240094
rect 234126 239850 234154 240108
rect 236072 240094 236408 240122
rect 234080 239822 234154 239850
rect 234080 235686 234108 239822
rect 236380 238474 236408 240094
rect 237392 240094 238004 240122
rect 240152 240094 240580 240122
rect 242268 240094 242512 240122
rect 244292 240094 244444 240122
rect 245672 240094 246376 240122
rect 248432 240094 248952 240122
rect 250548 240094 250884 240122
rect 252816 240094 253244 240122
rect 236368 238468 236420 238474
rect 236368 238410 236420 238416
rect 234068 235680 234120 235686
rect 234068 235622 234120 235628
rect 234080 233102 234108 235622
rect 234068 233096 234120 233102
rect 234068 233038 234120 233044
rect 231860 227792 231912 227798
rect 231860 227734 231912 227740
rect 233148 227792 233200 227798
rect 233148 227734 233200 227740
rect 229100 218816 229152 218822
rect 229100 218758 229152 218764
rect 229744 213444 229796 213450
rect 229744 213386 229796 213392
rect 227720 206916 227772 206922
rect 227720 206858 227772 206864
rect 229756 178838 229784 213386
rect 233160 200122 233188 227734
rect 236644 220312 236696 220318
rect 236644 220254 236696 220260
rect 233884 209092 233936 209098
rect 233884 209034 233936 209040
rect 233148 200116 233200 200122
rect 233148 200058 233200 200064
rect 232504 198212 232556 198218
rect 232504 198154 232556 198160
rect 232516 178945 232544 198154
rect 232502 178936 232558 178945
rect 232502 178871 232558 178880
rect 229744 178832 229796 178838
rect 229744 178774 229796 178780
rect 224960 178764 225012 178770
rect 224960 178706 225012 178712
rect 220084 178696 220136 178702
rect 220084 178638 220136 178644
rect 233896 176662 233924 209034
rect 236656 187202 236684 220254
rect 236736 195288 236788 195294
rect 236736 195230 236788 195236
rect 236644 187196 236696 187202
rect 236644 187138 236696 187144
rect 236748 180402 236776 195230
rect 236736 180396 236788 180402
rect 236736 180338 236788 180344
rect 237392 180334 237420 240094
rect 240152 238542 240180 240094
rect 240140 238536 240192 238542
rect 240140 238478 240192 238484
rect 240152 238338 240180 238478
rect 240140 238332 240192 238338
rect 240140 238274 240192 238280
rect 242268 237969 242296 240094
rect 242254 237960 242310 237969
rect 242254 237895 242310 237904
rect 242164 235272 242216 235278
rect 239402 235240 239458 235249
rect 242164 235214 242216 235220
rect 239402 235175 239458 235184
rect 239416 188630 239444 235175
rect 240784 221468 240836 221474
rect 240784 221410 240836 221416
rect 239496 209296 239548 209302
rect 239496 209238 239548 209244
rect 239404 188624 239456 188630
rect 239404 188566 239456 188572
rect 237380 180328 237432 180334
rect 237380 180270 237432 180276
rect 239508 177546 239536 209238
rect 239588 193996 239640 194002
rect 239588 193938 239640 193944
rect 239496 177540 239548 177546
rect 239496 177482 239548 177488
rect 239600 177410 239628 193938
rect 240796 178770 240824 221410
rect 242176 203862 242204 235214
rect 242268 227662 242296 237895
rect 243544 231260 243596 231266
rect 243544 231202 243596 231208
rect 242256 227656 242308 227662
rect 242256 227598 242308 227604
rect 242256 203924 242308 203930
rect 242256 203866 242308 203872
rect 242164 203856 242216 203862
rect 242164 203798 242216 203804
rect 242164 191208 242216 191214
rect 242164 191150 242216 191156
rect 242176 180470 242204 191150
rect 242164 180464 242216 180470
rect 242164 180406 242216 180412
rect 240784 178764 240836 178770
rect 240784 178706 240836 178712
rect 242268 177478 242296 203866
rect 243556 192778 243584 231202
rect 244292 229838 244320 240094
rect 244280 229832 244332 229838
rect 244280 229774 244332 229780
rect 245672 226370 245700 240094
rect 248432 231266 248460 240094
rect 250548 238678 250576 240094
rect 250536 238672 250588 238678
rect 250536 238614 250588 238620
rect 250548 235958 250576 238614
rect 253216 238406 253244 240094
rect 253952 240094 254748 240122
rect 257324 240094 257660 240122
rect 259256 240094 259408 240122
rect 261188 240094 261524 240122
rect 253204 238400 253256 238406
rect 253204 238342 253256 238348
rect 250536 235952 250588 235958
rect 250536 235894 250588 235900
rect 248420 231260 248472 231266
rect 248420 231202 248472 231208
rect 245660 226364 245712 226370
rect 245660 226306 245712 226312
rect 246948 226364 247000 226370
rect 246948 226306 247000 226312
rect 246304 202428 246356 202434
rect 246304 202370 246356 202376
rect 243544 192772 243596 192778
rect 243544 192714 243596 192720
rect 242348 185768 242400 185774
rect 242348 185710 242400 185716
rect 242256 177472 242308 177478
rect 242256 177414 242308 177420
rect 239588 177404 239640 177410
rect 239588 177346 239640 177352
rect 233884 176656 233936 176662
rect 233884 176598 233936 176604
rect 242360 176594 242388 185710
rect 245660 180192 245712 180198
rect 245660 180134 245712 180140
rect 245672 177585 245700 180134
rect 246316 178809 246344 202370
rect 246960 201482 246988 226306
rect 253216 224874 253244 238342
rect 253952 224913 253980 240094
rect 257632 238066 257660 240094
rect 257620 238060 257672 238066
rect 257620 238002 257672 238008
rect 259380 233209 259408 240094
rect 261496 236774 261524 240094
rect 263106 239850 263134 240108
rect 263060 239822 263134 239850
rect 265544 240094 265696 240122
rect 266372 240094 267628 240122
rect 269224 240094 269560 240122
rect 263060 239018 263088 239822
rect 263048 239012 263100 239018
rect 263048 238954 263100 238960
rect 262128 238060 262180 238066
rect 262128 238002 262180 238008
rect 261484 236768 261536 236774
rect 261484 236710 261536 236716
rect 259366 233200 259422 233209
rect 259366 233135 259422 233144
rect 262140 232529 262168 238002
rect 263060 235618 263088 238954
rect 264980 238672 265032 238678
rect 264980 238614 265032 238620
rect 264992 238513 265020 238614
rect 264978 238504 265034 238513
rect 264978 238439 265034 238448
rect 265544 237017 265572 240094
rect 265530 237008 265586 237017
rect 265530 236943 265586 236952
rect 265544 236065 265572 236943
rect 264058 236056 264114 236065
rect 264058 235991 264114 236000
rect 265530 236056 265586 236065
rect 265530 235991 265586 236000
rect 263048 235612 263100 235618
rect 263048 235554 263100 235560
rect 262126 232520 262182 232529
rect 262126 232455 262182 232464
rect 264072 231810 264100 235991
rect 264060 231804 264112 231810
rect 264060 231746 264112 231752
rect 266268 229832 266320 229838
rect 266268 229774 266320 229780
rect 261484 229764 261536 229770
rect 261484 229706 261536 229712
rect 253938 224904 253994 224913
rect 253204 224868 253256 224874
rect 253938 224839 253994 224848
rect 253204 224810 253256 224816
rect 249800 224324 249852 224330
rect 249800 224266 249852 224272
rect 247684 213376 247736 213382
rect 247684 213318 247736 213324
rect 246948 201476 247000 201482
rect 246948 201418 247000 201424
rect 246396 189916 246448 189922
rect 246396 189858 246448 189864
rect 246408 178906 246436 189858
rect 246396 178900 246448 178906
rect 246396 178842 246448 178848
rect 246948 178832 247000 178838
rect 246302 178800 246358 178809
rect 246948 178774 247000 178780
rect 246302 178735 246358 178744
rect 245658 177576 245714 177585
rect 245658 177511 245714 177520
rect 242348 176588 242400 176594
rect 242348 176530 242400 176536
rect 246960 175817 246988 178774
rect 247696 177954 247724 213318
rect 247776 205216 247828 205222
rect 247776 205158 247828 205164
rect 247684 177948 247736 177954
rect 247684 177890 247736 177896
rect 247788 175982 247816 205158
rect 247868 192704 247920 192710
rect 247868 192646 247920 192652
rect 247880 177857 247908 192646
rect 247960 188556 248012 188562
rect 247960 188498 248012 188504
rect 247972 178838 248000 188498
rect 249340 178900 249392 178906
rect 249340 178842 249392 178848
rect 247960 178832 248012 178838
rect 247960 178774 248012 178780
rect 249064 178832 249116 178838
rect 249064 178774 249116 178780
rect 247866 177848 247922 177857
rect 247866 177783 247922 177792
rect 247776 175976 247828 175982
rect 247776 175918 247828 175924
rect 246946 175808 247002 175817
rect 246946 175743 247002 175752
rect 249076 172553 249104 178774
rect 249248 177948 249300 177954
rect 249248 177890 249300 177896
rect 249156 176588 249208 176594
rect 249156 176530 249208 176536
rect 249062 172544 249118 172553
rect 249062 172479 249118 172488
rect 249168 171873 249196 176530
rect 249260 175273 249288 177890
rect 249246 175264 249302 175273
rect 249246 175199 249302 175208
rect 249154 171864 249210 171873
rect 249154 171799 249210 171808
rect 249352 171465 249380 178842
rect 249338 171456 249394 171465
rect 249338 171391 249394 171400
rect 249812 154465 249840 224266
rect 253940 221536 253992 221542
rect 253940 221478 253992 221484
rect 251180 220176 251232 220182
rect 251180 220118 251232 220124
rect 249892 183116 249944 183122
rect 249892 183058 249944 183064
rect 249798 154456 249854 154465
rect 249798 154391 249854 154400
rect 249904 149297 249932 183058
rect 250076 177540 250128 177546
rect 250076 177482 250128 177488
rect 249982 176080 250038 176089
rect 249982 176015 250038 176024
rect 249996 173777 250024 176015
rect 249982 173768 250038 173777
rect 249982 173703 250038 173712
rect 250088 170921 250116 177482
rect 250074 170912 250130 170921
rect 250074 170847 250130 170856
rect 251192 159633 251220 220118
rect 252560 215960 252612 215966
rect 252560 215902 252612 215908
rect 251272 205012 251324 205018
rect 251272 204954 251324 204960
rect 251178 159624 251234 159633
rect 251178 159559 251234 159568
rect 251180 154284 251232 154290
rect 251180 154226 251232 154232
rect 251192 153513 251220 154226
rect 251178 153504 251234 153513
rect 251178 153439 251234 153448
rect 250626 149696 250682 149705
rect 250626 149631 250682 149640
rect 249890 149288 249946 149297
rect 249890 149223 249946 149232
rect 250536 139460 250588 139466
rect 250536 139402 250588 139408
rect 250444 138032 250496 138038
rect 250444 137974 250496 137980
rect 249156 107908 249208 107914
rect 249156 107850 249208 107856
rect 249064 96688 249116 96694
rect 249064 96630 249116 96636
rect 242900 86284 242952 86290
rect 242900 86226 242952 86232
rect 238024 83564 238076 83570
rect 238024 83506 238076 83512
rect 216680 38004 216732 38010
rect 216680 37946 216732 37952
rect 215944 4140 215996 4146
rect 215944 4082 215996 4088
rect 214564 3596 214616 3602
rect 214564 3538 214616 3544
rect 238036 3534 238064 83506
rect 238760 82748 238812 82754
rect 238760 82690 238812 82696
rect 238772 16574 238800 82690
rect 241520 64320 241572 64326
rect 241520 64262 241572 64268
rect 240784 36712 240836 36718
rect 240784 36654 240836 36660
rect 238772 16546 239352 16574
rect 235816 3528 235868 3534
rect 235816 3470 235868 3476
rect 238024 3528 238076 3534
rect 238024 3470 238076 3476
rect 185584 3460 185636 3466
rect 185584 3402 185636 3408
rect 206284 3460 206336 3466
rect 206284 3402 206336 3408
rect 235828 480 235856 3470
rect 239324 480 239352 16546
rect 240796 15201 240824 36654
rect 241532 16574 241560 64262
rect 241532 16546 241744 16574
rect 240138 15192 240194 15201
rect 240138 15127 240194 15136
rect 240782 15192 240838 15201
rect 240782 15127 240838 15136
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 15127
rect 241716 480 241744 16546
rect 242912 3534 242940 86226
rect 245658 86184 245714 86193
rect 245658 86119 245714 86128
rect 245672 78674 245700 86119
rect 245660 78668 245712 78674
rect 245660 78610 245712 78616
rect 244924 51876 244976 51882
rect 244924 51818 244976 51824
rect 244936 19310 244964 51818
rect 244280 19304 244332 19310
rect 244280 19246 244332 19252
rect 244924 19304 244976 19310
rect 244924 19246 244976 19252
rect 244292 16574 244320 19246
rect 245672 16574 245700 78610
rect 247684 72480 247736 72486
rect 247684 72422 247736 72428
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 242992 3596 243044 3602
rect 242992 3538 243044 3544
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 243004 1850 243032 3538
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 242912 1822 243032 1850
rect 242912 480 242940 1822
rect 244108 480 244136 3470
rect 245212 480 245240 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247696 6914 247724 72422
rect 248420 45620 248472 45626
rect 248420 45562 248472 45568
rect 247604 6886 247724 6914
rect 247604 4146 247632 6886
rect 247592 4140 247644 4146
rect 247592 4082 247644 4088
rect 247604 480 247632 4082
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 45562
rect 249076 7614 249104 96630
rect 249168 68338 249196 107850
rect 249798 96656 249854 96665
rect 249798 96591 249854 96600
rect 249156 68332 249208 68338
rect 249156 68274 249208 68280
rect 249812 22098 249840 96591
rect 250456 24138 250484 137974
rect 250548 72554 250576 139402
rect 250640 137057 250668 149631
rect 251284 147937 251312 204954
rect 251364 192568 251416 192574
rect 251364 192510 251416 192516
rect 251376 161106 251404 192510
rect 251456 177336 251508 177342
rect 251456 177278 251508 177284
rect 251468 171134 251496 177278
rect 251468 171106 251680 171134
rect 251456 165232 251508 165238
rect 251456 165174 251508 165180
rect 251468 164393 251496 165174
rect 251454 164384 251510 164393
rect 251454 164319 251510 164328
rect 251376 161078 251588 161106
rect 251364 160880 251416 160886
rect 251364 160822 251416 160828
rect 251376 160585 251404 160822
rect 251362 160576 251418 160585
rect 251362 160511 251418 160520
rect 251560 156369 251588 161078
rect 251652 159225 251680 171106
rect 252468 170672 252520 170678
rect 252468 170614 252520 170620
rect 252480 170513 252508 170614
rect 252466 170504 252522 170513
rect 252466 170439 252522 170448
rect 252376 169584 252428 169590
rect 252376 169526 252428 169532
rect 252388 168609 252416 169526
rect 252468 169516 252520 169522
rect 252468 169458 252520 169464
rect 252480 169153 252508 169458
rect 252466 169144 252522 169153
rect 252466 169079 252522 169088
rect 252374 168600 252430 168609
rect 252374 168535 252430 168544
rect 252376 168360 252428 168366
rect 252376 168302 252428 168308
rect 252008 167748 252060 167754
rect 252008 167690 252060 167696
rect 252020 167249 252048 167690
rect 252388 167657 252416 168302
rect 252468 168292 252520 168298
rect 252468 168234 252520 168240
rect 252480 168201 252508 168234
rect 252466 168192 252522 168201
rect 252466 168127 252522 168136
rect 252374 167648 252430 167657
rect 252374 167583 252430 167592
rect 252006 167240 252062 167249
rect 252006 167175 252062 167184
rect 252376 167000 252428 167006
rect 252376 166942 252428 166948
rect 251916 166320 251968 166326
rect 251914 166288 251916 166297
rect 251968 166288 251970 166297
rect 251914 166223 251970 166232
rect 252388 165753 252416 166942
rect 252466 166696 252522 166705
rect 252466 166631 252522 166640
rect 252480 165918 252508 166631
rect 252468 165912 252520 165918
rect 252468 165854 252520 165860
rect 252374 165744 252430 165753
rect 252374 165679 252430 165688
rect 251916 165572 251968 165578
rect 251916 165514 251968 165520
rect 251928 164801 251956 165514
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 252480 164966 252508 165271
rect 252468 164960 252520 164966
rect 252468 164902 252520 164908
rect 251914 164792 251970 164801
rect 251914 164727 251970 164736
rect 252192 164212 252244 164218
rect 252192 164154 252244 164160
rect 251916 164144 251968 164150
rect 251916 164086 251968 164092
rect 251928 163441 251956 164086
rect 251914 163432 251970 163441
rect 251914 163367 251970 163376
rect 252204 163033 252232 164154
rect 252190 163024 252246 163033
rect 252190 162959 252246 162968
rect 252468 162852 252520 162858
rect 252468 162794 252520 162800
rect 252100 162784 252152 162790
rect 252100 162726 252152 162732
rect 252112 162489 252140 162726
rect 252098 162480 252154 162489
rect 252098 162415 252154 162424
rect 252480 162081 252508 162794
rect 252466 162072 252522 162081
rect 252466 162007 252522 162016
rect 252468 161560 252520 161566
rect 252466 161528 252468 161537
rect 252520 161528 252522 161537
rect 252466 161463 252522 161472
rect 252466 161120 252522 161129
rect 252466 161055 252522 161064
rect 252480 160750 252508 161055
rect 252468 160744 252520 160750
rect 252468 160686 252520 160692
rect 251916 160404 251968 160410
rect 251916 160346 251968 160352
rect 251928 160177 251956 160346
rect 251914 160168 251970 160177
rect 251914 160103 251970 160112
rect 251638 159216 251694 159225
rect 251638 159151 251694 159160
rect 252376 158704 252428 158710
rect 252376 158646 252428 158652
rect 252388 157865 252416 158646
rect 252468 158636 252520 158642
rect 252468 158578 252520 158584
rect 252480 158273 252508 158578
rect 252466 158264 252522 158273
rect 252466 158199 252522 158208
rect 252374 157856 252430 157865
rect 252374 157791 252430 157800
rect 252468 157344 252520 157350
rect 252468 157286 252520 157292
rect 252480 156913 252508 157286
rect 252466 156904 252522 156913
rect 252466 156839 252522 156848
rect 251546 156360 251602 156369
rect 251546 156295 251602 156304
rect 252466 155952 252522 155961
rect 252466 155887 252468 155896
rect 252520 155887 252522 155896
rect 252468 155858 252520 155864
rect 252376 155848 252428 155854
rect 252376 155790 252428 155796
rect 252388 155009 252416 155790
rect 252468 155780 252520 155786
rect 252468 155722 252520 155728
rect 252480 155417 252508 155722
rect 252466 155408 252522 155417
rect 252466 155343 252522 155352
rect 252374 155000 252430 155009
rect 252374 154935 252430 154944
rect 251732 154556 251784 154562
rect 251732 154498 251784 154504
rect 251744 154057 251772 154498
rect 251730 154048 251786 154057
rect 251730 153983 251786 153992
rect 252008 153196 252060 153202
rect 252008 153138 252060 153144
rect 252020 152153 252048 153138
rect 252468 153128 252520 153134
rect 252466 153096 252468 153105
rect 252520 153096 252522 153105
rect 252466 153031 252522 153040
rect 252006 152144 252062 152153
rect 252006 152079 252062 152088
rect 252466 151736 252522 151745
rect 252466 151671 252468 151680
rect 252520 151671 252522 151680
rect 252468 151642 252520 151648
rect 252376 151632 252428 151638
rect 252376 151574 252428 151580
rect 252388 150793 252416 151574
rect 252374 150784 252430 150793
rect 252374 150719 252430 150728
rect 251916 150408 251968 150414
rect 251916 150350 251968 150356
rect 251548 150340 251600 150346
rect 251548 150282 251600 150288
rect 251560 149841 251588 150282
rect 251928 150249 251956 150350
rect 251914 150240 251970 150249
rect 251914 150175 251970 150184
rect 251546 149832 251602 149841
rect 251546 149767 251602 149776
rect 252572 149138 252600 215902
rect 252744 207732 252796 207738
rect 252744 207674 252796 207680
rect 252652 206372 252704 206378
rect 252652 206314 252704 206320
rect 252664 151201 252692 206314
rect 252756 169561 252784 207674
rect 252836 202224 252888 202230
rect 252836 202166 252888 202172
rect 252742 169552 252798 169561
rect 252742 169487 252798 169496
rect 252848 165238 252876 202166
rect 252836 165232 252888 165238
rect 252836 165174 252888 165180
rect 253296 162920 253348 162926
rect 253296 162862 253348 162868
rect 252650 151192 252706 151201
rect 252650 151127 252706 151136
rect 252652 149796 252704 149802
rect 252652 149738 252704 149744
rect 252388 149110 252600 149138
rect 252388 148889 252416 149110
rect 252468 149048 252520 149054
rect 252468 148990 252520 148996
rect 252374 148880 252430 148889
rect 252374 148815 252430 148824
rect 252008 148368 252060 148374
rect 252480 148345 252508 148990
rect 252008 148310 252060 148316
rect 252466 148336 252522 148345
rect 251270 147928 251326 147937
rect 251270 147863 251326 147872
rect 251180 147008 251232 147014
rect 251178 146976 251180 146985
rect 251232 146976 251234 146985
rect 251178 146911 251234 146920
rect 251548 146940 251600 146946
rect 251548 146882 251600 146888
rect 251560 144673 251588 146882
rect 251732 146260 251784 146266
rect 251732 146202 251784 146208
rect 251546 144664 251602 144673
rect 251546 144599 251602 144608
rect 251744 143177 251772 146202
rect 251916 146192 251968 146198
rect 251916 146134 251968 146140
rect 251928 146033 251956 146134
rect 251914 146024 251970 146033
rect 251914 145959 251970 145968
rect 252020 145738 252048 148310
rect 252466 148271 252522 148280
rect 252376 147552 252428 147558
rect 252376 147494 252428 147500
rect 252466 147520 252522 147529
rect 252388 146577 252416 147494
rect 252466 147455 252468 147464
rect 252520 147455 252522 147464
rect 252468 147426 252520 147432
rect 252374 146568 252430 146577
rect 252374 146503 252430 146512
rect 252100 146124 252152 146130
rect 252100 146066 252152 146072
rect 251928 145710 252048 145738
rect 251730 143168 251786 143177
rect 251730 143103 251786 143112
rect 251824 142724 251876 142730
rect 251824 142666 251876 142672
rect 251086 142624 251142 142633
rect 251086 142559 251142 142568
rect 250626 137048 250682 137057
rect 250626 136983 250682 136992
rect 251100 109177 251128 142559
rect 251732 142112 251784 142118
rect 251732 142054 251784 142060
rect 251744 141409 251772 142054
rect 251730 141400 251786 141409
rect 251730 141335 251786 141344
rect 251732 139528 251784 139534
rect 251730 139496 251732 139505
rect 251784 139496 251786 139505
rect 251730 139431 251786 139440
rect 251732 139392 251784 139398
rect 251732 139334 251784 139340
rect 251744 138553 251772 139334
rect 251730 138544 251786 138553
rect 251730 138479 251786 138488
rect 251362 138000 251418 138009
rect 251362 137935 251418 137944
rect 251376 137902 251404 137935
rect 251364 137896 251416 137902
rect 251364 137838 251416 137844
rect 251732 136536 251784 136542
rect 251732 136478 251784 136484
rect 251744 135697 251772 136478
rect 251730 135688 251786 135697
rect 251730 135623 251786 135632
rect 251456 135244 251508 135250
rect 251456 135186 251508 135192
rect 251468 134745 251496 135186
rect 251454 134736 251510 134745
rect 251454 134671 251510 134680
rect 251364 133884 251416 133890
rect 251364 133826 251416 133832
rect 251376 133793 251404 133826
rect 251362 133784 251418 133793
rect 251362 133719 251418 133728
rect 251548 132388 251600 132394
rect 251548 132330 251600 132336
rect 251560 131889 251588 132330
rect 251546 131880 251602 131889
rect 251546 131815 251602 131824
rect 251456 129668 251508 129674
rect 251456 129610 251508 129616
rect 251468 129169 251496 129610
rect 251454 129160 251510 129169
rect 251454 129095 251510 129104
rect 251640 128308 251692 128314
rect 251640 128250 251692 128256
rect 251652 127673 251680 128250
rect 251638 127664 251694 127673
rect 251638 127599 251694 127608
rect 251364 126268 251416 126274
rect 251364 126210 251416 126216
rect 251376 124409 251404 126210
rect 251362 124400 251418 124409
rect 251362 124335 251418 124344
rect 251180 123548 251232 123554
rect 251180 123490 251232 123496
rect 251192 123049 251220 123490
rect 251178 123040 251234 123049
rect 251178 122975 251234 122984
rect 251836 122834 251864 142666
rect 251928 127265 251956 145710
rect 252008 145648 252060 145654
rect 252008 145590 252060 145596
rect 252020 142154 252048 145590
rect 252112 145081 252140 146066
rect 252466 145616 252522 145625
rect 252664 145602 252692 149738
rect 252522 145574 252692 145602
rect 252466 145551 252522 145560
rect 252098 145072 252154 145081
rect 252098 145007 252154 145016
rect 252192 144900 252244 144906
rect 252192 144842 252244 144848
rect 252204 143721 252232 144842
rect 252466 144120 252522 144129
rect 252466 144055 252468 144064
rect 252520 144055 252522 144064
rect 252650 144120 252706 144129
rect 252650 144055 252706 144064
rect 252468 144026 252520 144032
rect 252190 143712 252246 143721
rect 252190 143647 252246 143656
rect 252468 143540 252520 143546
rect 252468 143482 252520 143488
rect 252480 142769 252508 143482
rect 252466 142760 252522 142769
rect 252466 142695 252522 142704
rect 252664 142154 252692 144055
rect 252020 142126 252140 142154
rect 252008 131844 252060 131850
rect 252008 131786 252060 131792
rect 251914 127256 251970 127265
rect 251914 127191 251970 127200
rect 251916 125384 251968 125390
rect 251914 125352 251916 125361
rect 251968 125352 251970 125361
rect 251914 125287 251970 125296
rect 252020 122834 252048 131786
rect 252112 131481 252140 142126
rect 252572 142126 252692 142154
rect 252376 141432 252428 141438
rect 252376 141374 252428 141380
rect 252388 135289 252416 141374
rect 252468 139324 252520 139330
rect 252468 139266 252520 139272
rect 252480 138961 252508 139266
rect 252466 138952 252522 138961
rect 252466 138887 252522 138896
rect 252468 137964 252520 137970
rect 252468 137906 252520 137912
rect 252480 137601 252508 137906
rect 252466 137592 252522 137601
rect 252466 137527 252522 137536
rect 252468 136604 252520 136610
rect 252468 136546 252520 136552
rect 252480 136241 252508 136546
rect 252466 136232 252522 136241
rect 252466 136167 252522 136176
rect 252374 135280 252430 135289
rect 252374 135215 252430 135224
rect 252468 135176 252520 135182
rect 252468 135118 252520 135124
rect 252480 134337 252508 135118
rect 252466 134328 252522 134337
rect 252466 134263 252522 134272
rect 252376 133816 252428 133822
rect 252376 133758 252428 133764
rect 252388 133385 252416 133758
rect 252468 133748 252520 133754
rect 252468 133690 252520 133696
rect 252374 133376 252430 133385
rect 252374 133311 252430 133320
rect 252480 132841 252508 133690
rect 252466 132832 252522 132841
rect 252466 132767 252522 132776
rect 252468 132456 252520 132462
rect 252466 132424 252468 132433
rect 252520 132424 252522 132433
rect 252466 132359 252522 132368
rect 252098 131472 252154 131481
rect 252098 131407 252154 131416
rect 252376 131096 252428 131102
rect 252376 131038 252428 131044
rect 252388 130121 252416 131038
rect 252468 131028 252520 131034
rect 252468 130970 252520 130976
rect 252480 130937 252508 130970
rect 252466 130928 252522 130937
rect 252466 130863 252522 130872
rect 252468 130552 252520 130558
rect 252466 130520 252468 130529
rect 252520 130520 252522 130529
rect 252466 130455 252522 130464
rect 252374 130112 252430 130121
rect 252374 130047 252430 130056
rect 252468 129736 252520 129742
rect 252468 129678 252520 129684
rect 252376 129600 252428 129606
rect 252480 129577 252508 129678
rect 252376 129542 252428 129548
rect 252466 129568 252522 129577
rect 252388 128625 252416 129542
rect 252466 129503 252522 129512
rect 252374 128616 252430 128625
rect 252374 128551 252430 128560
rect 252468 128240 252520 128246
rect 252466 128208 252468 128217
rect 252520 128208 252522 128217
rect 252466 128143 252522 128152
rect 252192 127492 252244 127498
rect 252192 127434 252244 127440
rect 252100 126880 252152 126886
rect 252100 126822 252152 126828
rect 252112 125769 252140 126822
rect 252098 125760 252154 125769
rect 252098 125695 252154 125704
rect 252204 122834 252232 127434
rect 252468 126948 252520 126954
rect 252468 126890 252520 126896
rect 252480 126721 252508 126890
rect 252466 126712 252522 126721
rect 252466 126647 252522 126656
rect 252468 125044 252520 125050
rect 252468 124986 252520 124992
rect 252284 124908 252336 124914
rect 252284 124850 252336 124856
rect 251744 122806 251864 122834
rect 251928 122806 252048 122834
rect 252112 122806 252232 122834
rect 251364 122528 251416 122534
rect 251364 122470 251416 122476
rect 251376 122097 251404 122470
rect 251362 122088 251418 122097
rect 251362 122023 251418 122032
rect 251364 120012 251416 120018
rect 251364 119954 251416 119960
rect 251376 119649 251404 119954
rect 251362 119640 251418 119649
rect 251362 119575 251418 119584
rect 251744 117337 251772 122806
rect 251824 121372 251876 121378
rect 251824 121314 251876 121320
rect 251836 120601 251864 121314
rect 251822 120592 251878 120601
rect 251822 120527 251878 120536
rect 251824 118652 251876 118658
rect 251824 118594 251876 118600
rect 251836 117881 251864 118594
rect 251822 117872 251878 117881
rect 251822 117807 251878 117816
rect 251730 117328 251786 117337
rect 251364 117292 251416 117298
rect 251730 117263 251786 117272
rect 251364 117234 251416 117240
rect 251376 116929 251404 117234
rect 251362 116920 251418 116929
rect 251362 116855 251418 116864
rect 251928 115954 251956 122806
rect 252008 122732 252060 122738
rect 252008 122674 252060 122680
rect 252020 121553 252048 122674
rect 252006 121544 252062 121553
rect 252006 121479 252062 121488
rect 252008 116612 252060 116618
rect 252008 116554 252060 116560
rect 251744 115926 251956 115954
rect 251364 114504 251416 114510
rect 251744 114481 251772 115926
rect 251916 115864 251968 115870
rect 251916 115806 251968 115812
rect 251824 115252 251876 115258
rect 251824 115194 251876 115200
rect 251364 114446 251416 114452
rect 251730 114472 251786 114481
rect 251376 113529 251404 114446
rect 251730 114407 251786 114416
rect 251640 114232 251692 114238
rect 251640 114174 251692 114180
rect 251652 114073 251680 114174
rect 251638 114064 251694 114073
rect 251638 113999 251694 114008
rect 251362 113520 251418 113529
rect 251362 113455 251418 113464
rect 251836 113174 251864 115194
rect 251928 115025 251956 115806
rect 251914 115016 251970 115025
rect 251914 114951 251970 114960
rect 251744 113146 251864 113174
rect 251640 112260 251692 112266
rect 251640 112202 251692 112208
rect 251652 112169 251680 112202
rect 251638 112160 251694 112169
rect 251638 112095 251694 112104
rect 251086 109168 251142 109177
rect 251086 109103 251142 109112
rect 251364 106140 251416 106146
rect 251364 106082 251416 106088
rect 251376 105097 251404 106082
rect 251362 105088 251418 105097
rect 251362 105023 251418 105032
rect 251744 103737 251772 113146
rect 251824 111308 251876 111314
rect 251824 111250 251876 111256
rect 251836 107001 251864 111250
rect 252020 111217 252048 116554
rect 252112 111761 252140 122806
rect 252296 120193 252324 124850
rect 252480 124817 252508 124986
rect 252466 124808 252522 124817
rect 252466 124743 252522 124752
rect 252376 124160 252428 124166
rect 252376 124102 252428 124108
rect 252388 123457 252416 124102
rect 252468 124092 252520 124098
rect 252468 124034 252520 124040
rect 252480 124001 252508 124034
rect 252466 123992 252522 124001
rect 252466 123927 252522 123936
rect 252374 123448 252430 123457
rect 252374 123383 252430 123392
rect 252468 122800 252520 122806
rect 252468 122742 252520 122748
rect 252480 122505 252508 122742
rect 252466 122496 252522 122505
rect 252466 122431 252522 122440
rect 252468 121440 252520 121446
rect 252468 121382 252520 121388
rect 252480 121145 252508 121382
rect 252466 121136 252522 121145
rect 252466 121071 252522 121080
rect 252376 120284 252428 120290
rect 252376 120226 252428 120232
rect 252282 120184 252338 120193
rect 252282 120119 252338 120128
rect 252284 119332 252336 119338
rect 252284 119274 252336 119280
rect 252296 118833 252324 119274
rect 252282 118824 252338 118833
rect 252282 118759 252338 118768
rect 252388 116385 252416 120226
rect 252468 120080 252520 120086
rect 252468 120022 252520 120028
rect 252480 119241 252508 120022
rect 252466 119232 252522 119241
rect 252466 119167 252522 119176
rect 252468 118584 252520 118590
rect 252468 118526 252520 118532
rect 252480 118289 252508 118526
rect 252466 118280 252522 118289
rect 252466 118215 252522 118224
rect 252468 117224 252520 117230
rect 252468 117166 252520 117172
rect 252374 116376 252430 116385
rect 252374 116311 252430 116320
rect 252480 115977 252508 117166
rect 252466 115968 252522 115977
rect 252284 115932 252336 115938
rect 252466 115903 252522 115912
rect 252284 115874 252336 115880
rect 252296 115433 252324 115874
rect 252282 115424 252338 115433
rect 252282 115359 252338 115368
rect 252468 113824 252520 113830
rect 252468 113766 252520 113772
rect 252480 113121 252508 113766
rect 252466 113112 252522 113121
rect 252466 113047 252522 113056
rect 252468 112872 252520 112878
rect 252468 112814 252520 112820
rect 252480 112713 252508 112814
rect 252466 112704 252522 112713
rect 252466 112639 252522 112648
rect 252192 112532 252244 112538
rect 252192 112474 252244 112480
rect 252098 111752 252154 111761
rect 252098 111687 252154 111696
rect 252006 111208 252062 111217
rect 252006 111143 252062 111152
rect 251916 110424 251968 110430
rect 251916 110366 251968 110372
rect 251928 110265 251956 110366
rect 252100 110288 252152 110294
rect 251914 110256 251970 110265
rect 252100 110230 252152 110236
rect 251914 110191 251970 110200
rect 252112 109313 252140 110230
rect 252098 109304 252154 109313
rect 252098 109239 252154 109248
rect 252100 107636 252152 107642
rect 252100 107578 252152 107584
rect 251822 106992 251878 107001
rect 251822 106927 251878 106936
rect 252008 106956 252060 106962
rect 252008 106898 252060 106904
rect 251916 106208 251968 106214
rect 251916 106150 251968 106156
rect 251928 106049 251956 106150
rect 251914 106040 251970 106049
rect 251914 105975 251970 105984
rect 251916 104848 251968 104854
rect 251916 104790 251968 104796
rect 251928 104689 251956 104790
rect 251914 104680 251970 104689
rect 251914 104615 251970 104624
rect 251730 103728 251786 103737
rect 251730 103663 251786 103672
rect 252020 103514 252048 106898
rect 252112 106593 252140 107578
rect 252204 107545 252232 112474
rect 252284 111104 252336 111110
rect 252284 111046 252336 111052
rect 252296 107953 252324 111046
rect 252468 110356 252520 110362
rect 252468 110298 252520 110304
rect 252480 109857 252508 110298
rect 252466 109848 252522 109857
rect 252466 109783 252522 109792
rect 252376 108996 252428 109002
rect 252376 108938 252428 108944
rect 252388 108361 252416 108938
rect 252468 108928 252520 108934
rect 252466 108896 252468 108905
rect 252520 108896 252522 108905
rect 252466 108831 252522 108840
rect 252374 108352 252430 108361
rect 252374 108287 252430 108296
rect 252282 107944 252338 107953
rect 252282 107879 252338 107888
rect 252190 107536 252246 107545
rect 252190 107471 252246 107480
rect 252098 106584 252154 106593
rect 252098 106519 252154 106528
rect 252468 106276 252520 106282
rect 252468 106218 252520 106224
rect 252480 105641 252508 106218
rect 252466 105632 252522 105641
rect 252466 105567 252522 105576
rect 252468 104780 252520 104786
rect 252468 104722 252520 104728
rect 252284 104168 252336 104174
rect 252480 104145 252508 104722
rect 252284 104110 252336 104116
rect 252466 104136 252522 104145
rect 251928 103486 252048 103514
rect 251732 100700 251784 100706
rect 251732 100642 251784 100648
rect 251744 99929 251772 100642
rect 251730 99920 251786 99929
rect 251730 99855 251786 99864
rect 251548 99340 251600 99346
rect 251548 99282 251600 99288
rect 251180 99136 251232 99142
rect 251180 99078 251232 99084
rect 251192 98977 251220 99078
rect 251178 98968 251234 98977
rect 251178 98903 251234 98912
rect 251560 98025 251588 99282
rect 251824 99204 251876 99210
rect 251824 99146 251876 99152
rect 251836 98569 251864 99146
rect 251822 98560 251878 98569
rect 251822 98495 251878 98504
rect 251546 98016 251602 98025
rect 251546 97951 251602 97960
rect 251928 97073 251956 103486
rect 252008 103420 252060 103426
rect 252008 103362 252060 103368
rect 252020 103193 252048 103362
rect 252006 103184 252062 103193
rect 252006 103119 252062 103128
rect 252296 101833 252324 104110
rect 252466 104071 252522 104080
rect 252468 103488 252520 103494
rect 252468 103430 252520 103436
rect 252376 103012 252428 103018
rect 252376 102954 252428 102960
rect 252388 102785 252416 102954
rect 252374 102776 252430 102785
rect 252374 102711 252430 102720
rect 252480 102241 252508 103430
rect 252466 102232 252522 102241
rect 252466 102167 252522 102176
rect 252468 102128 252520 102134
rect 252468 102070 252520 102076
rect 252282 101824 252338 101833
rect 252282 101759 252338 101768
rect 252100 101448 252152 101454
rect 252480 101425 252508 102070
rect 252100 101390 252152 101396
rect 252466 101416 252522 101425
rect 252008 100904 252060 100910
rect 252006 100872 252008 100881
rect 252060 100872 252062 100881
rect 252006 100807 252062 100816
rect 251178 97064 251234 97073
rect 251178 96999 251234 97008
rect 251914 97064 251970 97073
rect 251914 96999 251970 97008
rect 250536 72548 250588 72554
rect 250536 72490 250588 72496
rect 251192 55214 251220 96999
rect 251916 96756 251968 96762
rect 251916 96698 251968 96704
rect 251270 96248 251326 96257
rect 251270 96183 251326 96192
rect 251284 83570 251312 96183
rect 251272 83564 251324 83570
rect 251272 83506 251324 83512
rect 251180 55208 251232 55214
rect 251180 55150 251232 55156
rect 251180 38004 251232 38010
rect 251180 37946 251232 37952
rect 250444 24132 250496 24138
rect 250444 24074 250496 24080
rect 249800 22092 249852 22098
rect 249800 22034 249852 22040
rect 249984 13252 250036 13258
rect 249984 13194 250036 13200
rect 249064 7608 249116 7614
rect 249064 7550 249116 7556
rect 249996 480 250024 13194
rect 251192 480 251220 37946
rect 251928 31074 251956 96698
rect 252112 96665 252140 101390
rect 252466 101351 252522 101360
rect 252468 100632 252520 100638
rect 252468 100574 252520 100580
rect 252376 100564 252428 100570
rect 252376 100506 252428 100512
rect 252388 99521 252416 100506
rect 252480 100473 252508 100574
rect 252466 100464 252522 100473
rect 252466 100399 252522 100408
rect 252374 99512 252430 99521
rect 252374 99447 252430 99456
rect 252192 97640 252244 97646
rect 252190 97608 252192 97617
rect 252244 97608 252246 97617
rect 252190 97543 252246 97552
rect 252098 96656 252154 96665
rect 252098 96591 252154 96600
rect 251916 31068 251968 31074
rect 251916 31010 251968 31016
rect 252572 6914 252600 142126
rect 253204 138100 253256 138106
rect 253204 138042 253256 138048
rect 253216 10334 253244 138042
rect 253308 123554 253336 162862
rect 253952 147014 253980 221478
rect 257344 206440 257396 206446
rect 257344 206382 257396 206388
rect 254124 203720 254176 203726
rect 254124 203662 254176 203668
rect 254032 196648 254084 196654
rect 254032 196590 254084 196596
rect 254044 154290 254072 196590
rect 254136 160886 254164 203662
rect 255596 200932 255648 200938
rect 255596 200874 255648 200880
rect 255412 199436 255464 199442
rect 255412 199378 255464 199384
rect 254584 161492 254636 161498
rect 254584 161434 254636 161440
rect 254124 160880 254176 160886
rect 254124 160822 254176 160828
rect 254032 154284 254084 154290
rect 254032 154226 254084 154232
rect 253940 147008 253992 147014
rect 253940 146950 253992 146956
rect 253388 145580 253440 145586
rect 253388 145522 253440 145528
rect 253296 123548 253348 123554
rect 253296 123490 253348 123496
rect 253296 110492 253348 110498
rect 253296 110434 253348 110440
rect 253308 14550 253336 110434
rect 253400 99142 253428 145522
rect 254596 122534 254624 161434
rect 254768 153876 254820 153882
rect 254768 153818 254820 153824
rect 254676 146328 254728 146334
rect 254676 146270 254728 146276
rect 254584 122528 254636 122534
rect 254584 122470 254636 122476
rect 254584 117564 254636 117570
rect 254584 117506 254636 117512
rect 253388 99136 253440 99142
rect 253388 99078 253440 99084
rect 253296 14544 253348 14550
rect 253296 14486 253348 14492
rect 253204 10328 253256 10334
rect 253204 10270 253256 10276
rect 252572 6886 253520 6914
rect 252374 3496 252430 3505
rect 252374 3431 252430 3440
rect 252388 480 252416 3431
rect 253492 480 253520 6886
rect 254596 4826 254624 117506
rect 254688 106146 254716 146270
rect 254780 114238 254808 153818
rect 255424 150346 255452 199378
rect 255504 175976 255556 175982
rect 255504 175918 255556 175924
rect 255516 160410 255544 175918
rect 255504 160404 255556 160410
rect 255504 160346 255556 160352
rect 255412 150340 255464 150346
rect 255412 150282 255464 150288
rect 254860 149728 254912 149734
rect 254860 149670 254912 149676
rect 254768 114232 254820 114238
rect 254768 114174 254820 114180
rect 254872 112266 254900 149670
rect 255608 139534 255636 200874
rect 256976 188692 257028 188698
rect 256976 188634 257028 188640
rect 256884 178696 256936 178702
rect 256884 178638 256936 178644
rect 256792 177404 256844 177410
rect 256792 177346 256844 177352
rect 256804 166326 256832 177346
rect 256896 167754 256924 178638
rect 256988 170678 257016 188634
rect 257356 180198 257384 206382
rect 259552 205080 259604 205086
rect 259552 205022 259604 205028
rect 258172 192636 258224 192642
rect 258172 192578 258224 192584
rect 258080 188488 258132 188494
rect 258080 188430 258132 188436
rect 257344 180192 257396 180198
rect 257344 180134 257396 180140
rect 256976 170672 257028 170678
rect 256976 170614 257028 170620
rect 257528 169788 257580 169794
rect 257528 169730 257580 169736
rect 256884 167748 256936 167754
rect 256884 167690 256936 167696
rect 256792 166320 256844 166326
rect 256792 166262 256844 166268
rect 257344 157412 257396 157418
rect 257344 157354 257396 157360
rect 256148 150476 256200 150482
rect 256148 150418 256200 150424
rect 255964 142180 256016 142186
rect 255964 142122 256016 142128
rect 255596 139528 255648 139534
rect 255596 139470 255648 139476
rect 254860 112260 254912 112266
rect 254860 112202 254912 112208
rect 254676 106140 254728 106146
rect 254676 106082 254728 106088
rect 255976 100910 256004 142122
rect 256056 139528 256108 139534
rect 256056 139470 256108 139476
rect 255964 100904 256016 100910
rect 255964 100846 256016 100852
rect 256068 97646 256096 139470
rect 256160 110294 256188 150418
rect 257356 142730 257384 157354
rect 257436 152516 257488 152522
rect 257436 152458 257488 152464
rect 257344 142724 257396 142730
rect 257344 142666 257396 142672
rect 256240 137284 256292 137290
rect 256240 137226 256292 137232
rect 256252 125390 256280 137226
rect 257344 130008 257396 130014
rect 257344 129950 257396 129956
rect 256240 125384 256292 125390
rect 256240 125326 256292 125332
rect 256148 110288 256200 110294
rect 256148 110230 256200 110236
rect 256056 97640 256108 97646
rect 256056 97582 256108 97588
rect 255964 96824 256016 96830
rect 255964 96766 256016 96772
rect 255320 56024 255372 56030
rect 255320 55966 255372 55972
rect 254676 35352 254728 35358
rect 254676 35294 254728 35300
rect 254688 34542 254716 35294
rect 254676 34536 254728 34542
rect 254676 34478 254728 34484
rect 254584 4820 254636 4826
rect 254584 4762 254636 4768
rect 254688 480 254716 34478
rect 255332 16574 255360 55966
rect 255976 36650 256004 96766
rect 256056 39432 256108 39438
rect 256056 39374 256108 39380
rect 255964 36644 256016 36650
rect 255964 36586 256016 36592
rect 256068 34542 256096 39374
rect 256056 34536 256108 34542
rect 256056 34478 256108 34484
rect 255332 16546 255912 16574
rect 255884 480 255912 16546
rect 257356 15978 257384 129950
rect 257448 112878 257476 152458
rect 257540 130558 257568 169730
rect 257620 165640 257672 165646
rect 257620 165582 257672 165588
rect 257632 152969 257660 165582
rect 257618 152960 257674 152969
rect 257618 152895 257674 152904
rect 257712 151972 257764 151978
rect 257712 151914 257764 151920
rect 257620 140820 257672 140826
rect 257620 140762 257672 140768
rect 257528 130552 257580 130558
rect 257528 130494 257580 130500
rect 257436 112872 257488 112878
rect 257436 112814 257488 112820
rect 257528 112464 257580 112470
rect 257528 112406 257580 112412
rect 257540 103018 257568 112406
rect 257528 103012 257580 103018
rect 257528 102954 257580 102960
rect 257436 102196 257488 102202
rect 257436 102138 257488 102144
rect 257448 40730 257476 102138
rect 257528 100972 257580 100978
rect 257528 100914 257580 100920
rect 257540 46306 257568 100914
rect 257632 99346 257660 140762
rect 257724 127498 257752 151914
rect 258092 144090 258120 188430
rect 258184 169522 258212 192578
rect 259460 189848 259512 189854
rect 259460 189790 259512 189796
rect 258356 180260 258408 180266
rect 258356 180202 258408 180208
rect 258264 177472 258316 177478
rect 258264 177414 258316 177420
rect 258172 169516 258224 169522
rect 258172 169458 258224 169464
rect 258276 160750 258304 177414
rect 258368 164966 258396 180202
rect 258356 164960 258408 164966
rect 258356 164902 258408 164908
rect 258908 164280 258960 164286
rect 258908 164222 258960 164228
rect 258264 160744 258316 160750
rect 258264 160686 258316 160692
rect 258816 155984 258868 155990
rect 258816 155926 258868 155932
rect 258080 144084 258132 144090
rect 258080 144026 258132 144032
rect 257712 127492 257764 127498
rect 257712 127434 257764 127440
rect 258724 124228 258776 124234
rect 258724 124170 258776 124176
rect 257620 99340 257672 99346
rect 257620 99282 257672 99288
rect 257528 46300 257580 46306
rect 257528 46242 257580 46248
rect 257436 40724 257488 40730
rect 257436 40666 257488 40672
rect 257344 15972 257396 15978
rect 257344 15914 257396 15920
rect 258736 13122 258764 124170
rect 258828 117230 258856 155926
rect 258920 125050 258948 164222
rect 259000 156052 259052 156058
rect 259000 155994 259052 156000
rect 258908 125044 258960 125050
rect 258908 124986 258960 124992
rect 259012 120290 259040 155994
rect 259472 142118 259500 189790
rect 259564 161566 259592 205022
rect 261024 198076 261076 198082
rect 261024 198018 261076 198024
rect 260840 191140 260892 191146
rect 260840 191082 260892 191088
rect 259644 184340 259696 184346
rect 259644 184282 259696 184288
rect 259552 161560 259604 161566
rect 259552 161502 259604 161508
rect 259656 146266 259684 184282
rect 259736 180464 259788 180470
rect 259736 180406 259788 180412
rect 259748 165918 259776 180406
rect 259736 165912 259788 165918
rect 259736 165854 259788 165860
rect 260288 158772 260340 158778
rect 260288 158714 260340 158720
rect 259644 146260 259696 146266
rect 259644 146202 259696 146208
rect 259460 142112 259512 142118
rect 259460 142054 259512 142060
rect 260196 127016 260248 127022
rect 260196 126958 260248 126964
rect 260104 122868 260156 122874
rect 260104 122810 260156 122816
rect 259000 120284 259052 120290
rect 259000 120226 259052 120232
rect 258816 117224 258868 117230
rect 258816 117166 258868 117172
rect 258816 109064 258868 109070
rect 258816 109006 258868 109012
rect 258828 17338 258856 109006
rect 259460 40724 259512 40730
rect 259460 40666 259512 40672
rect 258816 17332 258868 17338
rect 258816 17274 258868 17280
rect 258724 13116 258776 13122
rect 258724 13058 258776 13064
rect 256700 11892 256752 11898
rect 256700 11834 256752 11840
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 11834
rect 258262 3496 258318 3505
rect 258262 3431 258318 3440
rect 258276 480 258304 3431
rect 259472 480 259500 40666
rect 260116 29646 260144 122810
rect 260208 55894 260236 126958
rect 260300 119338 260328 158714
rect 260380 147688 260432 147694
rect 260380 147630 260432 147636
rect 260288 119332 260340 119338
rect 260288 119274 260340 119280
rect 260392 111314 260420 147630
rect 260852 139330 260880 191082
rect 260932 190052 260984 190058
rect 260932 189994 260984 190000
rect 260944 143546 260972 189994
rect 261036 167006 261064 198018
rect 261496 189854 261524 229706
rect 264244 222896 264296 222902
rect 264244 222838 264296 222844
rect 263600 205148 263652 205154
rect 263600 205090 263652 205096
rect 262312 194132 262364 194138
rect 262312 194074 262364 194080
rect 261484 189848 261536 189854
rect 261484 189790 261536 189796
rect 261116 184408 261168 184414
rect 261116 184350 261168 184356
rect 261024 167000 261076 167006
rect 261024 166942 261076 166948
rect 261128 162790 261156 184350
rect 262220 178764 262272 178770
rect 262220 178706 262272 178712
rect 261208 176656 261260 176662
rect 261206 176624 261208 176633
rect 261260 176624 261262 176633
rect 261206 176559 261262 176568
rect 261116 162784 261168 162790
rect 261116 162726 261168 162732
rect 261576 160132 261628 160138
rect 261576 160074 261628 160080
rect 260932 143540 260984 143546
rect 260932 143482 260984 143488
rect 260840 139324 260892 139330
rect 260840 139266 260892 139272
rect 261588 121378 261616 160074
rect 261668 155236 261720 155242
rect 261668 155178 261720 155184
rect 261576 121372 261628 121378
rect 261576 121314 261628 121320
rect 261484 120148 261536 120154
rect 261484 120090 261536 120096
rect 260380 111308 260432 111314
rect 260380 111250 260432 111256
rect 260196 55888 260248 55894
rect 260196 55830 260248 55836
rect 260104 29640 260156 29646
rect 260104 29582 260156 29588
rect 260840 18692 260892 18698
rect 260840 18634 260892 18640
rect 259552 17332 259604 17338
rect 259552 17274 259604 17280
rect 259564 16574 259592 17274
rect 260852 16574 260880 18634
rect 259564 16546 260696 16574
rect 260852 16546 261432 16574
rect 260668 480 260696 16546
rect 261404 3482 261432 16546
rect 261496 4894 261524 120090
rect 261680 117298 261708 155178
rect 262232 149802 262260 178706
rect 262324 168298 262352 194074
rect 262404 180396 262456 180402
rect 262404 180338 262456 180344
rect 262312 168292 262364 168298
rect 262312 168234 262364 168240
rect 262416 162858 262444 180338
rect 263048 162988 263100 162994
rect 263048 162930 263100 162936
rect 262404 162852 262456 162858
rect 262404 162794 262456 162800
rect 262864 157480 262916 157486
rect 262864 157422 262916 157428
rect 262220 149796 262272 149802
rect 262220 149738 262272 149744
rect 262876 118590 262904 157422
rect 262956 154624 263008 154630
rect 262956 154566 263008 154572
rect 262864 118584 262916 118590
rect 262864 118526 262916 118532
rect 261668 117292 261720 117298
rect 261668 117234 261720 117240
rect 262864 116000 262916 116006
rect 262864 115942 262916 115948
rect 262128 54596 262180 54602
rect 262128 54538 262180 54544
rect 262140 22001 262168 54538
rect 262876 42090 262904 115942
rect 262968 115870 262996 154566
rect 263060 124098 263088 162930
rect 263612 146946 263640 205090
rect 263692 196716 263744 196722
rect 263692 196658 263744 196664
rect 263704 168366 263732 196658
rect 264256 195294 264284 222838
rect 264980 210520 265032 210526
rect 264980 210462 265032 210468
rect 264244 195288 264296 195294
rect 264244 195230 264296 195236
rect 263784 189780 263836 189786
rect 263784 189722 263836 189728
rect 263796 169590 263824 189722
rect 264244 173936 264296 173942
rect 264244 173878 264296 173884
rect 263784 169584 263836 169590
rect 263784 169526 263836 169532
rect 263692 168360 263744 168366
rect 263692 168302 263744 168308
rect 263600 146940 263652 146946
rect 263600 146882 263652 146888
rect 264256 141438 264284 173878
rect 264336 167068 264388 167074
rect 264336 167010 264388 167016
rect 264244 141432 264296 141438
rect 264244 141374 264296 141380
rect 264348 128246 264376 167010
rect 264612 161560 264664 161566
rect 264612 161502 264664 161508
rect 264520 144220 264572 144226
rect 264520 144162 264572 144168
rect 264428 131164 264480 131170
rect 264428 131106 264480 131112
rect 264336 128240 264388 128246
rect 264336 128182 264388 128188
rect 264244 127084 264296 127090
rect 264244 127026 264296 127032
rect 263048 124092 263100 124098
rect 263048 124034 263100 124040
rect 262956 115864 263008 115870
rect 262956 115806 263008 115812
rect 263048 110560 263100 110566
rect 263048 110502 263100 110508
rect 262956 103556 263008 103562
rect 262956 103498 263008 103504
rect 262968 50454 262996 103498
rect 263060 65618 263088 110502
rect 263048 65612 263100 65618
rect 263048 65554 263100 65560
rect 262956 50448 263008 50454
rect 262956 50390 263008 50396
rect 262864 42084 262916 42090
rect 262864 42026 262916 42032
rect 262126 21992 262182 22001
rect 262126 21927 262182 21936
rect 262140 21570 262168 21927
rect 262140 21542 262260 21570
rect 262232 16574 262260 21542
rect 263600 18012 263652 18018
rect 263600 17954 263652 17960
rect 263612 16574 263640 17954
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 261484 4888 261536 4894
rect 261484 4830 261536 4836
rect 261404 3454 261800 3482
rect 261772 480 261800 3454
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 264256 11830 264284 127026
rect 264336 121508 264388 121514
rect 264336 121450 264388 121456
rect 264348 32434 264376 121450
rect 264440 54534 264468 131106
rect 264532 103426 264560 144162
rect 264624 122738 264652 161502
rect 264992 155786 265020 210462
rect 265072 207868 265124 207874
rect 265072 207810 265124 207816
rect 265084 158642 265112 207810
rect 265164 183184 265216 183190
rect 265164 183126 265216 183132
rect 265176 164150 265204 183126
rect 266280 176050 266308 229774
rect 266268 176044 266320 176050
rect 266268 175986 266320 175992
rect 266280 175953 266308 175986
rect 266266 175944 266322 175953
rect 266266 175879 266322 175888
rect 265624 169040 265676 169046
rect 265624 168982 265676 168988
rect 265164 164144 265216 164150
rect 265164 164086 265216 164092
rect 265072 158636 265124 158642
rect 265072 158578 265124 158584
rect 264980 155780 265032 155786
rect 264980 155722 265032 155728
rect 264978 149696 265034 149705
rect 264978 149631 265034 149640
rect 264612 122732 264664 122738
rect 264612 122674 264664 122680
rect 264520 103420 264572 103426
rect 264520 103362 264572 103368
rect 264428 54528 264480 54534
rect 264428 54470 264480 54476
rect 264336 32428 264388 32434
rect 264336 32370 264388 32376
rect 264244 11824 264296 11830
rect 264244 11766 264296 11772
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 149631
rect 265636 132394 265664 168982
rect 265624 132388 265676 132394
rect 265624 132330 265676 132336
rect 265716 131776 265768 131782
rect 265716 131718 265768 131724
rect 265624 114572 265676 114578
rect 265624 114514 265676 114520
rect 265636 33862 265664 114514
rect 265728 114510 265756 131718
rect 265716 114504 265768 114510
rect 265716 114446 265768 114452
rect 265624 33856 265676 33862
rect 265624 33798 265676 33804
rect 266372 15162 266400 240094
rect 269224 238882 269252 240094
rect 269212 238876 269264 238882
rect 269212 238818 269264 238824
rect 269120 238808 269172 238814
rect 269120 238750 269172 238756
rect 269132 235634 269160 238750
rect 269224 235822 269252 238818
rect 271800 238513 271828 240638
rect 284208 240644 284260 240650
rect 284208 240586 284260 240592
rect 274054 239850 274082 240108
rect 274008 239822 274082 239850
rect 275986 239850 276014 240108
rect 277918 239850 277946 240108
rect 279436 240094 279864 240122
rect 281552 240094 282440 240122
rect 275986 239822 276060 239850
rect 277918 239822 277992 239850
rect 274008 238785 274036 239822
rect 273994 238776 274050 238785
rect 273994 238711 274050 238720
rect 271786 238504 271842 238513
rect 271786 238439 271842 238448
rect 269212 235816 269264 235822
rect 269212 235758 269264 235764
rect 269304 235816 269356 235822
rect 269304 235758 269356 235764
rect 269316 235634 269344 235758
rect 274008 235754 274036 238711
rect 276032 237250 276060 239822
rect 277964 238241 277992 239822
rect 279436 238678 279464 240094
rect 279424 238672 279476 238678
rect 279424 238614 279476 238620
rect 279436 238377 279464 238614
rect 279422 238368 279478 238377
rect 279422 238303 279478 238312
rect 277950 238232 278006 238241
rect 277950 238167 278006 238176
rect 276020 237244 276072 237250
rect 276020 237186 276072 237192
rect 273996 235748 274048 235754
rect 273996 235690 274048 235696
rect 269132 235606 269344 235634
rect 276032 234394 276060 237186
rect 277964 234530 277992 238167
rect 277952 234524 278004 234530
rect 277952 234466 278004 234472
rect 276020 234388 276072 234394
rect 276020 234330 276072 234336
rect 271236 233980 271288 233986
rect 271236 233922 271288 233928
rect 271248 233102 271276 233922
rect 271236 233096 271288 233102
rect 271236 233038 271288 233044
rect 271248 232121 271276 233038
rect 278686 232520 278742 232529
rect 278686 232455 278742 232464
rect 271234 232112 271290 232121
rect 271234 232047 271290 232056
rect 270406 231160 270462 231169
rect 270406 231095 270462 231104
rect 270316 225684 270368 225690
rect 270316 225626 270368 225632
rect 270328 222902 270356 225626
rect 270316 222896 270368 222902
rect 270316 222838 270368 222844
rect 267832 203652 267884 203658
rect 267832 203594 267884 203600
rect 267740 195424 267792 195430
rect 267740 195366 267792 195372
rect 266544 185836 266596 185842
rect 266544 185778 266596 185784
rect 266452 181552 266504 181558
rect 266452 181494 266504 181500
rect 266464 146198 266492 181494
rect 266556 164218 266584 185778
rect 267096 167136 267148 167142
rect 267096 167078 267148 167084
rect 266544 164212 266596 164218
rect 266544 164154 266596 164160
rect 266452 146192 266504 146198
rect 266452 146134 266504 146140
rect 267004 135312 267056 135318
rect 267004 135254 267056 135260
rect 267016 60110 267044 135254
rect 267108 129606 267136 167078
rect 267752 144906 267780 195366
rect 267844 165578 267872 203594
rect 269212 198144 269264 198150
rect 269212 198086 269264 198092
rect 269120 196784 269172 196790
rect 269120 196726 269172 196732
rect 267924 189984 267976 189990
rect 267924 189926 267976 189932
rect 267832 165572 267884 165578
rect 267832 165514 267884 165520
rect 267936 157350 267964 189926
rect 268476 169856 268528 169862
rect 268476 169798 268528 169804
rect 268384 164892 268436 164898
rect 268384 164834 268436 164840
rect 267924 157344 267976 157350
rect 267924 157286 267976 157292
rect 267740 144900 267792 144906
rect 267740 144842 267792 144848
rect 268396 129674 268424 164834
rect 268488 145654 268516 169798
rect 268476 145648 268528 145654
rect 268476 145590 268528 145596
rect 268568 144968 268620 144974
rect 268568 144910 268620 144916
rect 268384 129668 268436 129674
rect 268384 129610 268436 129616
rect 267096 129600 267148 129606
rect 267096 129542 267148 129548
rect 268476 128376 268528 128382
rect 268476 128318 268528 128324
rect 268384 113212 268436 113218
rect 268384 113154 268436 113160
rect 267832 87644 267884 87650
rect 267832 87586 267884 87592
rect 267004 60104 267056 60110
rect 267004 60046 267056 60052
rect 266452 58812 266504 58818
rect 266452 58754 266504 58760
rect 266464 16574 266492 58754
rect 266464 16546 266584 16574
rect 266360 15156 266412 15162
rect 266360 15098 266412 15104
rect 266372 13258 266400 15098
rect 266360 13252 266412 13258
rect 266360 13194 266412 13200
rect 266556 480 266584 16546
rect 267844 6914 267872 87586
rect 268396 22778 268424 113154
rect 268488 73914 268516 128318
rect 268580 115258 268608 144910
rect 269132 137902 269160 196726
rect 269224 153134 269252 198086
rect 270420 181898 270448 231095
rect 275928 218816 275980 218822
rect 275928 218758 275980 218764
rect 270500 217320 270552 217326
rect 270500 217262 270552 217268
rect 269764 181892 269816 181898
rect 269764 181834 269816 181840
rect 270408 181892 270460 181898
rect 270408 181834 270460 181840
rect 269776 180878 269804 181834
rect 269764 180872 269816 180878
rect 269764 180814 269816 180820
rect 269212 153128 269264 153134
rect 269212 153070 269264 153076
rect 269120 137896 269172 137902
rect 269120 137838 269172 137844
rect 268568 115252 268620 115258
rect 268568 115194 268620 115200
rect 268476 73908 268528 73914
rect 268476 73850 268528 73856
rect 269120 60104 269172 60110
rect 269118 60072 269120 60081
rect 269172 60072 269174 60081
rect 269118 60007 269174 60016
rect 269776 56030 269804 180814
rect 269948 171148 270000 171154
rect 269948 171090 270000 171096
rect 269960 133754 269988 171090
rect 270512 151706 270540 217262
rect 271880 213376 271932 213382
rect 271880 213318 271932 213324
rect 270592 192500 270644 192506
rect 270592 192442 270644 192448
rect 270500 151700 270552 151706
rect 270500 151642 270552 151648
rect 270604 146130 270632 192442
rect 271236 172576 271288 172582
rect 271236 172518 271288 172524
rect 271144 153264 271196 153270
rect 271144 153206 271196 153212
rect 270592 146124 270644 146130
rect 270592 146066 270644 146072
rect 270038 134464 270094 134473
rect 270038 134399 270094 134408
rect 269948 133748 270000 133754
rect 269948 133690 270000 133696
rect 269856 132524 269908 132530
rect 269856 132466 269908 132472
rect 269868 62898 269896 132466
rect 270052 100570 270080 134399
rect 271156 113830 271184 153206
rect 271248 135182 271276 172518
rect 271328 147756 271380 147762
rect 271328 147698 271380 147704
rect 271236 135176 271288 135182
rect 271236 135118 271288 135124
rect 271144 113824 271196 113830
rect 271144 113766 271196 113772
rect 271340 112538 271368 147698
rect 271420 119400 271472 119406
rect 271420 119342 271472 119348
rect 271328 112532 271380 112538
rect 271328 112474 271380 112480
rect 271236 111852 271288 111858
rect 271236 111794 271288 111800
rect 270040 100564 270092 100570
rect 270040 100506 270092 100512
rect 271144 83496 271196 83502
rect 271144 83438 271196 83444
rect 271156 69834 271184 83438
rect 271144 69828 271196 69834
rect 271144 69770 271196 69776
rect 269856 62892 269908 62898
rect 269856 62834 269908 62840
rect 269764 56024 269816 56030
rect 269764 55966 269816 55972
rect 268384 22772 268436 22778
rect 268384 22714 268436 22720
rect 270776 12504 270828 12510
rect 270776 12446 270828 12452
rect 270406 11792 270462 11801
rect 270406 11727 270462 11736
rect 267752 6886 267872 6914
rect 267752 480 267780 6886
rect 268844 3460 268896 3466
rect 268844 3402 268896 3408
rect 268856 480 268884 3402
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 354 270122 480
rect 270420 354 270448 11727
rect 270010 326 270448 354
rect 270788 354 270816 12446
rect 271156 3058 271184 69770
rect 271248 39506 271276 111794
rect 271432 102134 271460 119342
rect 271786 113928 271842 113937
rect 271786 113863 271842 113872
rect 271420 102128 271472 102134
rect 271420 102070 271472 102076
rect 271696 46912 271748 46918
rect 271694 46880 271696 46889
rect 271748 46880 271750 46889
rect 271694 46815 271750 46824
rect 271708 45626 271736 46815
rect 271696 45620 271748 45626
rect 271696 45562 271748 45568
rect 271236 39500 271288 39506
rect 271236 39442 271288 39448
rect 271800 13802 271828 113863
rect 271892 16574 271920 213318
rect 273904 213308 273956 213314
rect 273904 213250 273956 213256
rect 271972 201000 272024 201006
rect 271972 200942 272024 200948
rect 271984 153202 272012 200942
rect 273260 199504 273312 199510
rect 273260 199446 273312 199452
rect 272064 182912 272116 182918
rect 272064 182854 272116 182860
rect 272076 158710 272104 182854
rect 272524 158840 272576 158846
rect 272524 158782 272576 158788
rect 272064 158704 272116 158710
rect 272064 158646 272116 158652
rect 271972 153196 272024 153202
rect 271972 153138 272024 153144
rect 272536 120018 272564 158782
rect 273272 151638 273300 199446
rect 273916 181393 273944 213250
rect 274640 211948 274692 211954
rect 274640 211890 274692 211896
rect 273902 181384 273958 181393
rect 273902 181319 273958 181328
rect 274088 169924 274140 169930
rect 274088 169866 274140 169872
rect 273996 165708 274048 165714
rect 273996 165650 274048 165656
rect 273260 151632 273312 151638
rect 273260 151574 273312 151580
rect 273904 150544 273956 150550
rect 273904 150486 273956 150492
rect 272616 149252 272668 149258
rect 272616 149194 272668 149200
rect 272524 120012 272576 120018
rect 272524 119954 272576 119960
rect 272524 116068 272576 116074
rect 272524 116010 272576 116016
rect 272536 35222 272564 116010
rect 272628 108934 272656 149194
rect 273916 110362 273944 150486
rect 274008 148374 274036 165650
rect 273996 148368 274048 148374
rect 273996 148310 274048 148316
rect 274100 131034 274128 169866
rect 274652 155854 274680 211890
rect 275836 192500 275888 192506
rect 275836 192442 275888 192448
rect 275376 164348 275428 164354
rect 275376 164290 275428 164296
rect 274640 155848 274692 155854
rect 274640 155790 274692 155796
rect 274180 147824 274232 147830
rect 274180 147766 274232 147772
rect 274088 131028 274140 131034
rect 274088 130970 274140 130976
rect 273996 129872 274048 129878
rect 273996 129814 274048 129820
rect 273904 110356 273956 110362
rect 273904 110298 273956 110304
rect 272616 108928 272668 108934
rect 272616 108870 272668 108876
rect 273904 107772 273956 107778
rect 273904 107714 273956 107720
rect 273260 61532 273312 61538
rect 273260 61474 273312 61480
rect 272524 35216 272576 35222
rect 272524 35158 272576 35164
rect 271892 16546 272472 16574
rect 271788 13796 271840 13802
rect 271788 13738 271840 13744
rect 271800 12510 271828 13738
rect 271788 12504 271840 12510
rect 271788 12446 271840 12452
rect 271144 3052 271196 3058
rect 271144 2994 271196 3000
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 270010 -960 270122 326
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 61474
rect 273916 25634 273944 107714
rect 274008 51814 274036 129814
rect 274192 107642 274220 147766
rect 275388 126886 275416 164290
rect 275376 126880 275428 126886
rect 275376 126822 275428 126828
rect 275284 125656 275336 125662
rect 275284 125598 275336 125604
rect 274180 107636 274232 107642
rect 274180 107578 274232 107584
rect 274088 106480 274140 106486
rect 274088 106422 274140 106428
rect 274100 61402 274128 106422
rect 274088 61396 274140 61402
rect 274088 61338 274140 61344
rect 273996 51808 274048 51814
rect 273996 51750 274048 51756
rect 273904 25628 273956 25634
rect 273904 25570 273956 25576
rect 274640 20664 274692 20670
rect 274640 20606 274692 20612
rect 274652 16574 274680 20606
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 275296 9110 275324 125598
rect 275376 109132 275428 109138
rect 275376 109074 275428 109080
rect 275388 66978 275416 109074
rect 275376 66972 275428 66978
rect 275376 66914 275428 66920
rect 275848 20670 275876 192442
rect 275836 20664 275888 20670
rect 275836 20606 275888 20612
rect 275940 15978 275968 218758
rect 276020 216028 276072 216034
rect 276020 215970 276072 215976
rect 276032 149054 276060 215970
rect 277492 207664 277544 207670
rect 277492 207606 277544 207612
rect 277400 203788 277452 203794
rect 277400 203730 277452 203736
rect 276112 181484 276164 181490
rect 276112 181426 276164 181432
rect 276020 149048 276072 149054
rect 276020 148990 276072 148996
rect 276124 147558 276152 181426
rect 276664 180328 276716 180334
rect 276664 180270 276716 180276
rect 276112 147552 276164 147558
rect 276112 147494 276164 147500
rect 276676 95062 276704 180270
rect 277412 147490 277440 203730
rect 277504 154562 277532 207606
rect 278044 175976 278096 175982
rect 278044 175918 278096 175924
rect 277492 154556 277544 154562
rect 277492 154498 277544 154504
rect 277400 147484 277452 147490
rect 277400 147426 277452 147432
rect 276756 136672 276808 136678
rect 276756 136614 276808 136620
rect 276664 95056 276716 95062
rect 276664 94998 276716 95004
rect 276664 79348 276716 79354
rect 276664 79290 276716 79296
rect 275928 15972 275980 15978
rect 275928 15914 275980 15920
rect 275284 9104 275336 9110
rect 275284 9046 275336 9052
rect 276676 3534 276704 79290
rect 276768 58750 276796 136614
rect 276756 58744 276808 58750
rect 276756 58686 276808 58692
rect 277952 15972 278004 15978
rect 277952 15914 278004 15920
rect 276664 3528 276716 3534
rect 276664 3470 276716 3476
rect 277964 3482 277992 15914
rect 278056 3602 278084 175918
rect 278136 151904 278188 151910
rect 278136 151846 278188 151852
rect 278148 113801 278176 151846
rect 278134 113792 278190 113801
rect 278134 113727 278190 113736
rect 278700 4010 278728 232455
rect 278780 231396 278832 231402
rect 278780 231338 278832 231344
rect 278792 16574 278820 231338
rect 279424 231328 279476 231334
rect 279424 231270 279476 231276
rect 278872 194064 278924 194070
rect 278872 194006 278924 194012
rect 278884 155922 278912 194006
rect 279436 178702 279464 231270
rect 281552 229770 281580 240094
rect 282184 231260 282236 231266
rect 282184 231202 282236 231208
rect 281540 229764 281592 229770
rect 281540 229706 281592 229712
rect 281448 224324 281500 224330
rect 281448 224266 281500 224272
rect 280160 206304 280212 206310
rect 280160 206246 280212 206252
rect 279424 178696 279476 178702
rect 279424 178638 279476 178644
rect 279424 174004 279476 174010
rect 279424 173946 279476 173952
rect 278872 155916 278924 155922
rect 278872 155858 278924 155864
rect 279436 136542 279464 173946
rect 279516 154692 279568 154698
rect 279516 154634 279568 154640
rect 279424 136536 279476 136542
rect 279424 136478 279476 136484
rect 279528 131850 279556 154634
rect 279608 142248 279660 142254
rect 279608 142190 279660 142196
rect 279516 131844 279568 131850
rect 279516 131786 279568 131792
rect 279516 120216 279568 120222
rect 279516 120158 279568 120164
rect 279424 113280 279476 113286
rect 279424 113222 279476 113228
rect 279436 37942 279464 113222
rect 279528 65550 279556 120158
rect 279620 100638 279648 142190
rect 280172 139398 280200 206246
rect 280896 160200 280948 160206
rect 280896 160142 280948 160148
rect 280160 139392 280212 139398
rect 280160 139334 280212 139340
rect 280804 135380 280856 135386
rect 280804 135322 280856 135328
rect 279608 100632 279660 100638
rect 279608 100574 279660 100580
rect 279516 65544 279568 65550
rect 279516 65486 279568 65492
rect 280816 61470 280844 135322
rect 280908 121446 280936 160142
rect 280896 121440 280948 121446
rect 280896 121382 280948 121388
rect 280804 61464 280856 61470
rect 280804 61406 280856 61412
rect 281460 53786 281488 224266
rect 281540 207800 281592 207806
rect 281540 207742 281592 207748
rect 281552 137970 281580 207742
rect 281632 195356 281684 195362
rect 281632 195298 281684 195304
rect 281644 150414 281672 195298
rect 281632 150408 281684 150414
rect 281632 150350 281684 150356
rect 281540 137964 281592 137970
rect 281540 137906 281592 137912
rect 281448 53780 281500 53786
rect 281448 53722 281500 53728
rect 281460 52494 281488 53722
rect 280160 52488 280212 52494
rect 280160 52430 280212 52436
rect 281448 52488 281500 52494
rect 281448 52430 281500 52436
rect 279424 37936 279476 37942
rect 279424 37878 279476 37884
rect 280172 16574 280200 52430
rect 281540 21480 281592 21486
rect 281540 21422 281592 21428
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 278688 4004 278740 4010
rect 278688 3946 278740 3952
rect 278044 3596 278096 3602
rect 278044 3538 278096 3544
rect 277964 3454 278360 3482
rect 277124 3324 277176 3330
rect 277124 3266 277176 3272
rect 276020 3052 276072 3058
rect 276020 2994 276072 3000
rect 276032 480 276060 2994
rect 277136 480 277164 3266
rect 278332 480 278360 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 21422
rect 282196 4078 282224 231202
rect 284116 227112 284168 227118
rect 284116 227054 284168 227060
rect 284128 200122 284156 227054
rect 284116 200116 284168 200122
rect 284116 200058 284168 200064
rect 284128 198762 284156 200058
rect 282920 198756 282972 198762
rect 282920 198698 282972 198704
rect 284116 198756 284168 198762
rect 284116 198698 284168 198704
rect 282368 171216 282420 171222
rect 282368 171158 282420 171164
rect 282276 138168 282328 138174
rect 282276 138110 282328 138116
rect 282288 26994 282316 138110
rect 282380 133822 282408 171158
rect 282368 133816 282420 133822
rect 282368 133758 282420 133764
rect 282460 132592 282512 132598
rect 282460 132534 282512 132540
rect 282368 118720 282420 118726
rect 282368 118662 282420 118668
rect 282276 26988 282328 26994
rect 282276 26930 282328 26936
rect 282380 15910 282408 118662
rect 282472 69766 282500 132534
rect 282460 69760 282512 69766
rect 282460 69702 282512 69708
rect 282932 16574 282960 198698
rect 283564 163056 283616 163062
rect 283564 162998 283616 163004
rect 283576 124166 283604 162998
rect 283564 124160 283616 124166
rect 283564 124102 283616 124108
rect 283564 121576 283616 121582
rect 283564 121518 283616 121524
rect 283576 18630 283604 121518
rect 283656 98048 283708 98054
rect 283656 97990 283708 97996
rect 283668 53106 283696 97990
rect 284220 64870 284248 240586
rect 292946 240544 293002 240553
rect 292744 240502 292946 240530
rect 292946 240479 293002 240488
rect 284372 240094 284708 240122
rect 286304 240094 286640 240122
rect 284680 237182 284708 240094
rect 284668 237176 284720 237182
rect 284668 237118 284720 237124
rect 285588 237176 285640 237182
rect 285588 237118 285640 237124
rect 285600 179450 285628 237118
rect 286612 235754 286640 240094
rect 288222 239850 288250 240108
rect 290812 240094 291148 240122
rect 288222 239822 288296 239850
rect 288268 237250 288296 239822
rect 291120 238754 291148 240094
rect 291120 238726 291240 238754
rect 291212 238066 291240 238726
rect 291200 238060 291252 238066
rect 291200 238002 291252 238008
rect 288256 237244 288308 237250
rect 288256 237186 288308 237192
rect 286600 235748 286652 235754
rect 286600 235690 286652 235696
rect 286876 235748 286928 235754
rect 286876 235690 286928 235696
rect 285588 179444 285640 179450
rect 285588 179386 285640 179392
rect 285600 174593 285628 179386
rect 285586 174584 285642 174593
rect 285586 174519 285642 174528
rect 284944 168428 284996 168434
rect 284944 168370 284996 168376
rect 284956 129742 284984 168370
rect 285128 156120 285180 156126
rect 285128 156062 285180 156068
rect 284944 129736 284996 129742
rect 284944 129678 284996 129684
rect 285036 128444 285088 128450
rect 285036 128386 285088 128392
rect 284944 125724 284996 125730
rect 284944 125666 284996 125672
rect 284208 64864 284260 64870
rect 284208 64806 284260 64812
rect 284220 64326 284248 64806
rect 284208 64320 284260 64326
rect 284208 64262 284260 64268
rect 284956 57254 284984 125666
rect 285048 64258 285076 128386
rect 285140 115938 285168 156062
rect 286324 139596 286376 139602
rect 286324 139538 286376 139544
rect 285128 115932 285180 115938
rect 285128 115874 285180 115880
rect 285128 106412 285180 106418
rect 285128 106354 285180 106360
rect 285140 76634 285168 106354
rect 285588 77240 285640 77246
rect 285588 77182 285640 77188
rect 285128 76628 285180 76634
rect 285128 76570 285180 76576
rect 285036 64252 285088 64258
rect 285036 64194 285088 64200
rect 284944 57248 284996 57254
rect 284944 57190 284996 57196
rect 283656 53100 283708 53106
rect 283656 53042 283708 53048
rect 284944 50448 284996 50454
rect 284944 50390 284996 50396
rect 283564 18624 283616 18630
rect 283564 18566 283616 18572
rect 282932 16546 283144 16574
rect 282368 15904 282420 15910
rect 282368 15846 282420 15852
rect 282184 4072 282236 4078
rect 282184 4014 282236 4020
rect 283116 480 283144 16546
rect 284956 13190 284984 50390
rect 284944 13184 284996 13190
rect 284944 13126 284996 13132
rect 284956 3534 284984 13126
rect 285600 6914 285628 77182
rect 286336 49026 286364 139538
rect 286416 115252 286468 115258
rect 286416 115194 286468 115200
rect 286428 103494 286456 115194
rect 286416 103488 286468 103494
rect 286416 103430 286468 103436
rect 286888 77246 286916 235690
rect 288268 230450 288296 237186
rect 288532 236700 288584 236706
rect 288532 236642 288584 236648
rect 288544 233209 288572 236642
rect 289820 234660 289872 234666
rect 289820 234602 289872 234608
rect 288530 233200 288586 233209
rect 288530 233135 288586 233144
rect 289084 231056 289136 231062
rect 289084 230998 289136 231004
rect 288256 230444 288308 230450
rect 288256 230386 288308 230392
rect 286966 218648 287022 218657
rect 286966 218583 287022 218592
rect 286876 77240 286928 77246
rect 286876 77182 286928 77188
rect 286324 49020 286376 49026
rect 286324 48962 286376 48968
rect 286980 12442 287008 218583
rect 287704 202156 287756 202162
rect 287704 202098 287756 202104
rect 287716 176662 287744 202098
rect 287704 176656 287756 176662
rect 287704 176598 287756 176604
rect 287704 174072 287756 174078
rect 287704 174014 287756 174020
rect 287716 136610 287744 174014
rect 287796 172644 287848 172650
rect 287796 172586 287848 172592
rect 287704 136604 287756 136610
rect 287704 136546 287756 136552
rect 287808 135250 287836 172586
rect 287888 161628 287940 161634
rect 287888 161570 287940 161576
rect 287796 135244 287848 135250
rect 287796 135186 287848 135192
rect 287704 131232 287756 131238
rect 287704 131174 287756 131180
rect 285680 12436 285732 12442
rect 285680 12378 285732 12384
rect 286968 12436 287020 12442
rect 286968 12378 287020 12384
rect 285692 11898 285720 12378
rect 285680 11892 285732 11898
rect 285680 11834 285732 11840
rect 285416 6886 285628 6914
rect 284300 3528 284352 3534
rect 284300 3470 284352 3476
rect 284944 3528 284996 3534
rect 284944 3470 284996 3476
rect 284312 480 284340 3470
rect 285416 480 285444 6886
rect 287716 6186 287744 131174
rect 287900 122806 287928 161570
rect 287980 145036 288032 145042
rect 287980 144978 288032 144984
rect 287888 122800 287940 122806
rect 287888 122742 287940 122748
rect 287796 121644 287848 121650
rect 287796 121586 287848 121592
rect 287808 28354 287836 121586
rect 287992 104786 288020 144978
rect 287980 104780 288032 104786
rect 287980 104722 288032 104728
rect 287888 103624 287940 103630
rect 287888 103566 287940 103572
rect 287796 28348 287848 28354
rect 287796 28290 287848 28296
rect 287900 19990 287928 103566
rect 287980 102264 288032 102270
rect 287980 102206 288032 102212
rect 287992 44878 288020 102206
rect 287980 44872 288032 44878
rect 287980 44814 288032 44820
rect 287978 32464 288034 32473
rect 287978 32399 288034 32408
rect 287888 19984 287940 19990
rect 287888 19926 287940 19932
rect 287992 9654 288020 32399
rect 287980 9648 288032 9654
rect 287980 9590 288032 9596
rect 287992 6914 288020 9590
rect 287808 6886 288020 6914
rect 287704 6180 287756 6186
rect 287704 6122 287756 6128
rect 286600 3868 286652 3874
rect 286600 3810 286652 3816
rect 286612 480 286640 3810
rect 287808 480 287836 6886
rect 288992 4004 289044 4010
rect 288992 3946 289044 3952
rect 289004 480 289032 3946
rect 289096 3874 289124 230998
rect 289360 150612 289412 150618
rect 289360 150554 289412 150560
rect 289268 133952 289320 133958
rect 289268 133894 289320 133900
rect 289176 122936 289228 122942
rect 289176 122878 289228 122884
rect 289188 17270 289216 122878
rect 289280 43518 289308 133894
rect 289372 110430 289400 150554
rect 289360 110424 289412 110430
rect 289360 110366 289412 110372
rect 289268 43512 289320 43518
rect 289268 43454 289320 43460
rect 289728 19304 289780 19310
rect 289726 19272 289728 19281
rect 289780 19272 289782 19281
rect 289726 19207 289782 19216
rect 289740 18018 289768 19207
rect 289728 18012 289780 18018
rect 289728 17954 289780 17960
rect 289176 17264 289228 17270
rect 289176 17206 289228 17212
rect 289728 4820 289780 4826
rect 289728 4762 289780 4768
rect 289740 4010 289768 4762
rect 289728 4004 289780 4010
rect 289728 3946 289780 3952
rect 289084 3868 289136 3874
rect 289084 3810 289136 3816
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 234602
rect 291212 215218 291240 238002
rect 291844 236768 291896 236774
rect 291844 236710 291896 236716
rect 291200 215212 291252 215218
rect 291200 215154 291252 215160
rect 290648 172712 290700 172718
rect 290648 172654 290700 172660
rect 290556 140888 290608 140894
rect 290556 140830 290608 140836
rect 290464 134020 290516 134026
rect 290464 133962 290516 133968
rect 290476 40798 290504 133962
rect 290568 99210 290596 140830
rect 290660 133890 290688 172654
rect 290648 133884 290700 133890
rect 290648 133826 290700 133832
rect 290556 99204 290608 99210
rect 290556 99146 290608 99152
rect 291856 48346 291884 236710
rect 292670 198112 292726 198121
rect 292670 198047 292672 198056
rect 292724 198047 292726 198056
rect 292672 198018 292724 198024
rect 293052 192506 293080 258839
rect 293144 213382 293172 325751
rect 293224 299532 293276 299538
rect 293224 299474 293276 299480
rect 293236 238513 293264 299474
rect 293868 259412 293920 259418
rect 293868 259354 293920 259360
rect 293880 259185 293908 259354
rect 293866 259176 293922 259185
rect 293866 259111 293922 259120
rect 293972 246265 294000 461586
rect 294052 362976 294104 362982
rect 294052 362918 294104 362924
rect 294064 305425 294092 362918
rect 294326 323096 294382 323105
rect 294326 323031 294382 323040
rect 294340 322998 294368 323031
rect 294328 322992 294380 322998
rect 294328 322934 294380 322940
rect 294340 316034 294368 322934
rect 294156 316006 294368 316034
rect 294050 305416 294106 305425
rect 294050 305351 294052 305360
rect 294104 305351 294106 305360
rect 294052 305322 294104 305328
rect 294064 305291 294092 305322
rect 294050 299296 294106 299305
rect 294050 299231 294106 299240
rect 294064 291174 294092 299231
rect 294052 291168 294104 291174
rect 294052 291110 294104 291116
rect 293958 246256 294014 246265
rect 293958 246191 294014 246200
rect 293314 241904 293370 241913
rect 293314 241839 293370 241848
rect 293328 241233 293356 241839
rect 293314 241224 293370 241233
rect 293314 241159 293370 241168
rect 293222 238504 293278 238513
rect 293222 238439 293278 238448
rect 293132 213376 293184 213382
rect 293132 213318 293184 213324
rect 293040 192500 293092 192506
rect 293040 192442 293092 192448
rect 293224 165776 293276 165782
rect 293224 165718 293276 165724
rect 292212 158908 292264 158914
rect 292212 158850 292264 158856
rect 292028 129940 292080 129946
rect 292028 129882 292080 129888
rect 291936 124296 291988 124302
rect 291936 124238 291988 124244
rect 291844 48340 291896 48346
rect 291844 48282 291896 48288
rect 290464 40792 290516 40798
rect 290464 40734 290516 40740
rect 291856 4146 291884 48282
rect 291948 9042 291976 124238
rect 292040 46238 292068 129882
rect 292224 120086 292252 158850
rect 293236 126954 293264 165718
rect 293408 157548 293460 157554
rect 293408 157490 293460 157496
rect 293316 136740 293368 136746
rect 293316 136682 293368 136688
rect 293224 126948 293276 126954
rect 293224 126890 293276 126896
rect 292212 120080 292264 120086
rect 292212 120022 292264 120028
rect 292120 118788 292172 118794
rect 292120 118730 292172 118736
rect 292132 53174 292160 118730
rect 293224 117428 293276 117434
rect 293224 117370 293276 117376
rect 292120 53168 292172 53174
rect 292120 53110 292172 53116
rect 292580 47728 292632 47734
rect 292580 47670 292632 47676
rect 292028 46232 292080 46238
rect 292028 46174 292080 46180
rect 292028 35216 292080 35222
rect 292028 35158 292080 35164
rect 291936 9036 291988 9042
rect 291936 8978 291988 8984
rect 291844 4140 291896 4146
rect 291844 4082 291896 4088
rect 292040 4078 292068 35158
rect 291384 4072 291436 4078
rect 291384 4014 291436 4020
rect 292028 4072 292080 4078
rect 292028 4014 292080 4020
rect 291396 480 291424 4014
rect 292592 480 292620 47670
rect 293236 22846 293264 117370
rect 293328 55962 293356 136682
rect 293420 118658 293448 157490
rect 293500 143608 293552 143614
rect 293500 143550 293552 143556
rect 293408 118652 293460 118658
rect 293408 118594 293460 118600
rect 293512 104174 293540 143550
rect 293500 104168 293552 104174
rect 293500 104110 293552 104116
rect 293408 103692 293460 103698
rect 293408 103634 293460 103640
rect 293420 62830 293448 103634
rect 294064 86290 294092 291110
rect 294156 234666 294184 316006
rect 295260 283665 295288 571270
rect 295352 325694 295380 584598
rect 297364 581052 297416 581058
rect 297364 580994 297416 581000
rect 297376 462398 297404 580994
rect 297916 469872 297968 469878
rect 297916 469814 297968 469820
rect 297364 462392 297416 462398
rect 297364 462334 297416 462340
rect 295432 374060 295484 374066
rect 295432 374002 295484 374008
rect 295444 354482 295472 374002
rect 296812 365832 296864 365838
rect 296812 365774 296864 365780
rect 295524 355360 295576 355366
rect 295524 355302 295576 355308
rect 295432 354476 295484 354482
rect 295432 354418 295484 354424
rect 295430 354376 295486 354385
rect 295430 354311 295486 354320
rect 295444 353326 295472 354311
rect 295432 353320 295484 353326
rect 295432 353262 295484 353268
rect 295432 352572 295484 352578
rect 295432 352514 295484 352520
rect 295444 352345 295472 352514
rect 295430 352336 295486 352345
rect 295430 352271 295486 352280
rect 295432 350532 295484 350538
rect 295432 350474 295484 350480
rect 295444 349625 295472 350474
rect 295430 349616 295486 349625
rect 295430 349551 295486 349560
rect 295430 347576 295486 347585
rect 295430 347511 295486 347520
rect 295444 347070 295472 347511
rect 295432 347064 295484 347070
rect 295432 347006 295484 347012
rect 295430 343496 295486 343505
rect 295430 343431 295486 343440
rect 295444 342922 295472 343431
rect 295432 342916 295484 342922
rect 295432 342858 295484 342864
rect 295432 340876 295484 340882
rect 295432 340818 295484 340824
rect 295444 340785 295472 340818
rect 295430 340776 295486 340785
rect 295430 340711 295486 340720
rect 295432 339448 295484 339454
rect 295432 339390 295484 339396
rect 295444 338745 295472 339390
rect 295430 338736 295486 338745
rect 295430 338671 295486 338680
rect 295430 334384 295486 334393
rect 295430 334319 295486 334328
rect 295444 333334 295472 334319
rect 295432 333328 295484 333334
rect 295432 333270 295484 333276
rect 295432 330540 295484 330546
rect 295432 330482 295484 330488
rect 295444 329905 295472 330482
rect 295430 329896 295486 329905
rect 295430 329831 295486 329840
rect 295536 327865 295564 355302
rect 296718 354648 296774 354657
rect 296718 354583 296774 354592
rect 295616 354476 295668 354482
rect 295616 354418 295668 354424
rect 295628 345710 295656 354418
rect 295800 347064 295852 347070
rect 295800 347006 295852 347012
rect 295616 345704 295668 345710
rect 295616 345646 295668 345652
rect 295628 345545 295656 345646
rect 295614 345536 295670 345545
rect 295614 345471 295670 345480
rect 295812 345014 295840 347006
rect 295628 344986 295840 345014
rect 295522 327856 295578 327865
rect 295522 327791 295578 327800
rect 295536 327758 295564 327791
rect 295524 327752 295576 327758
rect 295524 327694 295576 327700
rect 295352 325666 295472 325694
rect 295340 321564 295392 321570
rect 295340 321506 295392 321512
rect 295352 321065 295380 321506
rect 295338 321056 295394 321065
rect 295338 320991 295394 321000
rect 295338 319016 295394 319025
rect 295338 318951 295394 318960
rect 295352 318850 295380 318951
rect 295340 318844 295392 318850
rect 295340 318786 295392 318792
rect 295338 316976 295394 316985
rect 295338 316911 295394 316920
rect 295352 316742 295380 316911
rect 295340 316736 295392 316742
rect 295340 316678 295392 316684
rect 295340 314628 295392 314634
rect 295340 314570 295392 314576
rect 295352 314265 295380 314570
rect 295338 314256 295394 314265
rect 295338 314191 295394 314200
rect 295444 314106 295472 325666
rect 295352 314078 295472 314106
rect 295352 312594 295380 314078
rect 295340 312588 295392 312594
rect 295340 312530 295392 312536
rect 295352 312225 295380 312530
rect 295338 312216 295394 312225
rect 295338 312151 295394 312160
rect 295340 310480 295392 310486
rect 295340 310422 295392 310428
rect 295352 310185 295380 310422
rect 295338 310176 295394 310185
rect 295338 310111 295394 310120
rect 295338 307864 295394 307873
rect 295338 307799 295340 307808
rect 295392 307799 295394 307808
rect 295340 307770 295392 307776
rect 295340 305380 295392 305386
rect 295340 305322 295392 305328
rect 295352 304298 295380 305322
rect 295340 304292 295392 304298
rect 295340 304234 295392 304240
rect 295340 303612 295392 303618
rect 295340 303554 295392 303560
rect 295352 303385 295380 303554
rect 295338 303376 295394 303385
rect 295338 303311 295394 303320
rect 295338 301336 295394 301345
rect 295338 301271 295394 301280
rect 295352 300898 295380 301271
rect 295340 300892 295392 300898
rect 295340 300834 295392 300840
rect 295338 296576 295394 296585
rect 295338 296511 295394 296520
rect 295352 295390 295380 296511
rect 295340 295384 295392 295390
rect 295340 295326 295392 295332
rect 295340 292528 295392 292534
rect 295338 292496 295340 292505
rect 295392 292496 295394 292505
rect 295338 292431 295394 292440
rect 295338 290456 295394 290465
rect 295338 290391 295394 290400
rect 295352 289882 295380 290391
rect 295340 289876 295392 289882
rect 295340 289818 295392 289824
rect 294786 283656 294842 283665
rect 294786 283591 294842 283600
rect 295246 283656 295302 283665
rect 295246 283591 295302 283600
rect 294800 282946 294828 283591
rect 294788 282940 294840 282946
rect 294788 282882 294840 282888
rect 295338 281616 295394 281625
rect 295338 281551 295340 281560
rect 295392 281551 295394 281560
rect 295340 281522 295392 281528
rect 295338 274816 295394 274825
rect 295338 274751 295394 274760
rect 295352 274718 295380 274751
rect 295340 274712 295392 274718
rect 295340 274654 295392 274660
rect 295338 272776 295394 272785
rect 295338 272711 295394 272720
rect 295352 271930 295380 272711
rect 295340 271924 295392 271930
rect 295340 271866 295392 271872
rect 294236 268388 294288 268394
rect 294236 268330 294288 268336
rect 294248 268025 294276 268330
rect 294234 268016 294290 268025
rect 294234 267951 294290 267960
rect 294144 234660 294196 234666
rect 294144 234602 294196 234608
rect 294248 231402 294276 267951
rect 295338 261216 295394 261225
rect 295338 261151 295340 261160
rect 295392 261151 295394 261160
rect 295340 261122 295392 261128
rect 295338 257136 295394 257145
rect 295338 257071 295394 257080
rect 295352 256766 295380 257071
rect 295340 256760 295392 256766
rect 295340 256702 295392 256708
rect 295338 255096 295394 255105
rect 295338 255031 295394 255040
rect 295352 254590 295380 255031
rect 295340 254584 295392 254590
rect 295340 254526 295392 254532
rect 295338 252376 295394 252385
rect 295338 252311 295394 252320
rect 295352 251802 295380 252311
rect 295340 251796 295392 251802
rect 295340 251738 295392 251744
rect 295340 250504 295392 250510
rect 295340 250446 295392 250452
rect 295352 250345 295380 250446
rect 295338 250336 295394 250345
rect 295338 250271 295394 250280
rect 295340 248396 295392 248402
rect 295340 248338 295392 248344
rect 295352 248305 295380 248338
rect 295338 248296 295394 248305
rect 295338 248231 295394 248240
rect 294328 246356 294380 246362
rect 294328 246298 294380 246304
rect 294340 246265 294368 246298
rect 294326 246256 294382 246265
rect 294326 246191 294382 246200
rect 294236 231396 294288 231402
rect 294236 231338 294288 231344
rect 295628 231062 295656 344986
rect 295984 338768 296036 338774
rect 295984 338710 296036 338716
rect 295996 336705 296024 338710
rect 295706 336696 295762 336705
rect 295706 336631 295762 336640
rect 295982 336696 296038 336705
rect 295982 336631 296038 336640
rect 295720 334626 295748 336631
rect 295708 334620 295760 334626
rect 295708 334562 295760 334568
rect 296628 326392 296680 326398
rect 296628 326334 296680 326340
rect 296076 313948 296128 313954
rect 296076 313890 296128 313896
rect 296088 270473 296116 313890
rect 296640 296714 296668 326334
rect 296732 306374 296760 354583
rect 296824 342922 296852 365774
rect 297456 356788 297508 356794
rect 297456 356730 297508 356736
rect 296812 342916 296864 342922
rect 296812 342858 296864 342864
rect 296732 306346 296852 306374
rect 296548 296686 296668 296714
rect 296166 287192 296222 287201
rect 296166 287127 296222 287136
rect 296180 287094 296208 287127
rect 296168 287088 296220 287094
rect 296168 287030 296220 287036
rect 296548 279478 296576 296686
rect 296626 294536 296682 294545
rect 296682 294494 296760 294522
rect 296626 294471 296682 294480
rect 296732 293282 296760 294494
rect 296720 293276 296772 293282
rect 296720 293218 296772 293224
rect 296536 279472 296588 279478
rect 296536 279414 296588 279420
rect 296548 278905 296576 279414
rect 296534 278896 296590 278905
rect 296534 278831 296590 278840
rect 296824 277394 296852 306346
rect 296732 277366 296852 277394
rect 296536 271856 296588 271862
rect 296536 271798 296588 271804
rect 296074 270464 296130 270473
rect 296074 270399 296130 270408
rect 296352 263560 296404 263566
rect 296350 263528 296352 263537
rect 296404 263528 296406 263537
rect 296350 263463 296406 263472
rect 296258 243536 296314 243545
rect 296258 243471 296314 243480
rect 296272 242962 296300 243471
rect 296260 242956 296312 242962
rect 296260 242898 296312 242904
rect 296442 241496 296498 241505
rect 296442 241431 296444 241440
rect 296496 241431 296498 241440
rect 296444 241402 296496 241408
rect 296548 238678 296576 271798
rect 296628 251932 296680 251938
rect 296628 251874 296680 251880
rect 296640 250510 296668 251874
rect 296628 250504 296680 250510
rect 296628 250446 296680 250452
rect 296628 241460 296680 241466
rect 296628 241402 296680 241408
rect 296536 238672 296588 238678
rect 296536 238614 296588 238620
rect 296548 238474 296576 238614
rect 296536 238468 296588 238474
rect 296536 238410 296588 238416
rect 295616 231056 295668 231062
rect 295616 230998 295668 231004
rect 296640 176730 296668 241402
rect 296732 231305 296760 277366
rect 297468 251870 297496 356730
rect 297640 356244 297692 356250
rect 297640 356186 297692 356192
rect 297548 302932 297600 302938
rect 297548 302874 297600 302880
rect 297456 251864 297508 251870
rect 297456 251806 297508 251812
rect 297364 251796 297416 251802
rect 297364 251738 297416 251744
rect 296718 231296 296774 231305
rect 296718 231231 296774 231240
rect 296812 231260 296864 231266
rect 296812 231202 296864 231208
rect 296824 223446 296852 231202
rect 297376 230450 297404 251738
rect 297560 239018 297588 302874
rect 297652 295322 297680 356186
rect 297928 352578 297956 469814
rect 298020 358154 298048 601938
rect 299388 587172 299440 587178
rect 299388 587114 299440 587120
rect 298100 403028 298152 403034
rect 298100 402970 298152 402976
rect 298008 358148 298060 358154
rect 298008 358090 298060 358096
rect 298020 357921 298048 358090
rect 298006 357912 298062 357921
rect 298006 357847 298062 357856
rect 297916 352572 297968 352578
rect 297916 352514 297968 352520
rect 297640 295316 297692 295322
rect 297640 295258 297692 295264
rect 298112 271862 298140 402970
rect 298192 363860 298244 363866
rect 298192 363802 298244 363808
rect 298100 271856 298152 271862
rect 298100 271798 298152 271804
rect 298204 240825 298232 363802
rect 298744 356176 298796 356182
rect 298744 356118 298796 356124
rect 298756 283626 298784 356118
rect 299296 316736 299348 316742
rect 299296 316678 299348 316684
rect 299308 315994 299336 316678
rect 299296 315988 299348 315994
rect 299296 315930 299348 315936
rect 298744 283620 298796 283626
rect 298744 283562 298796 283568
rect 298284 281580 298336 281586
rect 298284 281522 298336 281528
rect 298190 240816 298246 240825
rect 298190 240751 298246 240760
rect 297548 239012 297600 239018
rect 297548 238954 297600 238960
rect 297364 230444 297416 230450
rect 297364 230386 297416 230392
rect 297376 229090 297404 230386
rect 297364 229084 297416 229090
rect 297364 229026 297416 229032
rect 298006 225584 298062 225593
rect 298006 225519 298062 225528
rect 296812 223440 296864 223446
rect 296812 223382 296864 223388
rect 298020 201482 298048 225519
rect 298296 222018 298324 281522
rect 299400 268394 299428 587114
rect 300124 525088 300176 525094
rect 300124 525030 300176 525036
rect 299478 353288 299534 353297
rect 299478 353223 299534 353232
rect 299388 268388 299440 268394
rect 299388 268330 299440 268336
rect 299388 261180 299440 261186
rect 299388 261122 299440 261128
rect 298284 222012 298336 222018
rect 298284 221954 298336 221960
rect 298008 201476 298060 201482
rect 298008 201418 298060 201424
rect 298020 200190 298048 201418
rect 298008 200184 298060 200190
rect 298008 200126 298060 200132
rect 295340 176724 295392 176730
rect 295340 176666 295392 176672
rect 296628 176724 296680 176730
rect 296628 176666 296680 176672
rect 295352 175982 295380 176666
rect 295340 175976 295392 175982
rect 295340 175918 295392 175924
rect 297364 175976 297416 175982
rect 297364 175918 297416 175924
rect 295984 167204 296036 167210
rect 295984 167146 296036 167152
rect 294696 144288 294748 144294
rect 294696 144230 294748 144236
rect 294604 114640 294656 114646
rect 294604 114582 294656 114588
rect 294052 86284 294104 86290
rect 294052 86226 294104 86232
rect 293408 62824 293460 62830
rect 293408 62766 293460 62772
rect 293316 55956 293368 55962
rect 293316 55898 293368 55904
rect 293224 22840 293276 22846
rect 293224 22782 293276 22788
rect 294616 11762 294644 114582
rect 294708 106214 294736 144230
rect 295996 128314 296024 167146
rect 296260 149184 296312 149190
rect 296260 149126 296312 149132
rect 296076 134088 296128 134094
rect 296076 134030 296128 134036
rect 295984 128308 296036 128314
rect 295984 128250 296036 128256
rect 295984 113348 296036 113354
rect 295984 113290 296036 113296
rect 294696 106208 294748 106214
rect 294696 106150 294748 106156
rect 294788 105052 294840 105058
rect 294788 104994 294840 105000
rect 294696 102332 294748 102338
rect 294696 102274 294748 102280
rect 294604 11756 294656 11762
rect 294604 11698 294656 11704
rect 293684 7608 293736 7614
rect 293684 7550 293736 7556
rect 293696 480 293724 7550
rect 294708 2106 294736 102274
rect 294800 47598 294828 104994
rect 295338 84280 295394 84289
rect 295338 84215 295394 84224
rect 295352 82754 295380 84215
rect 295340 82748 295392 82754
rect 295340 82690 295392 82696
rect 294788 47592 294840 47598
rect 294788 47534 294840 47540
rect 295340 43512 295392 43518
rect 295340 43454 295392 43460
rect 295352 16574 295380 43454
rect 295352 16546 295656 16574
rect 294880 16040 294932 16046
rect 294880 15982 294932 15988
rect 294696 2100 294748 2106
rect 294696 2042 294748 2048
rect 294892 480 294920 15982
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 295996 8974 296024 113290
rect 296088 49094 296116 134030
rect 296272 109002 296300 149126
rect 296260 108996 296312 109002
rect 296260 108938 296312 108944
rect 296168 107840 296220 107846
rect 296168 107782 296220 107788
rect 296180 58682 296208 107782
rect 297376 101454 297404 175918
rect 297456 132660 297508 132666
rect 297456 132602 297508 132608
rect 297364 101448 297416 101454
rect 297364 101390 297416 101396
rect 296260 100836 296312 100842
rect 296260 100778 296312 100784
rect 296168 58676 296220 58682
rect 296168 58618 296220 58624
rect 296168 57248 296220 57254
rect 296168 57190 296220 57196
rect 296076 49088 296128 49094
rect 296076 49030 296128 49036
rect 296180 16046 296208 57190
rect 296272 51746 296300 100778
rect 297364 99408 297416 99414
rect 297364 99350 297416 99356
rect 297376 73846 297404 99350
rect 297364 73840 297416 73846
rect 297364 73782 297416 73788
rect 296260 51740 296312 51746
rect 296260 51682 296312 51688
rect 297468 50386 297496 132602
rect 297548 127152 297600 127158
rect 297548 127094 297600 127100
rect 297560 75206 297588 127094
rect 297548 75200 297600 75206
rect 297548 75142 297600 75148
rect 297456 50380 297508 50386
rect 297456 50322 297508 50328
rect 297362 22672 297418 22681
rect 297362 22607 297418 22616
rect 296168 16040 296220 16046
rect 296168 15982 296220 15988
rect 295984 8968 296036 8974
rect 295984 8910 296036 8916
rect 297376 8265 297404 22607
rect 297362 8256 297418 8265
rect 297362 8191 297418 8200
rect 297376 6914 297404 8191
rect 297284 6886 297404 6914
rect 297284 480 297312 6886
rect 298020 3534 298048 200126
rect 299296 177336 299348 177342
rect 299296 177278 299348 177284
rect 298744 135448 298796 135454
rect 298744 135390 298796 135396
rect 298100 49020 298152 49026
rect 298100 48962 298152 48968
rect 298112 48346 298140 48962
rect 298100 48340 298152 48346
rect 298100 48282 298152 48288
rect 298756 47666 298784 135390
rect 298836 117496 298888 117502
rect 298836 117438 298888 117444
rect 298744 47660 298796 47666
rect 298744 47602 298796 47608
rect 298848 44946 298876 117438
rect 299308 95946 299336 177278
rect 299296 95940 299348 95946
rect 299296 95882 299348 95888
rect 298928 95260 298980 95266
rect 298928 95202 298980 95208
rect 298836 44940 298888 44946
rect 298836 44882 298888 44888
rect 298940 25566 298968 95202
rect 299400 86358 299428 261122
rect 299492 224330 299520 353223
rect 299940 342916 299992 342922
rect 299940 342858 299992 342864
rect 299952 336054 299980 342858
rect 299940 336048 299992 336054
rect 299940 335990 299992 335996
rect 299572 276752 299624 276758
rect 299572 276694 299624 276700
rect 299584 233170 299612 276694
rect 300136 254590 300164 525030
rect 300228 392630 300256 612750
rect 327908 611448 327960 611454
rect 327908 611390 327960 611396
rect 306288 607436 306340 607442
rect 306288 607378 306340 607384
rect 305644 601792 305696 601798
rect 305644 601734 305696 601740
rect 304264 568676 304316 568682
rect 304264 568618 304316 568624
rect 303526 522336 303582 522345
rect 303526 522271 303582 522280
rect 303540 521694 303568 522271
rect 303528 521688 303580 521694
rect 303528 521630 303580 521636
rect 301504 461644 301556 461650
rect 301504 461586 301556 461592
rect 300308 407176 300360 407182
rect 300308 407118 300360 407124
rect 300216 392624 300268 392630
rect 300216 392566 300268 392572
rect 300320 365702 300348 407118
rect 300860 367124 300912 367130
rect 300860 367066 300912 367072
rect 300308 365696 300360 365702
rect 300308 365638 300360 365644
rect 300768 365152 300820 365158
rect 300768 365094 300820 365100
rect 300308 357740 300360 357746
rect 300308 357682 300360 357688
rect 300216 322244 300268 322250
rect 300216 322186 300268 322192
rect 300124 254584 300176 254590
rect 300124 254526 300176 254532
rect 300124 250504 300176 250510
rect 300124 250446 300176 250452
rect 299572 233164 299624 233170
rect 299572 233106 299624 233112
rect 299480 224324 299532 224330
rect 299480 224266 299532 224272
rect 300136 222970 300164 250446
rect 300228 241466 300256 322186
rect 300320 307086 300348 357682
rect 300780 347070 300808 365094
rect 300768 347064 300820 347070
rect 300768 347006 300820 347012
rect 300308 307080 300360 307086
rect 300308 307022 300360 307028
rect 300872 303618 300900 367066
rect 301516 367062 301544 461586
rect 302976 383036 303028 383042
rect 302976 382978 303028 382984
rect 302240 369912 302292 369918
rect 302240 369854 302292 369860
rect 301044 367056 301096 367062
rect 301044 366998 301096 367004
rect 301504 367056 301556 367062
rect 301504 366998 301556 367004
rect 301056 365770 301084 366998
rect 301044 365764 301096 365770
rect 301044 365706 301096 365712
rect 300952 364472 301004 364478
rect 300952 364414 301004 364420
rect 300964 330546 300992 364414
rect 301056 339454 301084 365706
rect 301504 354884 301556 354890
rect 301504 354826 301556 354832
rect 301044 339448 301096 339454
rect 301044 339390 301096 339396
rect 301320 339448 301372 339454
rect 301320 339390 301372 339396
rect 301332 338842 301360 339390
rect 301320 338836 301372 338842
rect 301320 338778 301372 338784
rect 300952 330540 301004 330546
rect 300952 330482 301004 330488
rect 301320 330540 301372 330546
rect 301320 330482 301372 330488
rect 301332 329118 301360 330482
rect 301320 329112 301372 329118
rect 301320 329054 301372 329060
rect 300860 303612 300912 303618
rect 300860 303554 300912 303560
rect 300872 303006 300900 303554
rect 300860 303000 300912 303006
rect 300860 302942 300912 302948
rect 300308 300892 300360 300898
rect 300308 300834 300360 300840
rect 300320 289746 300348 300834
rect 300308 289740 300360 289746
rect 300308 289682 300360 289688
rect 300308 280832 300360 280838
rect 300308 280774 300360 280780
rect 300320 276758 300348 280774
rect 300308 276752 300360 276758
rect 300308 276694 300360 276700
rect 301320 275324 301372 275330
rect 301320 275266 301372 275272
rect 301332 274718 301360 275266
rect 300860 274712 300912 274718
rect 300860 274654 300912 274660
rect 301320 274712 301372 274718
rect 301320 274654 301372 274660
rect 300768 254584 300820 254590
rect 300768 254526 300820 254532
rect 300780 253230 300808 254526
rect 300768 253224 300820 253230
rect 300768 253166 300820 253172
rect 300216 241460 300268 241466
rect 300216 241402 300268 241408
rect 300872 230382 300900 274654
rect 301516 267714 301544 354826
rect 301596 300892 301648 300898
rect 301596 300834 301648 300840
rect 301504 267708 301556 267714
rect 301504 267650 301556 267656
rect 301608 246566 301636 300834
rect 301688 271924 301740 271930
rect 301688 271866 301740 271872
rect 301044 246560 301096 246566
rect 301044 246502 301096 246508
rect 301596 246560 301648 246566
rect 301596 246502 301648 246508
rect 301056 246362 301084 246502
rect 301044 246356 301096 246362
rect 301044 246298 301096 246304
rect 300952 242956 301004 242962
rect 300952 242898 301004 242904
rect 300860 230376 300912 230382
rect 300860 230318 300912 230324
rect 300124 222964 300176 222970
rect 300124 222906 300176 222912
rect 300124 218748 300176 218754
rect 300124 218690 300176 218696
rect 300136 180334 300164 218690
rect 300964 218006 300992 242898
rect 301056 231266 301084 246298
rect 301700 240786 301728 271866
rect 302252 241913 302280 369854
rect 302884 354816 302936 354822
rect 302884 354758 302936 354764
rect 302332 350532 302384 350538
rect 302332 350474 302384 350480
rect 302344 349858 302372 350474
rect 302332 349852 302384 349858
rect 302332 349794 302384 349800
rect 302896 262206 302924 354758
rect 302988 350538 303016 382978
rect 302976 350532 303028 350538
rect 302976 350474 303028 350480
rect 302884 262200 302936 262206
rect 302884 262142 302936 262148
rect 302332 256760 302384 256766
rect 302332 256702 302384 256708
rect 302238 241904 302294 241913
rect 302238 241839 302294 241848
rect 301136 240780 301188 240786
rect 301136 240722 301188 240728
rect 301688 240780 301740 240786
rect 301688 240722 301740 240728
rect 301148 240106 301176 240722
rect 301136 240100 301188 240106
rect 301136 240042 301188 240048
rect 301044 231260 301096 231266
rect 301044 231202 301096 231208
rect 302344 224942 302372 256702
rect 302332 224936 302384 224942
rect 302332 224878 302384 224884
rect 300952 218000 301004 218006
rect 300952 217942 301004 217948
rect 300124 180328 300176 180334
rect 300124 180270 300176 180276
rect 300124 171284 300176 171290
rect 300124 171226 300176 171232
rect 300136 132462 300164 171226
rect 300308 164280 300360 164286
rect 300308 164222 300360 164228
rect 300216 135516 300268 135522
rect 300216 135458 300268 135464
rect 300124 132456 300176 132462
rect 300124 132398 300176 132404
rect 300124 123004 300176 123010
rect 300124 122946 300176 122952
rect 299388 86352 299440 86358
rect 299388 86294 299440 86300
rect 299480 25696 299532 25702
rect 299480 25638 299532 25644
rect 298928 25560 298980 25566
rect 298928 25502 298980 25508
rect 298468 4140 298520 4146
rect 298468 4082 298520 4088
rect 298008 3528 298060 3534
rect 298008 3470 298060 3476
rect 298480 480 298508 4082
rect 299492 3482 299520 25638
rect 300136 20058 300164 122946
rect 300228 71126 300256 135458
rect 300320 126274 300348 164222
rect 302976 160268 303028 160274
rect 302976 160210 303028 160216
rect 301504 153332 301556 153338
rect 301504 153274 301556 153280
rect 301516 131782 301544 153274
rect 301688 140956 301740 140962
rect 301688 140898 301740 140904
rect 301504 131776 301556 131782
rect 301504 131718 301556 131724
rect 300308 126268 300360 126274
rect 300308 126210 300360 126216
rect 301504 120284 301556 120290
rect 301504 120226 301556 120232
rect 300400 109200 300452 109206
rect 300400 109142 300452 109148
rect 300308 98116 300360 98122
rect 300308 98058 300360 98064
rect 300216 71120 300268 71126
rect 300216 71062 300268 71068
rect 300320 43450 300348 98058
rect 300412 57322 300440 109142
rect 300400 57316 300452 57322
rect 300400 57258 300452 57264
rect 300308 43444 300360 43450
rect 300308 43386 300360 43392
rect 300768 25696 300820 25702
rect 300768 25638 300820 25644
rect 300780 24818 300808 25638
rect 300768 24812 300820 24818
rect 300768 24754 300820 24760
rect 300124 20052 300176 20058
rect 300124 19994 300176 20000
rect 301516 14482 301544 120226
rect 301596 111920 301648 111926
rect 301596 111862 301648 111868
rect 301608 42158 301636 111862
rect 301700 100706 301728 140898
rect 302988 124914 303016 160210
rect 303068 131300 303120 131306
rect 303068 131242 303120 131248
rect 302976 124908 303028 124914
rect 302976 124850 303028 124856
rect 302884 124364 302936 124370
rect 302884 124306 302936 124312
rect 301780 100768 301832 100774
rect 301780 100710 301832 100716
rect 301688 100700 301740 100706
rect 301688 100642 301740 100648
rect 301792 64190 301820 100710
rect 301780 64184 301832 64190
rect 301780 64126 301832 64132
rect 301596 42152 301648 42158
rect 301596 42094 301648 42100
rect 302238 25528 302294 25537
rect 302238 25463 302294 25472
rect 302252 16574 302280 25463
rect 302252 16546 302832 16574
rect 301504 14476 301556 14482
rect 301504 14418 301556 14424
rect 299570 11792 299626 11801
rect 299570 11727 299626 11736
rect 299584 3602 299612 11727
rect 302056 6316 302108 6322
rect 302056 6258 302108 6264
rect 302068 4146 302096 6258
rect 302056 4140 302108 4146
rect 302056 4082 302108 4088
rect 299572 3596 299624 3602
rect 299572 3538 299624 3544
rect 300768 3596 300820 3602
rect 300768 3538 300820 3544
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3538
rect 302068 3482 302096 4082
rect 301976 3454 302096 3482
rect 302804 3482 302832 16546
rect 302896 6254 302924 124306
rect 302976 118856 303028 118862
rect 302976 118798 303028 118804
rect 302988 31142 303016 118798
rect 303080 76566 303108 131242
rect 303540 102406 303568 521630
rect 303620 502988 303672 502994
rect 303620 502930 303672 502936
rect 303632 502382 303660 502930
rect 303620 502376 303672 502382
rect 303620 502318 303672 502324
rect 303620 307828 303672 307834
rect 303620 307770 303672 307776
rect 303632 234598 303660 307770
rect 303712 262200 303764 262206
rect 303712 262142 303764 262148
rect 303724 260914 303752 262142
rect 303712 260908 303764 260914
rect 303712 260850 303764 260856
rect 303620 234592 303672 234598
rect 303620 234534 303672 234540
rect 303724 226166 303752 260850
rect 304276 233102 304304 568618
rect 305656 568546 305684 601734
rect 305644 568540 305696 568546
rect 305644 568482 305696 568488
rect 304356 502376 304408 502382
rect 304356 502318 304408 502324
rect 304368 302938 304396 502318
rect 305000 363656 305052 363662
rect 305000 363598 305052 363604
rect 305012 363458 305040 363598
rect 305000 363452 305052 363458
rect 305000 363394 305052 363400
rect 304540 357468 304592 357474
rect 304540 357410 304592 357416
rect 304448 333260 304500 333266
rect 304448 333202 304500 333208
rect 304356 302932 304408 302938
rect 304356 302874 304408 302880
rect 304460 261186 304488 333202
rect 304552 316810 304580 357410
rect 304540 316804 304592 316810
rect 304540 316746 304592 316752
rect 305012 315994 305040 363394
rect 305090 354920 305146 354929
rect 305090 354855 305146 354864
rect 305000 315988 305052 315994
rect 305000 315930 305052 315936
rect 305012 315314 305040 315930
rect 305000 315308 305052 315314
rect 305000 315250 305052 315256
rect 305000 312588 305052 312594
rect 305000 312530 305052 312536
rect 305012 311914 305040 312530
rect 305000 311908 305052 311914
rect 305000 311850 305052 311856
rect 304448 261180 304500 261186
rect 304448 261122 304500 261128
rect 304264 233096 304316 233102
rect 304264 233038 304316 233044
rect 303712 226160 303764 226166
rect 303712 226102 303764 226108
rect 305012 223582 305040 311850
rect 305104 292534 305132 354855
rect 305092 292528 305144 292534
rect 305092 292470 305144 292476
rect 305552 292528 305604 292534
rect 305552 292470 305604 292476
rect 305564 291825 305592 292470
rect 305550 291816 305606 291825
rect 305550 291751 305606 291760
rect 305656 240281 305684 568482
rect 305736 513392 305788 513398
rect 305736 513334 305788 513340
rect 305748 458862 305776 513334
rect 305736 458856 305788 458862
rect 305736 458798 305788 458804
rect 305736 446412 305788 446418
rect 305736 446354 305788 446360
rect 305748 363458 305776 446354
rect 305736 363452 305788 363458
rect 305736 363394 305788 363400
rect 306300 321570 306328 607378
rect 319444 606144 319496 606150
rect 319444 606086 319496 606092
rect 308404 604648 308456 604654
rect 308404 604590 308456 604596
rect 307024 600704 307076 600710
rect 307024 600646 307076 600652
rect 306564 411324 306616 411330
rect 306564 411266 306616 411272
rect 306576 406434 306604 411266
rect 306564 406428 306616 406434
rect 306564 406370 306616 406376
rect 306472 387252 306524 387258
rect 306472 387194 306524 387200
rect 306380 357808 306432 357814
rect 306380 357750 306432 357756
rect 305736 321564 305788 321570
rect 305736 321506 305788 321512
rect 306288 321564 306340 321570
rect 306288 321506 306340 321512
rect 305748 320890 305776 321506
rect 305736 320884 305788 320890
rect 305736 320826 305788 320832
rect 306288 289808 306340 289814
rect 306288 289750 306340 289756
rect 305736 278044 305788 278050
rect 305736 277986 305788 277992
rect 305090 240272 305146 240281
rect 305090 240207 305146 240216
rect 305642 240272 305698 240281
rect 305642 240207 305698 240216
rect 305104 238785 305132 240207
rect 305090 238776 305146 238785
rect 305090 238711 305146 238720
rect 305748 229838 305776 277986
rect 306300 273970 306328 289750
rect 306288 273964 306340 273970
rect 306288 273906 306340 273912
rect 306392 240854 306420 357750
rect 306484 313954 306512 387194
rect 307036 383042 307064 600646
rect 307208 547936 307260 547942
rect 307208 547878 307260 547884
rect 307116 523048 307168 523054
rect 307116 522990 307168 522996
rect 307024 383036 307076 383042
rect 307024 382978 307076 382984
rect 306472 313948 306524 313954
rect 306472 313890 306524 313896
rect 307024 293276 307076 293282
rect 307024 293218 307076 293224
rect 306380 240848 306432 240854
rect 306380 240790 306432 240796
rect 305736 229832 305788 229838
rect 305736 229774 305788 229780
rect 305000 223576 305052 223582
rect 305000 223518 305052 223524
rect 304264 209228 304316 209234
rect 304264 209170 304316 209176
rect 304276 180266 304304 209170
rect 307036 189786 307064 293218
rect 307128 235754 307156 522990
rect 307220 420238 307248 547878
rect 307208 420232 307260 420238
rect 307208 420174 307260 420180
rect 307668 411936 307720 411942
rect 307668 411878 307720 411884
rect 307680 411398 307708 411878
rect 307208 411392 307260 411398
rect 307208 411334 307260 411340
rect 307668 411392 307720 411398
rect 307668 411334 307720 411340
rect 307220 238542 307248 411334
rect 307852 364404 307904 364410
rect 307852 364346 307904 364352
rect 307760 357536 307812 357542
rect 307760 357478 307812 357484
rect 307772 289814 307800 357478
rect 307864 310486 307892 364346
rect 307852 310480 307904 310486
rect 307852 310422 307904 310428
rect 307760 289808 307812 289814
rect 307760 289750 307812 289756
rect 308416 259418 308444 604590
rect 312544 604580 312596 604586
rect 312544 604522 312596 604528
rect 311808 599276 311860 599282
rect 311808 599218 311860 599224
rect 309048 596420 309100 596426
rect 309048 596362 309100 596368
rect 309060 527882 309088 596362
rect 309784 589348 309836 589354
rect 309784 589290 309836 589296
rect 309796 536790 309824 589290
rect 311164 542428 311216 542434
rect 311164 542370 311216 542376
rect 309784 536784 309836 536790
rect 309784 536726 309836 536732
rect 309048 527876 309100 527882
rect 309048 527818 309100 527824
rect 309060 527202 309088 527818
rect 309048 527196 309100 527202
rect 309048 527138 309100 527144
rect 309784 527196 309836 527202
rect 309784 527138 309836 527144
rect 308496 454096 308548 454102
rect 308496 454038 308548 454044
rect 308508 395962 308536 454038
rect 308496 395956 308548 395962
rect 308496 395898 308548 395904
rect 309048 395956 309100 395962
rect 309048 395898 309100 395904
rect 308956 310480 309008 310486
rect 308956 310422 309008 310428
rect 308968 309874 308996 310422
rect 308956 309868 309008 309874
rect 308956 309810 309008 309816
rect 308496 276684 308548 276690
rect 308496 276626 308548 276632
rect 308404 259412 308456 259418
rect 308404 259354 308456 259360
rect 307208 238536 307260 238542
rect 307208 238478 307260 238484
rect 308508 237182 308536 276626
rect 308496 237176 308548 237182
rect 308496 237118 308548 237124
rect 307116 235748 307168 235754
rect 307116 235690 307168 235696
rect 307024 189780 307076 189786
rect 307024 189722 307076 189728
rect 307036 189106 307064 189722
rect 307024 189100 307076 189106
rect 307024 189042 307076 189048
rect 307668 189100 307720 189106
rect 307668 189042 307720 189048
rect 304264 180260 304316 180266
rect 304264 180202 304316 180208
rect 307680 175982 307708 189042
rect 309060 182238 309088 395898
rect 309232 369980 309284 369986
rect 309232 369922 309284 369928
rect 309244 369889 309272 369922
rect 309230 369880 309286 369889
rect 309230 369815 309286 369824
rect 309048 182232 309100 182238
rect 309048 182174 309100 182180
rect 309796 180794 309824 527138
rect 310428 505776 310480 505782
rect 310428 505718 310480 505724
rect 310440 505170 310468 505718
rect 310428 505164 310480 505170
rect 310428 505106 310480 505112
rect 310440 489914 310468 505106
rect 310348 489886 310468 489914
rect 310244 371204 310296 371210
rect 310244 371146 310296 371152
rect 310256 369986 310284 371146
rect 310348 370530 310376 489886
rect 310428 474768 310480 474774
rect 310428 474710 310480 474716
rect 310336 370524 310388 370530
rect 310336 370466 310388 370472
rect 310244 369980 310296 369986
rect 310244 369922 310296 369928
rect 309968 367328 310020 367334
rect 309968 367270 310020 367276
rect 309876 295384 309928 295390
rect 309876 295326 309928 295332
rect 309704 180766 309824 180794
rect 308404 178152 308456 178158
rect 308404 178094 308456 178100
rect 307668 175976 307720 175982
rect 307668 175918 307720 175924
rect 307680 175681 307708 175918
rect 307666 175672 307722 175681
rect 307666 175607 307722 175616
rect 307022 175264 307078 175273
rect 307022 175199 307078 175208
rect 306930 173224 306986 173233
rect 306930 173159 306986 173168
rect 306944 172582 306972 173159
rect 306932 172576 306984 172582
rect 306932 172518 306984 172524
rect 306562 170640 306618 170649
rect 306562 170575 306618 170584
rect 306576 169862 306604 170575
rect 306564 169856 306616 169862
rect 306564 169798 306616 169804
rect 306562 169280 306618 169289
rect 306562 169215 306618 169224
rect 306576 168502 306604 169215
rect 304264 168496 304316 168502
rect 304264 168438 304316 168444
rect 306564 168496 306616 168502
rect 306564 168438 306616 168444
rect 304276 131102 304304 168438
rect 306562 166832 306618 166841
rect 306562 166767 306618 166776
rect 306378 166424 306434 166433
rect 306378 166359 306434 166368
rect 306392 165782 306420 166359
rect 306470 165880 306526 165889
rect 306470 165815 306526 165824
rect 306380 165776 306432 165782
rect 306380 165718 306432 165724
rect 306484 165646 306512 165815
rect 306576 165714 306604 166767
rect 306564 165708 306616 165714
rect 306564 165650 306616 165656
rect 306472 165640 306524 165646
rect 306472 165582 306524 165588
rect 306470 165472 306526 165481
rect 306470 165407 306526 165416
rect 306378 164656 306434 164665
rect 306378 164591 306434 164600
rect 306392 164422 306420 164591
rect 306484 164490 306512 165407
rect 306472 164484 306524 164490
rect 306472 164426 306524 164432
rect 306380 164416 306432 164422
rect 306380 164358 306432 164364
rect 306380 164280 306432 164286
rect 306378 164248 306380 164257
rect 306432 164248 306434 164257
rect 306378 164183 306434 164192
rect 306562 163840 306618 163849
rect 306562 163775 306618 163784
rect 306378 163432 306434 163441
rect 306378 163367 306434 163376
rect 306392 163062 306420 163367
rect 306380 163056 306432 163062
rect 306380 162998 306432 163004
rect 306470 163024 306526 163033
rect 306576 162994 306604 163775
rect 306470 162959 306526 162968
rect 306564 162988 306616 162994
rect 306484 162926 306512 162959
rect 306564 162930 306616 162936
rect 306472 162920 306524 162926
rect 306472 162862 306524 162868
rect 306470 162480 306526 162489
rect 306470 162415 306526 162424
rect 306378 161664 306434 161673
rect 306484 161634 306512 162415
rect 306562 162072 306618 162081
rect 306562 162007 306618 162016
rect 306378 161599 306434 161608
rect 306472 161628 306524 161634
rect 306392 161566 306420 161599
rect 306472 161570 306524 161576
rect 306380 161560 306432 161566
rect 306380 161502 306432 161508
rect 306576 161498 306604 162007
rect 306564 161492 306616 161498
rect 306564 161434 306616 161440
rect 306470 161256 306526 161265
rect 306470 161191 306526 161200
rect 306378 160848 306434 160857
rect 306378 160783 306434 160792
rect 306392 160138 306420 160783
rect 306484 160206 306512 161191
rect 306562 160440 306618 160449
rect 306562 160375 306618 160384
rect 306576 160274 306604 160375
rect 306564 160268 306616 160274
rect 306564 160210 306616 160216
rect 306472 160200 306524 160206
rect 306472 160142 306524 160148
rect 306380 160132 306432 160138
rect 306380 160074 306432 160080
rect 306562 160032 306618 160041
rect 306562 159967 306618 159976
rect 306378 159624 306434 159633
rect 306378 159559 306434 159568
rect 306392 158914 306420 159559
rect 306470 159080 306526 159089
rect 306470 159015 306526 159024
rect 306380 158908 306432 158914
rect 306380 158850 306432 158856
rect 306484 158778 306512 159015
rect 306576 158846 306604 159967
rect 306564 158840 306616 158846
rect 306564 158782 306616 158788
rect 306472 158772 306524 158778
rect 306472 158714 306524 158720
rect 306562 158672 306618 158681
rect 306562 158607 306618 158616
rect 306378 158264 306434 158273
rect 306378 158199 306434 158208
rect 306392 157554 306420 158199
rect 306470 157856 306526 157865
rect 306470 157791 306526 157800
rect 306380 157548 306432 157554
rect 306380 157490 306432 157496
rect 306484 157418 306512 157791
rect 306576 157486 306604 158607
rect 306564 157480 306616 157486
rect 306564 157422 306616 157428
rect 306930 157448 306986 157457
rect 306472 157412 306524 157418
rect 306930 157383 306986 157392
rect 306472 157354 306524 157360
rect 306746 155680 306802 155689
rect 306746 155615 306802 155624
rect 306760 154630 306788 155615
rect 306944 155242 306972 157383
rect 306932 155236 306984 155242
rect 306932 155178 306984 155184
rect 306748 154624 306800 154630
rect 306748 154566 306800 154572
rect 306654 153232 306710 153241
rect 306654 153167 306710 153176
rect 306562 152688 306618 152697
rect 306562 152623 306618 152632
rect 305734 152280 305790 152289
rect 305734 152215 305790 152224
rect 305642 149288 305698 149297
rect 305642 149223 305698 149232
rect 304540 146396 304592 146402
rect 304540 146338 304592 146344
rect 304264 131096 304316 131102
rect 304264 131038 304316 131044
rect 304356 129804 304408 129810
rect 304356 129746 304408 129752
rect 304264 110628 304316 110634
rect 304264 110570 304316 110576
rect 303528 102400 303580 102406
rect 303528 102342 303580 102348
rect 303160 99476 303212 99482
rect 303160 99418 303212 99424
rect 303068 76560 303120 76566
rect 303068 76502 303120 76508
rect 303172 60042 303200 99418
rect 303620 71120 303672 71126
rect 303620 71062 303672 71068
rect 303160 60036 303212 60042
rect 303160 59978 303212 59984
rect 302976 31136 303028 31142
rect 302976 31078 303028 31084
rect 303632 16574 303660 71062
rect 303632 16546 303936 16574
rect 302884 6248 302936 6254
rect 302884 6190 302936 6196
rect 302804 3454 303200 3482
rect 301976 480 302004 3454
rect 303172 480 303200 3454
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 304276 7682 304304 110570
rect 304368 33794 304396 129746
rect 304448 117360 304500 117366
rect 304448 117302 304500 117308
rect 304460 66910 304488 117302
rect 304552 106282 304580 146338
rect 305656 111110 305684 149223
rect 305748 116618 305776 152215
rect 306576 151978 306604 152623
rect 306564 151972 306616 151978
rect 306564 151914 306616 151920
rect 306668 149734 306696 153167
rect 306656 149728 306708 149734
rect 306656 149670 306708 149676
rect 307036 145586 307064 175199
rect 307482 174856 307538 174865
rect 307482 174791 307538 174800
rect 307496 174078 307524 174791
rect 307574 174448 307630 174457
rect 307574 174383 307630 174392
rect 307484 174072 307536 174078
rect 307484 174014 307536 174020
rect 307588 174010 307616 174383
rect 307666 174040 307722 174049
rect 307576 174004 307628 174010
rect 307666 173975 307722 173984
rect 307576 173946 307628 173952
rect 307680 173942 307708 173975
rect 307668 173936 307720 173942
rect 307668 173878 307720 173884
rect 307666 173632 307722 173641
rect 307666 173567 307722 173576
rect 307300 172712 307352 172718
rect 307298 172680 307300 172689
rect 307352 172680 307354 172689
rect 307680 172650 307708 173567
rect 307298 172615 307354 172624
rect 307668 172644 307720 172650
rect 307668 172586 307720 172592
rect 307574 172272 307630 172281
rect 307574 172207 307630 172216
rect 307482 171456 307538 171465
rect 307482 171391 307538 171400
rect 307496 171290 307524 171391
rect 307484 171284 307536 171290
rect 307484 171226 307536 171232
rect 307588 171222 307616 172207
rect 307666 171864 307722 171873
rect 307666 171799 307722 171808
rect 307576 171216 307628 171222
rect 307576 171158 307628 171164
rect 307680 171154 307708 171799
rect 307668 171148 307720 171154
rect 307668 171090 307720 171096
rect 307298 171048 307354 171057
rect 307298 170983 307354 170992
rect 307312 169046 307340 170983
rect 307666 170232 307722 170241
rect 307666 170167 307722 170176
rect 307680 169930 307708 170167
rect 307668 169924 307720 169930
rect 307668 169866 307720 169872
rect 307666 169824 307722 169833
rect 307666 169759 307668 169768
rect 307720 169759 307722 169768
rect 307668 169730 307720 169736
rect 307300 169040 307352 169046
rect 307300 168982 307352 168988
rect 307666 168872 307722 168881
rect 307666 168807 307722 168816
rect 307298 168464 307354 168473
rect 307680 168434 307708 168807
rect 307298 168399 307354 168408
rect 307668 168428 307720 168434
rect 307114 165064 307170 165073
rect 307114 164999 307170 165008
rect 307024 145580 307076 145586
rect 307024 145522 307076 145528
rect 306562 145072 306618 145081
rect 306562 145007 306618 145016
rect 306576 144226 306604 145007
rect 306564 144220 306616 144226
rect 306564 144162 306616 144168
rect 306562 140040 306618 140049
rect 306562 139975 306618 139984
rect 306576 139602 306604 139975
rect 306564 139596 306616 139602
rect 306564 139538 306616 139544
rect 306746 137864 306802 137873
rect 306746 137799 306802 137808
rect 306760 136746 306788 137799
rect 307128 137290 307156 164999
rect 307312 164898 307340 168399
rect 307668 168370 307720 168376
rect 307482 168056 307538 168065
rect 307482 167991 307538 168000
rect 307496 167142 307524 167991
rect 307574 167648 307630 167657
rect 307574 167583 307630 167592
rect 307484 167136 307536 167142
rect 307484 167078 307536 167084
rect 307588 167074 307616 167583
rect 307666 167240 307722 167249
rect 307666 167175 307668 167184
rect 307720 167175 307722 167184
rect 307668 167146 307720 167152
rect 307576 167068 307628 167074
rect 307576 167010 307628 167016
rect 307300 164892 307352 164898
rect 307300 164834 307352 164840
rect 307482 157040 307538 157049
rect 307482 156975 307538 156984
rect 307496 156058 307524 156975
rect 307574 156632 307630 156641
rect 307574 156567 307630 156576
rect 307484 156052 307536 156058
rect 307484 155994 307536 156000
rect 307588 155990 307616 156567
rect 307666 156224 307722 156233
rect 307666 156159 307722 156168
rect 307680 156126 307708 156159
rect 307668 156120 307720 156126
rect 307668 156062 307720 156068
rect 307576 155984 307628 155990
rect 307576 155926 307628 155932
rect 307482 155272 307538 155281
rect 307482 155207 307538 155216
rect 307390 154864 307446 154873
rect 307390 154799 307446 154808
rect 307404 153882 307432 154799
rect 307496 154698 307524 155207
rect 307484 154692 307536 154698
rect 307484 154634 307536 154640
rect 307574 154456 307630 154465
rect 307574 154391 307630 154400
rect 307392 153876 307444 153882
rect 307392 153818 307444 153824
rect 307482 153640 307538 153649
rect 307482 153575 307538 153584
rect 307496 152522 307524 153575
rect 307588 153338 307616 154391
rect 307666 154048 307722 154057
rect 307666 153983 307722 153992
rect 307576 153332 307628 153338
rect 307576 153274 307628 153280
rect 307680 153270 307708 153983
rect 307668 153264 307720 153270
rect 307668 153206 307720 153212
rect 307484 152516 307536 152522
rect 307484 152458 307536 152464
rect 307668 151904 307720 151910
rect 307666 151872 307668 151881
rect 307720 151872 307722 151881
rect 307666 151807 307722 151816
rect 307482 151464 307538 151473
rect 307482 151399 307538 151408
rect 307298 151056 307354 151065
rect 307298 150991 307354 151000
rect 307312 150550 307340 150991
rect 307496 150618 307524 151399
rect 307666 150648 307722 150657
rect 307484 150612 307536 150618
rect 307666 150583 307722 150592
rect 307484 150554 307536 150560
rect 307300 150544 307352 150550
rect 307300 150486 307352 150492
rect 307680 150482 307708 150583
rect 307668 150476 307720 150482
rect 307668 150418 307720 150424
rect 307482 150240 307538 150249
rect 307482 150175 307538 150184
rect 307496 149258 307524 150175
rect 307666 149832 307722 149841
rect 307666 149767 307722 149776
rect 307484 149252 307536 149258
rect 307484 149194 307536 149200
rect 307680 149190 307708 149767
rect 307668 149184 307720 149190
rect 307668 149126 307720 149132
rect 307574 148880 307630 148889
rect 307574 148815 307630 148824
rect 307482 148064 307538 148073
rect 307482 147999 307538 148008
rect 307496 147830 307524 147999
rect 307484 147824 307536 147830
rect 307484 147766 307536 147772
rect 307588 147762 307616 148815
rect 307666 148472 307722 148481
rect 307666 148407 307722 148416
rect 307576 147756 307628 147762
rect 307576 147698 307628 147704
rect 307680 147694 307708 148407
rect 307668 147688 307720 147694
rect 307574 147656 307630 147665
rect 307668 147630 307720 147636
rect 307574 147591 307630 147600
rect 307482 147248 307538 147257
rect 307482 147183 307538 147192
rect 307496 146402 307524 147183
rect 307484 146396 307536 146402
rect 307484 146338 307536 146344
rect 307482 145888 307538 145897
rect 307482 145823 307538 145832
rect 307496 145042 307524 145823
rect 307484 145036 307536 145042
rect 307484 144978 307536 144984
rect 307206 144664 307262 144673
rect 307206 144599 307262 144608
rect 307116 137284 307168 137290
rect 307116 137226 307168 137232
rect 306748 136740 306800 136746
rect 306748 136682 306800 136688
rect 306746 136640 306802 136649
rect 306746 136575 306802 136584
rect 306562 136232 306618 136241
rect 306562 136167 306618 136176
rect 306576 135386 306604 136167
rect 306564 135380 306616 135386
rect 306564 135322 306616 135328
rect 306760 135318 306788 136575
rect 306930 135688 306986 135697
rect 306930 135623 306986 135632
rect 306944 135454 306972 135623
rect 306932 135448 306984 135454
rect 306932 135390 306984 135396
rect 306748 135312 306800 135318
rect 306748 135254 306800 135260
rect 307114 131064 307170 131073
rect 307114 130999 307170 131008
rect 307128 129810 307156 130999
rect 307116 129804 307168 129810
rect 307116 129746 307168 129752
rect 306562 129296 306618 129305
rect 306562 129231 306618 129240
rect 306576 128450 306604 129231
rect 307114 128888 307170 128897
rect 307114 128823 307170 128832
rect 306564 128444 306616 128450
rect 306564 128386 306616 128392
rect 307128 128382 307156 128823
rect 307116 128376 307168 128382
rect 307116 128318 307168 128324
rect 307114 127664 307170 127673
rect 307114 127599 307170 127608
rect 306746 127256 306802 127265
rect 306746 127191 306802 127200
rect 306760 127022 306788 127191
rect 307128 127158 307156 127599
rect 307116 127152 307168 127158
rect 307116 127094 307168 127100
rect 306748 127016 306800 127022
rect 306748 126958 306800 126964
rect 306746 125896 306802 125905
rect 306746 125831 306802 125840
rect 306760 125662 306788 125831
rect 306748 125656 306800 125662
rect 306748 125598 306800 125604
rect 306746 125488 306802 125497
rect 306746 125423 306802 125432
rect 306760 124302 306788 125423
rect 307022 124672 307078 124681
rect 307022 124607 307078 124616
rect 306748 124296 306800 124302
rect 306748 124238 306800 124244
rect 306562 123856 306618 123865
rect 306562 123791 306618 123800
rect 306576 122942 306604 123791
rect 306564 122936 306616 122942
rect 306564 122878 306616 122884
rect 306746 121272 306802 121281
rect 306746 121207 306802 121216
rect 306760 120290 306788 121207
rect 306748 120284 306800 120290
rect 306748 120226 306800 120232
rect 306562 118280 306618 118289
rect 306562 118215 306618 118224
rect 306576 117502 306604 118215
rect 306564 117496 306616 117502
rect 306564 117438 306616 117444
rect 306746 117056 306802 117065
rect 306746 116991 306802 117000
rect 305736 116612 305788 116618
rect 305736 116554 305788 116560
rect 306760 116074 306788 116991
rect 306748 116068 306800 116074
rect 306748 116010 306800 116016
rect 306930 114472 306986 114481
rect 306930 114407 306986 114416
rect 306562 114064 306618 114073
rect 306562 113999 306618 114008
rect 306576 113354 306604 113999
rect 306564 113348 306616 113354
rect 306564 113290 306616 113296
rect 306944 113286 306972 114407
rect 306932 113280 306984 113286
rect 306932 113222 306984 113228
rect 305644 111104 305696 111110
rect 305644 111046 305696 111052
rect 305642 107672 305698 107681
rect 305642 107607 305698 107616
rect 304540 106276 304592 106282
rect 304540 106218 304592 106224
rect 304632 104916 304684 104922
rect 304632 104858 304684 104864
rect 304644 71058 304672 104858
rect 304632 71052 304684 71058
rect 304632 70994 304684 71000
rect 304448 66904 304500 66910
rect 304448 66846 304500 66852
rect 304356 33788 304408 33794
rect 304356 33730 304408 33736
rect 305656 28286 305684 107607
rect 305734 106312 305790 106321
rect 305734 106247 305790 106256
rect 305644 28280 305696 28286
rect 305644 28222 305696 28228
rect 305748 26926 305776 106247
rect 305918 105496 305974 105505
rect 305918 105431 305974 105440
rect 305826 101144 305882 101153
rect 305826 101079 305882 101088
rect 305840 36582 305868 101079
rect 305932 69698 305960 105431
rect 306746 101688 306802 101697
rect 306746 101623 306802 101632
rect 306760 100774 306788 101623
rect 306748 100768 306800 100774
rect 306748 100710 306800 100716
rect 305920 69692 305972 69698
rect 305920 69634 305972 69640
rect 305828 36576 305880 36582
rect 305828 36518 305880 36524
rect 305736 26920 305788 26926
rect 305736 26862 305788 26868
rect 305644 25560 305696 25566
rect 305644 25502 305696 25508
rect 304264 7676 304316 7682
rect 304264 7618 304316 7624
rect 305656 5545 305684 25502
rect 307036 21418 307064 124607
rect 307114 124264 307170 124273
rect 307114 124199 307116 124208
rect 307168 124199 307170 124208
rect 307116 124170 307168 124176
rect 307114 123448 307170 123457
rect 307114 123383 307170 123392
rect 307128 123010 307156 123383
rect 307116 123004 307168 123010
rect 307116 122946 307168 122952
rect 307114 115696 307170 115705
rect 307114 115631 307170 115640
rect 307128 39370 307156 115631
rect 307220 112470 307248 144599
rect 307588 144294 307616 147591
rect 307666 146840 307722 146849
rect 307666 146775 307722 146784
rect 307680 146334 307708 146775
rect 307668 146328 307720 146334
rect 307668 146270 307720 146276
rect 307666 145480 307722 145489
rect 307666 145415 307722 145424
rect 307680 144974 307708 145415
rect 307668 144968 307720 144974
rect 307668 144910 307720 144916
rect 307576 144288 307628 144294
rect 307390 144256 307446 144265
rect 307576 144230 307628 144236
rect 307390 144191 307446 144200
rect 307298 143440 307354 143449
rect 307298 143375 307354 143384
rect 307312 119406 307340 143375
rect 307300 119400 307352 119406
rect 307300 119342 307352 119348
rect 307298 116240 307354 116249
rect 307298 116175 307354 116184
rect 307208 112464 307260 112470
rect 307208 112406 307260 112412
rect 307206 98696 307262 98705
rect 307206 98631 307262 98640
rect 307220 80714 307248 98631
rect 307312 90370 307340 116175
rect 307404 115258 307432 144191
rect 307482 143848 307538 143857
rect 307482 143783 307538 143792
rect 307496 143614 307524 143783
rect 307484 143608 307536 143614
rect 307484 143550 307536 143556
rect 307666 143032 307722 143041
rect 307666 142967 307722 142976
rect 307482 142488 307538 142497
rect 307482 142423 307538 142432
rect 307496 142254 307524 142423
rect 307484 142248 307536 142254
rect 307484 142190 307536 142196
rect 307680 142186 307708 142967
rect 307668 142180 307720 142186
rect 307668 142122 307720 142128
rect 307666 142080 307722 142089
rect 307666 142015 307722 142024
rect 307574 141264 307630 141273
rect 307574 141199 307630 141208
rect 307588 140894 307616 141199
rect 307680 140962 307708 142015
rect 307668 140956 307720 140962
rect 307668 140898 307720 140904
rect 307576 140888 307628 140894
rect 307576 140830 307628 140836
rect 307666 140856 307722 140865
rect 307666 140791 307668 140800
rect 307720 140791 307722 140800
rect 307668 140762 307720 140768
rect 307574 140448 307630 140457
rect 307574 140383 307630 140392
rect 307588 139534 307616 140383
rect 307666 139632 307722 139641
rect 307666 139567 307722 139576
rect 307576 139528 307628 139534
rect 307576 139470 307628 139476
rect 307680 139466 307708 139567
rect 307668 139460 307720 139466
rect 307668 139402 307720 139408
rect 307482 139088 307538 139097
rect 307482 139023 307538 139032
rect 307496 138106 307524 139023
rect 307666 138680 307722 138689
rect 307666 138615 307722 138624
rect 307574 138272 307630 138281
rect 307574 138207 307630 138216
rect 307484 138100 307536 138106
rect 307484 138042 307536 138048
rect 307588 138038 307616 138207
rect 307680 138174 307708 138615
rect 307668 138168 307720 138174
rect 307668 138110 307720 138116
rect 307576 138032 307628 138038
rect 307576 137974 307628 137980
rect 307666 137456 307722 137465
rect 307666 137391 307722 137400
rect 307680 136678 307708 137391
rect 307668 136672 307720 136678
rect 307668 136614 307720 136620
rect 307668 135516 307720 135522
rect 307668 135458 307720 135464
rect 307680 135289 307708 135458
rect 307666 135280 307722 135289
rect 307666 135215 307722 135224
rect 307482 134872 307538 134881
rect 307482 134807 307538 134816
rect 307496 134026 307524 134807
rect 307574 134464 307630 134473
rect 307574 134399 307630 134408
rect 307484 134020 307536 134026
rect 307484 133962 307536 133968
rect 307588 133958 307616 134399
rect 307668 134088 307720 134094
rect 307666 134056 307668 134065
rect 307720 134056 307722 134065
rect 307666 133991 307722 134000
rect 307576 133952 307628 133958
rect 307576 133894 307628 133900
rect 307482 133648 307538 133657
rect 307482 133583 307538 133592
rect 307496 132598 307524 133583
rect 307574 133240 307630 133249
rect 307574 133175 307630 133184
rect 307484 132592 307536 132598
rect 307484 132534 307536 132540
rect 307588 132530 307616 133175
rect 307666 132696 307722 132705
rect 307666 132631 307668 132640
rect 307720 132631 307722 132640
rect 307668 132602 307720 132608
rect 307576 132524 307628 132530
rect 307576 132466 307628 132472
rect 307482 132288 307538 132297
rect 307482 132223 307538 132232
rect 307496 131306 307524 132223
rect 307574 131880 307630 131889
rect 307574 131815 307630 131824
rect 307484 131300 307536 131306
rect 307484 131242 307536 131248
rect 307588 131238 307616 131815
rect 307666 131472 307722 131481
rect 307666 131407 307722 131416
rect 307576 131232 307628 131238
rect 307576 131174 307628 131180
rect 307680 131170 307708 131407
rect 307668 131164 307720 131170
rect 307668 131106 307720 131112
rect 307574 130656 307630 130665
rect 307574 130591 307630 130600
rect 307482 130248 307538 130257
rect 307482 130183 307538 130192
rect 307496 129878 307524 130183
rect 307588 130014 307616 130591
rect 307576 130008 307628 130014
rect 307576 129950 307628 129956
rect 307668 129940 307720 129946
rect 307668 129882 307720 129888
rect 307484 129872 307536 129878
rect 307680 129849 307708 129882
rect 307484 129814 307536 129820
rect 307666 129840 307722 129849
rect 307666 129775 307722 129784
rect 307666 128072 307722 128081
rect 307666 128007 307722 128016
rect 307680 127090 307708 128007
rect 307668 127084 307720 127090
rect 307668 127026 307720 127032
rect 307666 126848 307722 126857
rect 307666 126783 307722 126792
rect 307680 125730 307708 126783
rect 307668 125724 307720 125730
rect 307668 125666 307720 125672
rect 307666 125080 307722 125089
rect 307666 125015 307722 125024
rect 307680 124370 307708 125015
rect 307668 124364 307720 124370
rect 307668 124306 307720 124312
rect 307666 123040 307722 123049
rect 307666 122975 307722 122984
rect 307680 122874 307708 122975
rect 307668 122868 307720 122874
rect 307668 122810 307720 122816
rect 307482 122496 307538 122505
rect 307482 122431 307538 122440
rect 307496 121582 307524 122431
rect 307574 122088 307630 122097
rect 307574 122023 307630 122032
rect 307484 121576 307536 121582
rect 307484 121518 307536 121524
rect 307588 121514 307616 122023
rect 307666 121680 307722 121689
rect 307666 121615 307668 121624
rect 307720 121615 307722 121624
rect 307668 121586 307720 121592
rect 307576 121508 307628 121514
rect 307576 121450 307628 121456
rect 307574 120864 307630 120873
rect 307574 120799 307630 120808
rect 307588 120222 307616 120799
rect 307666 120456 307722 120465
rect 307666 120391 307722 120400
rect 307576 120216 307628 120222
rect 307576 120158 307628 120164
rect 307680 120154 307708 120391
rect 307668 120148 307720 120154
rect 307668 120090 307720 120096
rect 307574 120048 307630 120057
rect 307574 119983 307630 119992
rect 307482 119640 307538 119649
rect 307482 119575 307538 119584
rect 307496 118726 307524 119575
rect 307588 118794 307616 119983
rect 307666 119096 307722 119105
rect 307666 119031 307722 119040
rect 307680 118862 307708 119031
rect 307668 118856 307720 118862
rect 307668 118798 307720 118804
rect 307576 118788 307628 118794
rect 307576 118730 307628 118736
rect 307484 118720 307536 118726
rect 307484 118662 307536 118668
rect 307574 118688 307630 118697
rect 307574 118623 307630 118632
rect 307588 117366 307616 118623
rect 307666 117872 307722 117881
rect 307666 117807 307722 117816
rect 307680 117570 307708 117807
rect 307668 117564 307720 117570
rect 307668 117506 307720 117512
rect 307666 117464 307722 117473
rect 307666 117399 307668 117408
rect 307720 117399 307722 117408
rect 307668 117370 307720 117376
rect 307576 117360 307628 117366
rect 307576 117302 307628 117308
rect 307482 116648 307538 116657
rect 307482 116583 307538 116592
rect 307496 116006 307524 116583
rect 307484 116000 307536 116006
rect 307484 115942 307536 115948
rect 307574 115288 307630 115297
rect 307392 115252 307444 115258
rect 307574 115223 307630 115232
rect 307392 115194 307444 115200
rect 307588 114646 307616 115223
rect 307666 114880 307722 114889
rect 307666 114815 307722 114824
rect 307576 114640 307628 114646
rect 307576 114582 307628 114588
rect 307680 114578 307708 114815
rect 307668 114572 307720 114578
rect 307668 114514 307720 114520
rect 307666 113248 307722 113257
rect 307666 113183 307668 113192
rect 307720 113183 307722 113192
rect 307668 113154 307720 113160
rect 307482 112296 307538 112305
rect 307482 112231 307538 112240
rect 307496 111858 307524 112231
rect 307668 111920 307720 111926
rect 307666 111888 307668 111897
rect 307720 111888 307722 111897
rect 307484 111852 307536 111858
rect 307666 111823 307722 111832
rect 307484 111794 307536 111800
rect 307482 111480 307538 111489
rect 307482 111415 307538 111424
rect 307496 110634 307524 111415
rect 307574 111072 307630 111081
rect 307574 111007 307630 111016
rect 307484 110628 307536 110634
rect 307484 110570 307536 110576
rect 307588 110566 307616 111007
rect 307666 110664 307722 110673
rect 307666 110599 307722 110608
rect 307576 110560 307628 110566
rect 307576 110502 307628 110508
rect 307680 110498 307708 110599
rect 307668 110492 307720 110498
rect 307668 110434 307720 110440
rect 307482 110256 307538 110265
rect 307482 110191 307538 110200
rect 307496 109206 307524 110191
rect 307574 109848 307630 109857
rect 307574 109783 307630 109792
rect 307484 109200 307536 109206
rect 307484 109142 307536 109148
rect 307588 109138 307616 109783
rect 307666 109304 307722 109313
rect 307666 109239 307722 109248
rect 307576 109132 307628 109138
rect 307576 109074 307628 109080
rect 307680 109070 307708 109239
rect 307668 109064 307720 109070
rect 307668 109006 307720 109012
rect 307482 108896 307538 108905
rect 307482 108831 307538 108840
rect 307496 107681 307524 108831
rect 307666 108488 307722 108497
rect 307666 108423 307722 108432
rect 307574 108080 307630 108089
rect 307574 108015 307630 108024
rect 307588 107846 307616 108015
rect 307680 107914 307708 108423
rect 307668 107908 307720 107914
rect 307668 107850 307720 107856
rect 307576 107840 307628 107846
rect 307576 107782 307628 107788
rect 307668 107772 307720 107778
rect 307668 107714 307720 107720
rect 307680 107681 307708 107714
rect 307482 107672 307538 107681
rect 307482 107607 307538 107616
rect 307666 107672 307722 107681
rect 307666 107607 307722 107616
rect 307482 107264 307538 107273
rect 307482 107199 307538 107208
rect 307496 106321 307524 107199
rect 308416 106962 308444 178094
rect 309704 178090 309732 180766
rect 309692 178084 309744 178090
rect 309692 178026 309744 178032
rect 309784 176792 309836 176798
rect 309784 176734 309836 176740
rect 308494 146432 308550 146441
rect 308494 146367 308550 146376
rect 308404 106956 308456 106962
rect 308404 106898 308456 106904
rect 307574 106856 307630 106865
rect 307574 106791 307630 106800
rect 307588 106418 307616 106791
rect 307668 106480 307720 106486
rect 307666 106448 307668 106457
rect 307720 106448 307722 106457
rect 307576 106412 307628 106418
rect 307666 106383 307722 106392
rect 307576 106354 307628 106360
rect 307482 106312 307538 106321
rect 307482 106247 307538 106256
rect 307574 105904 307630 105913
rect 307574 105839 307630 105848
rect 307588 104922 307616 105839
rect 307666 105088 307722 105097
rect 307666 105023 307668 105032
rect 307720 105023 307722 105032
rect 307668 104994 307720 105000
rect 307576 104916 307628 104922
rect 307576 104858 307628 104864
rect 308508 104854 308536 146367
rect 308496 104848 308548 104854
rect 308496 104790 308548 104796
rect 307482 104680 307538 104689
rect 307482 104615 307538 104624
rect 307496 103630 307524 104615
rect 307666 104272 307722 104281
rect 307666 104207 307722 104216
rect 307574 103864 307630 103873
rect 307574 103799 307630 103808
rect 307484 103624 307536 103630
rect 307484 103566 307536 103572
rect 307588 103562 307616 103799
rect 307680 103698 307708 104207
rect 307668 103692 307720 103698
rect 307668 103634 307720 103640
rect 307576 103556 307628 103562
rect 307576 103498 307628 103504
rect 307574 103456 307630 103465
rect 307574 103391 307630 103400
rect 307482 103048 307538 103057
rect 307482 102983 307538 102992
rect 307496 102270 307524 102983
rect 307484 102264 307536 102270
rect 307484 102206 307536 102212
rect 307588 102202 307616 103391
rect 307666 102504 307722 102513
rect 307666 102439 307722 102448
rect 307680 102338 307708 102439
rect 308404 102400 308456 102406
rect 308404 102342 308456 102348
rect 307668 102332 307720 102338
rect 307668 102274 307720 102280
rect 307576 102196 307628 102202
rect 307576 102138 307628 102144
rect 307482 102096 307538 102105
rect 307482 102031 307538 102040
rect 307496 101153 307524 102031
rect 307574 101280 307630 101289
rect 307574 101215 307630 101224
rect 307482 101144 307538 101153
rect 307482 101079 307538 101088
rect 307588 100842 307616 101215
rect 307668 100972 307720 100978
rect 307668 100914 307720 100920
rect 307680 100881 307708 100914
rect 307666 100872 307722 100881
rect 307576 100836 307628 100842
rect 307666 100807 307722 100816
rect 307576 100778 307628 100784
rect 307574 100464 307630 100473
rect 307574 100399 307630 100408
rect 307588 99414 307616 100399
rect 307666 99648 307722 99657
rect 307666 99583 307722 99592
rect 307680 99482 307708 99583
rect 307668 99476 307720 99482
rect 307668 99418 307720 99424
rect 307576 99408 307628 99414
rect 307576 99350 307628 99356
rect 307574 99104 307630 99113
rect 307574 99039 307630 99048
rect 307588 98122 307616 99039
rect 307666 98288 307722 98297
rect 307666 98223 307722 98232
rect 307576 98116 307628 98122
rect 307576 98058 307628 98064
rect 307680 98054 307708 98223
rect 307668 98048 307720 98054
rect 307668 97990 307720 97996
rect 307666 97472 307722 97481
rect 307666 97407 307722 97416
rect 307574 97064 307630 97073
rect 307574 96999 307630 97008
rect 307588 96762 307616 96999
rect 307680 96830 307708 97407
rect 307668 96824 307720 96830
rect 307668 96766 307720 96772
rect 307576 96756 307628 96762
rect 307576 96698 307628 96704
rect 307668 96688 307720 96694
rect 307666 96656 307668 96665
rect 307720 96656 307722 96665
rect 307666 96591 307722 96600
rect 307666 96248 307722 96257
rect 307666 96183 307722 96192
rect 307680 95266 307708 96183
rect 307668 95260 307720 95266
rect 307668 95202 307720 95208
rect 308416 93838 308444 102342
rect 309230 100192 309286 100201
rect 309230 100127 309286 100136
rect 308404 93832 308456 93838
rect 308404 93774 308456 93780
rect 307300 90364 307352 90370
rect 307300 90306 307352 90312
rect 308416 82822 308444 93774
rect 308404 82816 308456 82822
rect 308404 82758 308456 82764
rect 307208 80708 307260 80714
rect 307208 80650 307260 80656
rect 307758 42120 307814 42129
rect 307758 42055 307814 42064
rect 307116 39364 307168 39370
rect 307116 39306 307168 39312
rect 307024 21412 307076 21418
rect 307024 21354 307076 21360
rect 307772 16574 307800 42055
rect 309140 27668 309192 27674
rect 309140 27610 309192 27616
rect 307772 16546 307984 16574
rect 305642 5536 305698 5545
rect 305642 5471 305698 5480
rect 305656 4078 305684 5471
rect 305644 4072 305696 4078
rect 305644 4014 305696 4020
rect 306748 4072 306800 4078
rect 306748 4014 306800 4020
rect 305552 3460 305604 3466
rect 305552 3402 305604 3408
rect 305564 480 305592 3402
rect 306760 480 306788 4014
rect 307956 480 307984 16546
rect 309152 6914 309180 27610
rect 309244 7614 309272 100127
rect 309796 80034 309824 176734
rect 309784 80028 309836 80034
rect 309784 79970 309836 79976
rect 309888 32434 309916 295326
rect 309980 177410 310008 367270
rect 310440 335354 310468 474710
rect 310348 335326 310468 335354
rect 310348 327078 310376 335326
rect 310428 327752 310480 327758
rect 310428 327694 310480 327700
rect 310336 327072 310388 327078
rect 310336 327014 310388 327020
rect 310348 326466 310376 327014
rect 310336 326460 310388 326466
rect 310336 326402 310388 326408
rect 310336 324964 310388 324970
rect 310336 324906 310388 324912
rect 310348 316034 310376 324906
rect 310440 321570 310468 327694
rect 310428 321564 310480 321570
rect 310428 321506 310480 321512
rect 310348 316006 310468 316034
rect 310336 295384 310388 295390
rect 310336 295326 310388 295332
rect 310348 295254 310376 295326
rect 310336 295248 310388 295254
rect 310336 295190 310388 295196
rect 310440 240106 310468 316006
rect 310520 282940 310572 282946
rect 310520 282882 310572 282888
rect 310428 240100 310480 240106
rect 310428 240042 310480 240048
rect 310532 230314 310560 282882
rect 311176 251938 311204 542370
rect 311716 536104 311768 536110
rect 311716 536046 311768 536052
rect 311256 347064 311308 347070
rect 311256 347006 311308 347012
rect 311164 251932 311216 251938
rect 311164 251874 311216 251880
rect 310612 240100 310664 240106
rect 310612 240042 310664 240048
rect 310520 230308 310572 230314
rect 310520 230250 310572 230256
rect 310624 187134 310652 240042
rect 311268 213314 311296 347006
rect 311728 281654 311756 536046
rect 311820 340882 311848 599218
rect 311900 504416 311952 504422
rect 311900 504358 311952 504364
rect 311912 503742 311940 504358
rect 311900 503736 311952 503742
rect 311900 503678 311952 503684
rect 311900 380180 311952 380186
rect 311900 380122 311952 380128
rect 311912 379642 311940 380122
rect 311900 379636 311952 379642
rect 311900 379578 311952 379584
rect 311808 340876 311860 340882
rect 311808 340818 311860 340824
rect 311820 340202 311848 340818
rect 311808 340196 311860 340202
rect 311808 340138 311860 340144
rect 311900 289740 311952 289746
rect 311900 289682 311952 289688
rect 311912 289134 311940 289682
rect 312556 289134 312584 604522
rect 317236 601860 317288 601866
rect 317236 601802 317288 601808
rect 313922 599176 313978 599185
rect 313922 599111 313978 599120
rect 312636 503736 312688 503742
rect 312636 503678 312688 503684
rect 311900 289128 311952 289134
rect 311900 289070 311952 289076
rect 312544 289128 312596 289134
rect 312544 289070 312596 289076
rect 311716 281648 311768 281654
rect 311716 281590 311768 281596
rect 312648 238474 312676 503678
rect 312728 379636 312780 379642
rect 312728 379578 312780 379584
rect 312636 238468 312688 238474
rect 312636 238410 312688 238416
rect 312648 238066 312676 238410
rect 312636 238060 312688 238066
rect 312636 238002 312688 238008
rect 311900 234388 311952 234394
rect 311900 234330 311952 234336
rect 311912 233986 311940 234330
rect 312740 233986 312768 379578
rect 313280 368484 313332 368490
rect 313280 368426 313332 368432
rect 313292 367266 313320 368426
rect 313280 367260 313332 367266
rect 313280 367202 313332 367208
rect 311900 233980 311952 233986
rect 311900 233922 311952 233928
rect 312728 233980 312780 233986
rect 312728 233922 312780 233928
rect 313186 217424 313242 217433
rect 313186 217359 313242 217368
rect 313200 216753 313228 217359
rect 313186 216744 313242 216753
rect 313186 216679 313242 216688
rect 311256 213308 311308 213314
rect 311256 213250 311308 213256
rect 311164 208412 311216 208418
rect 311164 208354 311216 208360
rect 310612 187128 310664 187134
rect 310612 187070 310664 187076
rect 309968 177404 310020 177410
rect 309968 177346 310020 177352
rect 311176 177342 311204 208354
rect 313200 180402 313228 216679
rect 313188 180396 313240 180402
rect 313188 180338 313240 180344
rect 311164 177336 311216 177342
rect 311164 177278 311216 177284
rect 313292 176798 313320 367202
rect 313372 319456 313424 319462
rect 313372 319398 313424 319404
rect 313384 318850 313412 319398
rect 313372 318844 313424 318850
rect 313372 318786 313424 318792
rect 313372 281648 313424 281654
rect 313372 281590 313424 281596
rect 313384 237250 313412 281590
rect 313936 243545 313964 599111
rect 314936 576156 314988 576162
rect 314936 576098 314988 576104
rect 314948 575550 314976 576098
rect 314752 575544 314804 575550
rect 314752 575486 314804 575492
rect 314936 575544 314988 575550
rect 314936 575486 314988 575492
rect 314660 565888 314712 565894
rect 314660 565830 314712 565836
rect 314016 520328 314068 520334
rect 314016 520270 314068 520276
rect 314028 368490 314056 520270
rect 314016 368484 314068 368490
rect 314016 368426 314068 368432
rect 314016 365220 314068 365226
rect 314016 365162 314068 365168
rect 314028 297430 314056 365162
rect 314568 319456 314620 319462
rect 314568 319398 314620 319404
rect 314016 297424 314068 297430
rect 314016 297366 314068 297372
rect 313922 243536 313978 243545
rect 313922 243471 313978 243480
rect 313372 237244 313424 237250
rect 313372 237186 313424 237192
rect 314476 231804 314528 231810
rect 314476 231746 314528 231752
rect 314488 231198 314516 231746
rect 314476 231192 314528 231198
rect 314476 231134 314528 231140
rect 313922 187232 313978 187241
rect 313922 187167 313978 187176
rect 313280 176792 313332 176798
rect 313280 176734 313332 176740
rect 313936 175982 313964 187167
rect 314488 178945 314516 231134
rect 314580 228546 314608 319398
rect 314568 228540 314620 228546
rect 314568 228482 314620 228488
rect 314672 216753 314700 565830
rect 314764 231810 314792 575486
rect 315304 566500 315356 566506
rect 315304 566442 315356 566448
rect 315316 565894 315344 566442
rect 315304 565888 315356 565894
rect 315304 565830 315356 565836
rect 317248 527134 317276 601802
rect 317418 597952 317474 597961
rect 317418 597887 317474 597896
rect 317432 595474 317460 597887
rect 317420 595468 317472 595474
rect 317420 595410 317472 595416
rect 318064 594924 318116 594930
rect 318064 594866 318116 594872
rect 317328 562352 317380 562358
rect 317328 562294 317380 562300
rect 317340 561746 317368 562294
rect 317328 561740 317380 561746
rect 317328 561682 317380 561688
rect 317236 527128 317288 527134
rect 317236 527070 317288 527076
rect 314844 526448 314896 526454
rect 314844 526390 314896 526396
rect 314856 525842 314884 526390
rect 317248 525842 317276 527070
rect 314844 525836 314896 525842
rect 314844 525778 314896 525784
rect 315304 525836 315356 525842
rect 315304 525778 315356 525784
rect 317236 525836 317288 525842
rect 317236 525778 317288 525784
rect 315316 238338 315344 525778
rect 317236 388476 317288 388482
rect 317236 388418 317288 388424
rect 317248 387870 317276 388418
rect 316040 387864 316092 387870
rect 316040 387806 316092 387812
rect 317236 387864 317288 387870
rect 317236 387806 317288 387812
rect 315396 363044 315448 363050
rect 315396 362986 315448 362992
rect 315304 238332 315356 238338
rect 315304 238274 315356 238280
rect 315316 238066 315344 238274
rect 315304 238060 315356 238066
rect 315304 238002 315356 238008
rect 314752 231804 314804 231810
rect 314752 231746 314804 231752
rect 314658 216744 314714 216753
rect 314658 216679 314714 216688
rect 315408 182918 315436 362986
rect 315948 222896 316000 222902
rect 315948 222838 316000 222844
rect 315396 182912 315448 182918
rect 315396 182854 315448 182860
rect 314474 178936 314530 178945
rect 314474 178871 314530 178880
rect 315960 177449 315988 222838
rect 316052 208418 316080 387806
rect 316132 360868 316184 360874
rect 316132 360810 316184 360816
rect 316144 248402 316172 360810
rect 316132 248396 316184 248402
rect 316132 248338 316184 248344
rect 317236 248396 317288 248402
rect 317236 248338 317288 248344
rect 317248 247722 317276 248338
rect 317236 247716 317288 247722
rect 317236 247658 317288 247664
rect 317340 239086 317368 561682
rect 317420 525836 317472 525842
rect 317420 525778 317472 525784
rect 316132 239080 316184 239086
rect 316132 239022 316184 239028
rect 317328 239080 317380 239086
rect 317328 239022 317380 239028
rect 316144 235958 316172 239022
rect 316132 235952 316184 235958
rect 316132 235894 316184 235900
rect 317432 235822 317460 525778
rect 317512 431996 317564 432002
rect 317512 431938 317564 431944
rect 317524 360330 317552 431938
rect 318076 411942 318104 594866
rect 318156 587988 318208 587994
rect 318156 587930 318208 587936
rect 318168 560250 318196 587930
rect 318800 582412 318852 582418
rect 318800 582354 318852 582360
rect 318156 560244 318208 560250
rect 318156 560186 318208 560192
rect 318708 468512 318760 468518
rect 318708 468454 318760 468460
rect 318064 411936 318116 411942
rect 318064 411878 318116 411884
rect 317512 360324 317564 360330
rect 317512 360266 317564 360272
rect 317524 325694 317552 360266
rect 318616 345704 318668 345710
rect 318616 345646 318668 345652
rect 317524 325666 317644 325694
rect 317616 314634 317644 325666
rect 317604 314628 317656 314634
rect 317604 314570 317656 314576
rect 318524 314628 318576 314634
rect 318524 314570 318576 314576
rect 318536 313954 318564 314570
rect 318524 313948 318576 313954
rect 318524 313890 318576 313896
rect 318628 256018 318656 345646
rect 318616 256012 318668 256018
rect 318616 255954 318668 255960
rect 318720 246362 318748 468454
rect 318708 246356 318760 246362
rect 318708 246298 318760 246304
rect 318720 245682 318748 246298
rect 318064 245676 318116 245682
rect 318064 245618 318116 245624
rect 318708 245676 318760 245682
rect 318708 245618 318760 245624
rect 317420 235816 317472 235822
rect 317420 235758 317472 235764
rect 318076 235686 318104 245618
rect 318156 242956 318208 242962
rect 318156 242898 318208 242904
rect 318168 235929 318196 242898
rect 318154 235920 318210 235929
rect 318154 235855 318210 235864
rect 318064 235680 318116 235686
rect 318064 235622 318116 235628
rect 318706 226944 318762 226953
rect 318706 226879 318762 226888
rect 318064 220244 318116 220250
rect 318064 220186 318116 220192
rect 316040 208412 316092 208418
rect 316040 208354 316092 208360
rect 316684 202292 316736 202298
rect 316684 202234 316736 202240
rect 316040 178152 316092 178158
rect 316040 178094 316092 178100
rect 315946 177440 316002 177449
rect 315946 177375 316002 177384
rect 313924 175976 313976 175982
rect 316052 175930 316080 178094
rect 316696 177614 316724 202234
rect 316684 177608 316736 177614
rect 316684 177550 316736 177556
rect 318076 177478 318104 220186
rect 318156 189848 318208 189854
rect 318156 189790 318208 189796
rect 318064 177472 318116 177478
rect 318064 177414 318116 177420
rect 318168 176225 318196 189790
rect 318720 177342 318748 226879
rect 318812 222902 318840 582354
rect 319456 295254 319484 606086
rect 324228 606076 324280 606082
rect 324228 606018 324280 606024
rect 321468 603356 321520 603362
rect 321468 603298 321520 603304
rect 320086 582992 320142 583001
rect 320086 582927 320142 582936
rect 320100 582418 320128 582927
rect 320088 582412 320140 582418
rect 320088 582354 320140 582360
rect 320824 411324 320876 411330
rect 320824 411266 320876 411272
rect 320836 385014 320864 411266
rect 321480 392766 321508 603298
rect 323584 596556 323636 596562
rect 323584 596498 323636 596504
rect 322202 583944 322258 583953
rect 322202 583879 322258 583888
rect 322216 539578 322244 583879
rect 322204 539572 322256 539578
rect 322204 539514 322256 539520
rect 321560 529236 321612 529242
rect 321560 529178 321612 529184
rect 321468 392760 321520 392766
rect 321468 392702 321520 392708
rect 320824 385008 320876 385014
rect 320824 384950 320876 384956
rect 321468 385008 321520 385014
rect 321468 384950 321520 384956
rect 320180 370592 320232 370598
rect 320180 370534 320232 370540
rect 319536 367804 319588 367810
rect 319536 367746 319588 367752
rect 319444 295248 319496 295254
rect 319444 295190 319496 295196
rect 318800 222896 318852 222902
rect 318800 222838 318852 222844
rect 319444 209160 319496 209166
rect 319444 209102 319496 209108
rect 318708 177336 318760 177342
rect 318708 177278 318760 177284
rect 319456 176526 319484 209102
rect 319548 183122 319576 367746
rect 319628 320884 319680 320890
rect 319628 320826 319680 320832
rect 319640 225622 319668 320826
rect 320192 229094 320220 370534
rect 320822 356144 320878 356153
rect 320822 356079 320878 356088
rect 320836 314634 320864 356079
rect 320824 314628 320876 314634
rect 320824 314570 320876 314576
rect 321376 234592 321428 234598
rect 321376 234534 321428 234540
rect 321388 233918 321416 234534
rect 321376 233912 321428 233918
rect 321376 233854 321428 233860
rect 320100 229066 320220 229094
rect 320100 228478 320128 229066
rect 320088 228472 320140 228478
rect 320088 228414 320140 228420
rect 319628 225616 319680 225622
rect 319628 225558 319680 225564
rect 319536 183116 319588 183122
rect 319536 183058 319588 183064
rect 320100 177546 320128 228414
rect 321284 184204 321336 184210
rect 321284 184146 321336 184152
rect 320088 177540 320140 177546
rect 320088 177482 320140 177488
rect 319444 176520 319496 176526
rect 319444 176462 319496 176468
rect 318154 176216 318210 176225
rect 318154 176151 318210 176160
rect 313924 175918 313976 175924
rect 316020 175902 316080 175930
rect 321296 165073 321324 184146
rect 321388 176118 321416 233854
rect 321480 186318 321508 384950
rect 321572 233238 321600 529178
rect 322940 501628 322992 501634
rect 322940 501570 322992 501576
rect 322204 434784 322256 434790
rect 322204 434726 322256 434732
rect 322216 395894 322244 434726
rect 322296 420980 322348 420986
rect 322296 420922 322348 420928
rect 322308 397322 322336 420922
rect 322296 397316 322348 397322
rect 322296 397258 322348 397264
rect 322756 397316 322808 397322
rect 322756 397258 322808 397264
rect 322204 395888 322256 395894
rect 322204 395830 322256 395836
rect 321560 233232 321612 233238
rect 321560 233174 321612 233180
rect 321468 186312 321520 186318
rect 321468 186254 321520 186260
rect 321468 176656 321520 176662
rect 321468 176598 321520 176604
rect 321376 176112 321428 176118
rect 321480 176089 321508 176598
rect 321376 176054 321428 176060
rect 321466 176080 321522 176089
rect 321466 176015 321522 176024
rect 321282 165064 321338 165073
rect 321282 164999 321338 165008
rect 321572 142905 321600 233174
rect 322768 230489 322796 397258
rect 322848 395888 322900 395894
rect 322848 395830 322900 395836
rect 322754 230480 322810 230489
rect 322754 230415 322810 230424
rect 322860 209817 322888 395830
rect 322846 209808 322902 209817
rect 322846 209743 322848 209752
rect 322900 209743 322902 209752
rect 322848 209714 322900 209720
rect 322952 208350 322980 501570
rect 323596 402966 323624 596498
rect 323676 427848 323728 427854
rect 323676 427790 323728 427796
rect 323584 402960 323636 402966
rect 323584 402902 323636 402908
rect 323688 394466 323716 427790
rect 323676 394460 323728 394466
rect 323676 394402 323728 394408
rect 323688 393314 323716 394402
rect 323596 393286 323716 393314
rect 323124 383104 323176 383110
rect 323124 383046 323176 383052
rect 323136 226953 323164 383046
rect 323400 239420 323452 239426
rect 323400 239362 323452 239368
rect 323412 235278 323440 239362
rect 323400 235272 323452 235278
rect 323400 235214 323452 235220
rect 323596 227594 323624 393286
rect 324240 392698 324268 606018
rect 327816 599208 327868 599214
rect 327816 599150 327868 599156
rect 327724 599140 327776 599146
rect 327724 599082 327776 599088
rect 326436 597780 326488 597786
rect 326436 597722 326488 597728
rect 325056 595128 325108 595134
rect 325056 595070 325108 595076
rect 324964 587920 325016 587926
rect 324964 587862 325016 587868
rect 324228 392692 324280 392698
rect 324228 392634 324280 392640
rect 323584 227588 323636 227594
rect 323584 227530 323636 227536
rect 323122 226944 323178 226953
rect 323122 226879 323178 226888
rect 323596 226370 323624 227530
rect 323032 226364 323084 226370
rect 323032 226306 323084 226312
rect 323584 226364 323636 226370
rect 323584 226306 323636 226312
rect 322940 208344 322992 208350
rect 322940 208286 322992 208292
rect 322952 207097 322980 208286
rect 322938 207088 322994 207097
rect 322938 207023 322994 207032
rect 322940 200796 322992 200802
rect 322940 200738 322992 200744
rect 321652 182844 321704 182850
rect 321652 182786 321704 182792
rect 321558 142896 321614 142905
rect 321558 142831 321614 142840
rect 321664 133210 321692 182786
rect 321744 176112 321796 176118
rect 321744 176054 321796 176060
rect 321756 171426 321784 176054
rect 321744 171420 321796 171426
rect 321744 171362 321796 171368
rect 322952 137902 322980 200738
rect 323044 149433 323072 226306
rect 324976 218822 325004 587862
rect 325068 319462 325096 595070
rect 325148 568608 325200 568614
rect 325148 568550 325200 568556
rect 325160 399566 325188 568550
rect 326344 532772 326396 532778
rect 326344 532714 326396 532720
rect 325148 399560 325200 399566
rect 325148 399502 325200 399508
rect 325148 349852 325200 349858
rect 325148 349794 325200 349800
rect 325056 319456 325108 319462
rect 325056 319398 325108 319404
rect 325160 237250 325188 349794
rect 325240 338836 325292 338842
rect 325240 338778 325292 338784
rect 325252 286346 325280 338778
rect 325240 286340 325292 286346
rect 325240 286282 325292 286288
rect 326356 237318 326384 532714
rect 326448 356114 326476 597722
rect 327736 571334 327764 599082
rect 327724 571328 327776 571334
rect 327724 571270 327776 571276
rect 327724 485852 327776 485858
rect 327724 485794 327776 485800
rect 326528 431248 326580 431254
rect 326528 431190 326580 431196
rect 326436 356108 326488 356114
rect 326436 356050 326488 356056
rect 326448 309806 326476 356050
rect 326436 309800 326488 309806
rect 326436 309742 326488 309748
rect 325700 237312 325752 237318
rect 325700 237254 325752 237260
rect 326344 237312 326396 237318
rect 326344 237254 326396 237260
rect 325148 237244 325200 237250
rect 325148 237186 325200 237192
rect 324964 218816 325016 218822
rect 324964 218758 325016 218764
rect 324410 191040 324466 191049
rect 324410 190975 324466 190984
rect 323124 188352 323176 188358
rect 323124 188294 323176 188300
rect 323136 151814 323164 188294
rect 323216 185632 323268 185638
rect 323216 185574 323268 185580
rect 323228 153241 323256 185574
rect 324320 172440 324372 172446
rect 324318 172408 324320 172417
rect 324372 172408 324374 172417
rect 324318 172343 324374 172352
rect 324320 171080 324372 171086
rect 324320 171022 324372 171028
rect 324332 170105 324360 171022
rect 324318 170096 324374 170105
rect 324318 170031 324374 170040
rect 324424 169810 324452 190975
rect 324596 188420 324648 188426
rect 324596 188362 324648 188368
rect 324504 180124 324556 180130
rect 324504 180066 324556 180072
rect 324240 169782 324452 169810
rect 324240 169266 324268 169782
rect 324320 169720 324372 169726
rect 324320 169662 324372 169668
rect 324332 169425 324360 169662
rect 324412 169652 324464 169658
rect 324412 169594 324464 169600
rect 324318 169416 324374 169425
rect 324318 169351 324374 169360
rect 324240 169238 324360 169266
rect 324332 167793 324360 169238
rect 324424 168609 324452 169594
rect 324410 168600 324466 168609
rect 324410 168535 324466 168544
rect 324318 167784 324374 167793
rect 324318 167719 324374 167728
rect 324320 165572 324372 165578
rect 324320 165514 324372 165520
rect 324332 165481 324360 165514
rect 324318 165472 324374 165481
rect 324318 165407 324374 165416
rect 324412 164212 324464 164218
rect 324412 164154 324464 164160
rect 324320 164076 324372 164082
rect 324320 164018 324372 164024
rect 324332 163985 324360 164018
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324424 163169 324452 164154
rect 324410 163160 324466 163169
rect 324410 163095 324466 163104
rect 324320 161424 324372 161430
rect 324320 161366 324372 161372
rect 324332 160857 324360 161366
rect 324318 160848 324374 160857
rect 324318 160783 324374 160792
rect 324516 160177 324544 180066
rect 324608 174729 324636 188362
rect 324688 187060 324740 187066
rect 324688 187002 324740 187008
rect 324594 174720 324650 174729
rect 324594 174655 324650 174664
rect 324502 160168 324558 160177
rect 324502 160103 324558 160112
rect 324320 160064 324372 160070
rect 324320 160006 324372 160012
rect 324332 159361 324360 160006
rect 324318 159352 324374 159361
rect 324318 159287 324374 159296
rect 324412 158704 324464 158710
rect 324412 158646 324464 158652
rect 324320 158636 324372 158642
rect 324320 158578 324372 158584
rect 324332 158545 324360 158578
rect 324318 158536 324374 158545
rect 324318 158471 324374 158480
rect 324424 157865 324452 158646
rect 324410 157856 324466 157865
rect 324410 157791 324466 157800
rect 324412 157344 324464 157350
rect 324412 157286 324464 157292
rect 324320 157072 324372 157078
rect 324318 157040 324320 157049
rect 324372 157040 324374 157049
rect 324318 156975 324374 156984
rect 324424 156369 324452 157286
rect 324410 156360 324466 156369
rect 324410 156295 324466 156304
rect 324320 155916 324372 155922
rect 324320 155858 324372 155864
rect 324332 154737 324360 155858
rect 324700 155553 324728 187002
rect 324686 155544 324742 155553
rect 324686 155479 324742 155488
rect 324318 154728 324374 154737
rect 324318 154663 324374 154672
rect 324320 154352 324372 154358
rect 324320 154294 324372 154300
rect 324332 154057 324360 154294
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 323214 153232 323270 153241
rect 323214 153167 323270 153176
rect 324320 153196 324372 153202
rect 324320 153138 324372 153144
rect 324332 152425 324360 153138
rect 324318 152416 324374 152425
rect 324318 152351 324374 152360
rect 323136 151786 323440 151814
rect 323030 149424 323086 149433
rect 323030 149359 323086 149368
rect 322940 137896 322992 137902
rect 322940 137838 322992 137844
rect 323308 137896 323360 137902
rect 323308 137838 323360 137844
rect 323320 137057 323348 137838
rect 323306 137048 323362 137057
rect 323306 136983 323362 136992
rect 323412 136610 323440 151786
rect 324320 151768 324372 151774
rect 324318 151736 324320 151745
rect 324372 151736 324374 151745
rect 324318 151671 324374 151680
rect 324320 151360 324372 151366
rect 324320 151302 324372 151308
rect 324332 150929 324360 151302
rect 324318 150920 324374 150929
rect 324318 150855 324374 150864
rect 325606 150104 325662 150113
rect 325712 150090 325740 237254
rect 326540 234598 326568 431190
rect 327354 405648 327410 405657
rect 327354 405583 327410 405592
rect 327368 404977 327396 405583
rect 327354 404968 327410 404977
rect 327354 404903 327410 404912
rect 327172 387116 327224 387122
rect 327172 387058 327224 387064
rect 326528 234592 326580 234598
rect 326528 234534 326580 234540
rect 327080 192772 327132 192778
rect 327080 192714 327132 192720
rect 325884 186312 325936 186318
rect 325884 186254 325936 186260
rect 325792 177608 325844 177614
rect 325792 177550 325844 177556
rect 325804 171737 325832 177550
rect 325790 171728 325846 171737
rect 325790 171663 325846 171672
rect 325792 171420 325844 171426
rect 325792 171362 325844 171368
rect 325662 150062 325740 150090
rect 325606 150039 325662 150048
rect 324412 149048 324464 149054
rect 324412 148990 324464 148996
rect 324320 148980 324372 148986
rect 324320 148922 324372 148928
rect 324332 148617 324360 148922
rect 324318 148608 324374 148617
rect 324318 148543 324374 148552
rect 324424 147801 324452 148990
rect 324410 147792 324466 147801
rect 324410 147727 324466 147736
rect 324320 147552 324372 147558
rect 324320 147494 324372 147500
rect 324332 147121 324360 147494
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 324318 146296 324374 146305
rect 324318 146231 324320 146240
rect 324372 146231 324374 146240
rect 324320 146202 324372 146208
rect 324412 146192 324464 146198
rect 324412 146134 324464 146140
rect 324424 145489 324452 146134
rect 324410 145480 324466 145489
rect 324410 145415 324466 145424
rect 324412 144900 324464 144906
rect 324412 144842 324464 144848
rect 324320 144832 324372 144838
rect 324318 144800 324320 144809
rect 324372 144800 324374 144809
rect 324318 144735 324374 144744
rect 324424 143993 324452 144842
rect 324410 143984 324466 143993
rect 324410 143919 324466 143928
rect 324964 143608 325016 143614
rect 324964 143550 325016 143556
rect 324320 143540 324372 143546
rect 324320 143482 324372 143488
rect 324332 143177 324360 143482
rect 324318 143168 324374 143177
rect 324318 143103 324374 143112
rect 324412 142112 324464 142118
rect 324412 142054 324464 142060
rect 324320 141840 324372 141846
rect 324320 141782 324372 141788
rect 324332 141681 324360 141782
rect 324318 141672 324374 141681
rect 324318 141607 324374 141616
rect 324424 140865 324452 142054
rect 324410 140856 324466 140865
rect 324410 140791 324466 140800
rect 324320 140752 324372 140758
rect 324320 140694 324372 140700
rect 324332 140185 324360 140694
rect 324318 140176 324374 140185
rect 324318 140111 324374 140120
rect 324320 139324 324372 139330
rect 324320 139266 324372 139272
rect 324332 138553 324360 139266
rect 324318 138544 324374 138553
rect 324318 138479 324374 138488
rect 324320 137964 324372 137970
rect 324320 137906 324372 137912
rect 324332 137873 324360 137906
rect 324318 137864 324374 137873
rect 324318 137799 324374 137808
rect 323400 136604 323452 136610
rect 323400 136546 323452 136552
rect 323412 136377 323440 136546
rect 324320 136536 324372 136542
rect 324320 136478 324372 136484
rect 323398 136368 323454 136377
rect 323398 136303 323454 136312
rect 324332 135561 324360 136478
rect 324318 135552 324374 135561
rect 324318 135487 324374 135496
rect 324412 135244 324464 135250
rect 324412 135186 324464 135192
rect 324320 135176 324372 135182
rect 324320 135118 324372 135124
rect 324332 134745 324360 135118
rect 324318 134736 324374 134745
rect 324318 134671 324374 134680
rect 324424 134065 324452 135186
rect 324410 134056 324466 134065
rect 324410 133991 324466 134000
rect 324320 133884 324372 133890
rect 324320 133826 324372 133832
rect 324332 133249 324360 133826
rect 324318 133240 324374 133249
rect 321652 133204 321704 133210
rect 324318 133175 324374 133184
rect 321652 133146 321704 133152
rect 321664 122233 321692 133146
rect 323490 131880 323546 131889
rect 323490 131815 323546 131824
rect 323504 131209 323532 131815
rect 323490 131200 323546 131209
rect 323490 131135 323546 131144
rect 324412 131096 324464 131102
rect 324412 131038 324464 131044
rect 324320 131028 324372 131034
rect 324320 130970 324372 130976
rect 324332 130937 324360 130970
rect 324318 130928 324374 130937
rect 324318 130863 324374 130872
rect 324424 130121 324452 131038
rect 324410 130112 324466 130121
rect 324410 130047 324466 130056
rect 324412 129736 324464 129742
rect 324412 129678 324464 129684
rect 324320 129464 324372 129470
rect 324318 129432 324320 129441
rect 324372 129432 324374 129441
rect 324318 129367 324374 129376
rect 324424 128625 324452 129678
rect 324410 128616 324466 128625
rect 324410 128551 324466 128560
rect 324320 128308 324372 128314
rect 324320 128250 324372 128256
rect 324332 127809 324360 128250
rect 324412 128240 324464 128246
rect 324412 128182 324464 128188
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324424 127129 324452 128182
rect 324410 127120 324466 127129
rect 324410 127055 324466 127064
rect 324320 125588 324372 125594
rect 324320 125530 324372 125536
rect 324332 124817 324360 125530
rect 324318 124808 324374 124817
rect 324318 124743 324374 124752
rect 323490 123448 323546 123457
rect 323490 123383 323546 123392
rect 323504 122913 323532 123383
rect 323490 122904 323546 122913
rect 323490 122839 323546 122848
rect 324320 122800 324372 122806
rect 324320 122742 324372 122748
rect 324332 122505 324360 122742
rect 324318 122496 324374 122505
rect 324318 122431 324374 122440
rect 321650 122224 321706 122233
rect 321650 122159 321706 122168
rect 324320 121440 324372 121446
rect 324320 121382 324372 121388
rect 324332 120873 324360 121382
rect 324412 121372 324464 121378
rect 324412 121314 324464 121320
rect 324318 120864 324374 120873
rect 324318 120799 324374 120808
rect 324424 120193 324452 121314
rect 324410 120184 324466 120193
rect 324410 120119 324466 120128
rect 324320 120080 324372 120086
rect 324320 120022 324372 120028
rect 324332 119377 324360 120022
rect 324318 119368 324374 119377
rect 324318 119303 324374 119312
rect 324320 118652 324372 118658
rect 324320 118594 324372 118600
rect 324332 117881 324360 118594
rect 324976 118561 325004 143550
rect 325606 126304 325662 126313
rect 325804 126290 325832 171362
rect 325896 161673 325924 186254
rect 327092 184210 327120 192714
rect 327080 184204 327132 184210
rect 327080 184146 327132 184152
rect 325974 177304 326030 177313
rect 325974 177239 326030 177248
rect 325882 161664 325938 161673
rect 325882 161599 325938 161608
rect 325988 157078 326016 177239
rect 327080 176520 327132 176526
rect 327080 176462 327132 176468
rect 327092 172446 327120 176462
rect 327080 172440 327132 172446
rect 327080 172382 327132 172388
rect 327184 164082 327212 387058
rect 327264 226228 327316 226234
rect 327264 226170 327316 226176
rect 327172 164076 327224 164082
rect 327172 164018 327224 164024
rect 326436 160744 326488 160750
rect 326436 160686 326488 160692
rect 325976 157072 326028 157078
rect 325976 157014 326028 157020
rect 326448 154358 326476 160686
rect 326436 154352 326488 154358
rect 326436 154294 326488 154300
rect 327276 141846 327304 226170
rect 327368 151366 327396 404903
rect 327736 226234 327764 485794
rect 327828 456074 327856 599150
rect 327920 591326 327948 611390
rect 331126 601760 331182 601769
rect 331126 601695 331182 601704
rect 328366 600536 328422 600545
rect 328366 600471 328422 600480
rect 327908 591320 327960 591326
rect 327908 591262 327960 591268
rect 328276 491360 328328 491366
rect 328276 491302 328328 491308
rect 328288 485858 328316 491302
rect 328276 485852 328328 485858
rect 328276 485794 328328 485800
rect 327908 479528 327960 479534
rect 327908 479470 327960 479476
rect 327816 456068 327868 456074
rect 327816 456010 327868 456016
rect 327816 451920 327868 451926
rect 327816 451862 327868 451868
rect 327828 405657 327856 451862
rect 327814 405648 327870 405657
rect 327814 405583 327870 405592
rect 327920 387122 327948 479470
rect 328380 396681 328408 600471
rect 329196 596488 329248 596494
rect 329196 596430 329248 596436
rect 329102 594824 329158 594833
rect 329102 594759 329158 594768
rect 329116 543726 329144 594759
rect 329208 561678 329236 596430
rect 331036 596284 331088 596290
rect 331036 596226 331088 596232
rect 329748 576904 329800 576910
rect 329748 576846 329800 576852
rect 329196 561672 329248 561678
rect 329196 561614 329248 561620
rect 329104 543720 329156 543726
rect 329104 543662 329156 543668
rect 329104 528964 329156 528970
rect 329104 528906 329156 528912
rect 328460 405680 328512 405686
rect 328460 405622 328512 405628
rect 328472 405006 328500 405622
rect 328460 405000 328512 405006
rect 328460 404942 328512 404948
rect 328366 396672 328422 396681
rect 328366 396607 328422 396616
rect 327908 387116 327960 387122
rect 327908 387058 327960 387064
rect 327724 226228 327776 226234
rect 327724 226170 327776 226176
rect 328472 169658 328500 404942
rect 328552 222080 328604 222086
rect 328552 222022 328604 222028
rect 328460 169652 328512 169658
rect 328460 169594 328512 169600
rect 327816 168428 327868 168434
rect 327816 168370 327868 168376
rect 327356 151360 327408 151366
rect 327356 151302 327408 151308
rect 327724 146940 327776 146946
rect 327724 146882 327776 146888
rect 327264 141840 327316 141846
rect 327264 141782 327316 141788
rect 327080 134564 327132 134570
rect 327080 134506 327132 134512
rect 327092 129470 327120 134506
rect 327080 129464 327132 129470
rect 327080 129406 327132 129412
rect 325662 126262 325832 126290
rect 325606 126239 325662 126248
rect 325056 119400 325108 119406
rect 325056 119342 325108 119348
rect 324962 118552 325018 118561
rect 324962 118487 325018 118496
rect 324318 117872 324374 117881
rect 324318 117807 324374 117816
rect 324320 116612 324372 116618
rect 324320 116554 324372 116560
rect 324332 116385 324360 116554
rect 324318 116376 324374 116385
rect 324318 116311 324374 116320
rect 324320 115932 324372 115938
rect 324320 115874 324372 115880
rect 324332 115569 324360 115874
rect 324318 115560 324374 115569
rect 324318 115495 324374 115504
rect 324964 115320 325016 115326
rect 324964 115262 325016 115268
rect 323584 115252 323636 115258
rect 323584 115194 323636 115200
rect 321558 109168 321614 109177
rect 321558 109103 321614 109112
rect 321466 97336 321522 97345
rect 321466 97271 321522 97280
rect 321480 96626 321508 97271
rect 321468 96620 321520 96626
rect 321468 96562 321520 96568
rect 314660 95940 314712 95946
rect 314660 95882 314712 95888
rect 311164 90364 311216 90370
rect 311164 90306 311216 90312
rect 310520 89004 310572 89010
rect 310520 88946 310572 88952
rect 310428 80028 310480 80034
rect 310428 79970 310480 79976
rect 310440 79354 310468 79970
rect 310428 79348 310480 79354
rect 310428 79290 310480 79296
rect 309876 32428 309928 32434
rect 309876 32370 309928 32376
rect 310532 16574 310560 88946
rect 310532 16546 311112 16574
rect 309876 8220 309928 8226
rect 309876 8162 309928 8168
rect 309888 7614 309916 8162
rect 309232 7608 309284 7614
rect 309232 7550 309284 7556
rect 309876 7608 309928 7614
rect 309876 7550 309928 7556
rect 309152 6886 309824 6914
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 309060 480 309088 3538
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 6886
rect 311084 3482 311112 16546
rect 311176 3602 311204 90306
rect 312544 86284 312596 86290
rect 312544 86226 312596 86232
rect 312556 27606 312584 86226
rect 313738 84824 313794 84833
rect 313738 84759 313794 84768
rect 313752 84182 313780 84759
rect 313740 84176 313792 84182
rect 313740 84118 313792 84124
rect 313752 82890 313780 84118
rect 313280 82884 313332 82890
rect 313280 82826 313332 82832
rect 313740 82884 313792 82890
rect 313740 82826 313792 82832
rect 311900 27600 311952 27606
rect 311900 27542 311952 27548
rect 312544 27600 312596 27606
rect 312544 27542 312596 27548
rect 311912 16574 311940 27542
rect 313292 16574 313320 82826
rect 314672 22098 314700 95882
rect 317420 94512 317472 94518
rect 317420 94454 317472 94460
rect 316038 91760 316094 91769
rect 316038 91695 316094 91704
rect 316052 88262 316080 91695
rect 316040 88256 316092 88262
rect 316040 88198 316092 88204
rect 315304 67040 315356 67046
rect 315304 66982 315356 66988
rect 314660 22092 314712 22098
rect 314660 22034 314712 22040
rect 314672 21486 314700 22034
rect 314660 21480 314712 21486
rect 314660 21422 314712 21428
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 311164 3596 311216 3602
rect 311164 3538 311216 3544
rect 311084 3454 311480 3482
rect 311452 480 311480 3454
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 315316 3534 315344 66982
rect 316052 3602 316080 88198
rect 317432 16574 317460 94454
rect 318800 93152 318852 93158
rect 318800 93094 318852 93100
rect 317512 90432 317564 90438
rect 317512 90374 317564 90380
rect 317524 28966 317552 90374
rect 317512 28960 317564 28966
rect 317512 28902 317564 28908
rect 318708 28960 318760 28966
rect 318708 28902 318760 28908
rect 318720 27674 318748 28902
rect 318708 27668 318760 27674
rect 318708 27610 318760 27616
rect 318812 16574 318840 93094
rect 321572 92478 321600 109103
rect 323308 107636 323360 107642
rect 323308 107578 323360 107584
rect 323320 106321 323348 107578
rect 322938 106312 322994 106321
rect 322938 106247 322994 106256
rect 323306 106312 323362 106321
rect 323306 106247 323362 106256
rect 321652 103488 321704 103494
rect 321652 103430 321704 103436
rect 321664 102785 321692 103430
rect 321650 102776 321706 102785
rect 321650 102711 321706 102720
rect 321664 95130 321692 102711
rect 321742 101144 321798 101153
rect 321742 101079 321798 101088
rect 321652 95124 321704 95130
rect 321652 95066 321704 95072
rect 321756 93838 321784 101079
rect 322952 95198 322980 106247
rect 322940 95192 322992 95198
rect 322940 95134 322992 95140
rect 321744 93832 321796 93838
rect 321744 93774 321796 93780
rect 321560 92472 321612 92478
rect 321560 92414 321612 92420
rect 320824 86352 320876 86358
rect 320824 86294 320876 86300
rect 320836 31754 320864 86294
rect 323596 75274 323624 115194
rect 324320 114504 324372 114510
rect 324320 114446 324372 114452
rect 324332 114073 324360 114446
rect 324412 114436 324464 114442
rect 324412 114378 324464 114384
rect 324318 114064 324374 114073
rect 324318 113999 324374 114008
rect 324424 113257 324452 114378
rect 324410 113248 324466 113257
rect 324410 113183 324466 113192
rect 324976 110945 325004 115262
rect 324962 110936 325018 110945
rect 324962 110871 325018 110880
rect 324320 110424 324372 110430
rect 324320 110366 324372 110372
rect 324332 110129 324360 110366
rect 324318 110120 324374 110129
rect 324318 110055 324374 110064
rect 324412 108996 324464 109002
rect 324412 108938 324464 108944
rect 324320 108928 324372 108934
rect 324320 108870 324372 108876
rect 324332 108361 324360 108870
rect 324424 108633 324452 108938
rect 324410 108624 324466 108633
rect 324410 108559 324466 108568
rect 324318 108352 324374 108361
rect 324318 108287 324374 108296
rect 325068 107137 325096 119342
rect 326342 112432 326398 112441
rect 326342 112367 326398 112376
rect 325054 107128 325110 107137
rect 325054 107063 325110 107072
rect 324320 106276 324372 106282
rect 324320 106218 324372 106224
rect 324332 105505 324360 106218
rect 324318 105496 324374 105505
rect 324318 105431 324374 105440
rect 324320 104848 324372 104854
rect 324320 104790 324372 104796
rect 324502 104816 324558 104825
rect 324332 104009 324360 104790
rect 324502 104751 324558 104760
rect 324516 104174 324544 104751
rect 324504 104168 324556 104174
rect 324504 104110 324556 104116
rect 324318 104000 324374 104009
rect 324318 103935 324374 103944
rect 324318 102504 324374 102513
rect 324318 102439 324374 102448
rect 324332 102134 324360 102439
rect 324320 102128 324372 102134
rect 324320 102070 324372 102076
rect 324412 102060 324464 102066
rect 324412 102002 324464 102008
rect 324424 100881 324452 102002
rect 324410 100872 324466 100881
rect 324410 100807 324466 100816
rect 324320 100700 324372 100706
rect 324320 100642 324372 100648
rect 324332 100201 324360 100642
rect 324318 100192 324374 100201
rect 324318 100127 324374 100136
rect 324410 99376 324466 99385
rect 324410 99311 324466 99320
rect 324318 97064 324374 97073
rect 324318 96999 324374 97008
rect 324332 92449 324360 96999
rect 324424 93673 324452 99311
rect 324516 93809 324544 104110
rect 326356 95062 326384 112367
rect 327080 101448 327132 101454
rect 327080 101390 327132 101396
rect 325700 95056 325752 95062
rect 325700 94998 325752 95004
rect 326344 95056 326396 95062
rect 326344 94998 326396 95004
rect 324502 93800 324558 93809
rect 324502 93735 324558 93744
rect 324410 93664 324466 93673
rect 324410 93599 324466 93608
rect 324318 92440 324374 92449
rect 324318 92375 324374 92384
rect 323584 75268 323636 75274
rect 323584 75210 323636 75216
rect 324964 66904 325016 66910
rect 324964 66846 325016 66852
rect 322940 40792 322992 40798
rect 322940 40734 322992 40740
rect 320824 31748 320876 31754
rect 320824 31690 320876 31696
rect 320836 31278 320864 31690
rect 320180 31272 320232 31278
rect 320180 31214 320232 31220
rect 320824 31272 320876 31278
rect 320824 31214 320876 31220
rect 320192 16574 320220 31214
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 316040 3596 316092 3602
rect 316040 3538 316092 3544
rect 317328 3596 317380 3602
rect 317328 3538 317380 3544
rect 315028 3528 315080 3534
rect 315028 3470 315080 3476
rect 315304 3528 315356 3534
rect 315304 3470 315356 3476
rect 316224 3528 316276 3534
rect 316224 3470 316276 3476
rect 315040 480 315068 3470
rect 316236 480 316264 3470
rect 317340 480 317368 3538
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322112 3596 322164 3602
rect 322112 3538 322164 3544
rect 322124 480 322152 3538
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 40734
rect 324976 38622 325004 66846
rect 324320 38616 324372 38622
rect 324320 38558 324372 38564
rect 324964 38616 325016 38622
rect 324964 38558 325016 38564
rect 324332 3398 324360 38558
rect 324964 32428 325016 32434
rect 324964 32370 325016 32376
rect 324976 6866 325004 32370
rect 325712 16574 325740 94998
rect 327092 16574 327120 101390
rect 325712 16546 326384 16574
rect 327092 16546 327672 16574
rect 324964 6860 325016 6866
rect 324964 6802 325016 6808
rect 324976 5574 325004 6802
rect 324412 5568 324464 5574
rect 324412 5510 324464 5516
rect 324964 5568 325016 5574
rect 324964 5510 325016 5516
rect 324320 3392 324372 3398
rect 324320 3334 324372 3340
rect 324424 480 324452 5510
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 327080 7608 327132 7614
rect 327080 7550 327132 7556
rect 327092 3602 327120 7550
rect 327080 3596 327132 3602
rect 327080 3538 327132 3544
rect 327644 3482 327672 16546
rect 327736 3602 327764 146882
rect 327828 143614 327856 168370
rect 328564 144838 328592 222022
rect 328552 144832 328604 144838
rect 328552 144774 328604 144780
rect 327816 143608 327868 143614
rect 327816 143550 327868 143556
rect 329116 104174 329144 528906
rect 329288 474156 329340 474162
rect 329288 474098 329340 474104
rect 329196 438932 329248 438938
rect 329196 438874 329248 438880
rect 329208 222086 329236 438874
rect 329300 405686 329328 474098
rect 329288 405680 329340 405686
rect 329288 405622 329340 405628
rect 329760 392834 329788 576846
rect 331048 572694 331076 596226
rect 331036 572688 331088 572694
rect 331036 572630 331088 572636
rect 330576 510672 330628 510678
rect 330576 510614 330628 510620
rect 330484 454096 330536 454102
rect 330484 454038 330536 454044
rect 329748 392828 329800 392834
rect 329748 392770 329800 392776
rect 329196 222080 329248 222086
rect 329196 222022 329248 222028
rect 329840 197736 329892 197742
rect 329840 197678 329892 197684
rect 329196 177404 329248 177410
rect 329196 177346 329248 177352
rect 329208 153270 329236 177346
rect 329196 153264 329248 153270
rect 329196 153206 329248 153212
rect 329208 151814 329236 153206
rect 329208 151786 329328 151814
rect 329196 144968 329248 144974
rect 329196 144910 329248 144916
rect 329104 104168 329156 104174
rect 329104 104110 329156 104116
rect 328460 86352 328512 86358
rect 328460 86294 328512 86300
rect 328472 16574 328500 86294
rect 328472 16546 328776 16574
rect 327724 3596 327776 3602
rect 327724 3538 327776 3544
rect 327644 3454 328040 3482
rect 328012 480 328040 3454
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 329208 4146 329236 144910
rect 329300 43518 329328 151786
rect 329852 128246 329880 197678
rect 330024 183116 330076 183122
rect 330024 183058 330076 183064
rect 329932 177540 329984 177546
rect 329932 177482 329984 177488
rect 329944 148986 329972 177482
rect 330036 158642 330064 183058
rect 330024 158636 330076 158642
rect 330024 158578 330076 158584
rect 329932 148980 329984 148986
rect 329932 148922 329984 148928
rect 330496 137902 330524 454038
rect 330588 198694 330616 510614
rect 331140 396817 331168 601695
rect 331864 599344 331916 599350
rect 331864 599286 331916 599292
rect 331876 482322 331904 599286
rect 331956 594856 332008 594862
rect 331956 594798 332008 594804
rect 331968 549234 331996 594798
rect 331956 549228 332008 549234
rect 331956 549170 332008 549176
rect 331864 482316 331916 482322
rect 331864 482258 331916 482264
rect 331956 467492 332008 467498
rect 331956 467434 332008 467440
rect 331864 456816 331916 456822
rect 331864 456758 331916 456764
rect 331220 398132 331272 398138
rect 331220 398074 331272 398080
rect 331126 396808 331182 396817
rect 331126 396743 331182 396752
rect 330576 198688 330628 198694
rect 330576 198630 330628 198636
rect 330588 197742 330616 198630
rect 330576 197736 330628 197742
rect 330576 197678 330628 197684
rect 331232 164218 331260 398074
rect 331312 397248 331364 397254
rect 331312 397190 331364 397196
rect 331324 396846 331352 397190
rect 331312 396840 331364 396846
rect 331312 396782 331364 396788
rect 331312 234592 331364 234598
rect 331312 234534 331364 234540
rect 331324 234462 331352 234534
rect 331312 234456 331364 234462
rect 331312 234398 331364 234404
rect 331876 219434 331904 456758
rect 331968 398138 331996 467434
rect 331956 398132 332008 398138
rect 331956 398074 332008 398080
rect 332428 396846 332456 700266
rect 348804 699718 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 359464 700392 359516 700398
rect 359464 700334 359516 700340
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 351184 699712 351236 699718
rect 351184 699654 351236 699660
rect 348804 698970 348832 699654
rect 348792 698964 348844 698970
rect 348792 698906 348844 698912
rect 338764 643136 338816 643142
rect 338764 643078 338816 643084
rect 337936 630692 337988 630698
rect 337936 630634 337988 630640
rect 333336 606008 333388 606014
rect 333336 605950 333388 605956
rect 332508 604784 332560 604790
rect 332508 604726 332560 604732
rect 332416 396840 332468 396846
rect 332416 396782 332468 396788
rect 332520 234598 332548 604726
rect 333244 585200 333296 585206
rect 333244 585142 333296 585148
rect 332598 236056 332654 236065
rect 332598 235991 332654 236000
rect 332508 234592 332560 234598
rect 332508 234534 332560 234540
rect 331864 219428 331916 219434
rect 331864 219370 331916 219376
rect 331876 218822 331904 219370
rect 331312 218816 331364 218822
rect 331312 218758 331364 218764
rect 331864 218816 331916 218822
rect 331864 218758 331916 218764
rect 331220 164212 331272 164218
rect 331220 164154 331272 164160
rect 331324 146198 331352 218758
rect 331402 198792 331458 198801
rect 331402 198727 331458 198736
rect 331312 146192 331364 146198
rect 331312 146134 331364 146140
rect 331416 143546 331444 198727
rect 331496 178084 331548 178090
rect 331496 178026 331548 178032
rect 331508 144906 331536 178026
rect 332416 163532 332468 163538
rect 332416 163474 332468 163480
rect 332428 160070 332456 163474
rect 332416 160064 332468 160070
rect 332416 160006 332468 160012
rect 331864 146396 331916 146402
rect 331864 146338 331916 146344
rect 331496 144900 331548 144906
rect 331496 144842 331548 144848
rect 331404 143540 331456 143546
rect 331404 143482 331456 143488
rect 330484 137896 330536 137902
rect 330484 137838 330536 137844
rect 329840 128240 329892 128246
rect 329840 128182 329892 128188
rect 329288 43512 329340 43518
rect 329288 43454 329340 43460
rect 329840 37936 329892 37942
rect 329840 37878 329892 37884
rect 329852 16574 329880 37878
rect 331220 23452 331272 23458
rect 331220 23394 331272 23400
rect 331232 22982 331260 23394
rect 331220 22976 331272 22982
rect 331220 22918 331272 22924
rect 329852 16546 330432 16574
rect 329196 4140 329248 4146
rect 329196 4082 329248 4088
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 22918
rect 331876 3670 331904 146338
rect 331956 142180 332008 142186
rect 331956 142122 332008 142128
rect 331968 33930 331996 142122
rect 332612 115326 332640 235991
rect 333256 197305 333284 585142
rect 333348 566506 333376 605950
rect 336094 601896 336150 601905
rect 336094 601831 336150 601840
rect 334808 600568 334860 600574
rect 334808 600510 334860 600516
rect 334716 599072 334768 599078
rect 334716 599014 334768 599020
rect 333428 597848 333480 597854
rect 333428 597790 333480 597796
rect 333336 566500 333388 566506
rect 333336 566442 333388 566448
rect 333336 495508 333388 495514
rect 333336 495450 333388 495456
rect 333348 237289 333376 495450
rect 333440 388482 333468 597790
rect 334622 595096 334678 595105
rect 334622 595031 334678 595040
rect 333980 405680 334032 405686
rect 333980 405622 334032 405628
rect 333992 404394 334020 405622
rect 333980 404388 334032 404394
rect 333980 404330 334032 404336
rect 333428 388476 333480 388482
rect 333428 388418 333480 388424
rect 333334 237280 333390 237289
rect 333334 237215 333390 237224
rect 333348 236065 333376 237215
rect 333334 236056 333390 236065
rect 333334 235991 333390 236000
rect 333980 215552 334032 215558
rect 333980 215494 334032 215500
rect 333242 197296 333298 197305
rect 333242 197231 333298 197240
rect 333256 196081 333284 197231
rect 333242 196072 333298 196081
rect 333242 196007 333298 196016
rect 332692 187196 332744 187202
rect 332692 187138 332744 187144
rect 332704 135182 332732 187138
rect 332782 181520 332838 181529
rect 332782 181455 332838 181464
rect 332796 142118 332824 181455
rect 332876 177472 332928 177478
rect 332876 177414 332928 177420
rect 332888 157350 332916 177414
rect 332876 157344 332928 157350
rect 332876 157286 332928 157292
rect 332784 142112 332836 142118
rect 332784 142054 332836 142060
rect 332692 135176 332744 135182
rect 332692 135118 332744 135124
rect 333992 119406 334020 215494
rect 334636 206961 334664 595031
rect 334728 534070 334756 599014
rect 334820 559570 334848 600510
rect 336002 597680 336058 597689
rect 336002 597615 336058 597624
rect 334808 559564 334860 559570
rect 334808 559506 334860 559512
rect 334716 534064 334768 534070
rect 334716 534006 334768 534012
rect 336016 528562 336044 597615
rect 336108 580990 336136 601831
rect 336648 600636 336700 600642
rect 336648 600578 336700 600584
rect 336554 594552 336610 594561
rect 336554 594487 336610 594496
rect 336568 589966 336596 594487
rect 336556 589960 336608 589966
rect 336556 589902 336608 589908
rect 336096 580984 336148 580990
rect 336096 580926 336148 580932
rect 336004 528556 336056 528562
rect 336004 528498 336056 528504
rect 336004 518968 336056 518974
rect 336004 518910 336056 518916
rect 335268 459604 335320 459610
rect 335268 459546 335320 459552
rect 335176 407176 335228 407182
rect 335176 407118 335228 407124
rect 334808 404388 334860 404394
rect 334808 404330 334860 404336
rect 334716 222964 334768 222970
rect 334716 222906 334768 222912
rect 334622 206952 334678 206961
rect 334622 206887 334678 206896
rect 334636 205737 334664 206887
rect 334622 205728 334678 205737
rect 334622 205663 334678 205672
rect 334164 184204 334216 184210
rect 334164 184146 334216 184152
rect 334072 178696 334124 178702
rect 334072 178638 334124 178644
rect 334084 158710 334112 178638
rect 334176 168434 334204 184146
rect 334164 168428 334216 168434
rect 334164 168370 334216 168376
rect 334072 158704 334124 158710
rect 334072 158646 334124 158652
rect 333980 119400 334032 119406
rect 333980 119342 334032 119348
rect 332600 115320 332652 115326
rect 332600 115262 332652 115268
rect 332600 98660 332652 98666
rect 332600 98602 332652 98608
rect 332046 84824 332102 84833
rect 332046 84759 332102 84768
rect 331956 33924 332008 33930
rect 331956 33866 332008 33872
rect 332060 22982 332088 84759
rect 332048 22976 332100 22982
rect 332048 22918 332100 22924
rect 331864 3664 331916 3670
rect 331864 3606 331916 3612
rect 332612 3534 332640 98602
rect 334728 77314 334756 222906
rect 334820 216578 334848 404330
rect 335188 394602 335216 407118
rect 335280 396914 335308 459546
rect 335360 408536 335412 408542
rect 335360 408478 335412 408484
rect 335372 405686 335400 408478
rect 335360 405680 335412 405686
rect 335360 405622 335412 405628
rect 335372 402974 335400 405622
rect 335372 402946 335492 402974
rect 335268 396908 335320 396914
rect 335268 396850 335320 396856
rect 335176 394596 335228 394602
rect 335176 394538 335228 394544
rect 335360 393984 335412 393990
rect 335360 393926 335412 393932
rect 334808 216572 334860 216578
rect 334808 216514 334860 216520
rect 334820 215558 334848 216514
rect 334808 215552 334860 215558
rect 334808 215494 334860 215500
rect 335372 102066 335400 393926
rect 335464 211138 335492 402946
rect 336016 398546 336044 518910
rect 336096 443148 336148 443154
rect 336096 443090 336148 443096
rect 336004 398540 336056 398546
rect 336004 398482 336056 398488
rect 336108 393990 336136 443090
rect 336096 393984 336148 393990
rect 336096 393926 336148 393932
rect 336660 363730 336688 600578
rect 337844 594992 337896 594998
rect 337844 594934 337896 594940
rect 337106 591832 337162 591841
rect 337106 591767 337162 591776
rect 337120 587178 337148 591767
rect 337658 589112 337714 589121
rect 337658 589047 337714 589056
rect 337672 587926 337700 589047
rect 337660 587920 337712 587926
rect 337660 587862 337712 587868
rect 337108 587172 337160 587178
rect 337108 587114 337160 587120
rect 337658 586392 337714 586401
rect 337658 586327 337714 586336
rect 337672 585206 337700 586327
rect 337660 585200 337712 585206
rect 337660 585142 337712 585148
rect 337658 584352 337714 584361
rect 337658 584287 337714 584296
rect 337672 583778 337700 584287
rect 337660 583772 337712 583778
rect 337660 583714 337712 583720
rect 337658 581632 337714 581641
rect 337658 581567 337714 581576
rect 337672 581058 337700 581567
rect 337660 581052 337712 581058
rect 337660 580994 337712 581000
rect 337658 578912 337714 578921
rect 337658 578847 337714 578856
rect 337672 578270 337700 578847
rect 337660 578264 337712 578270
rect 337660 578206 337712 578212
rect 337660 576904 337712 576910
rect 337658 576872 337660 576881
rect 337712 576872 337714 576881
rect 337658 576807 337714 576816
rect 337856 574161 337884 594934
rect 337842 574152 337898 574161
rect 337842 574087 337898 574096
rect 337660 572688 337712 572694
rect 337660 572630 337712 572636
rect 337672 571441 337700 572630
rect 337658 571432 337714 571441
rect 337658 571367 337714 571376
rect 337844 570580 337896 570586
rect 337844 570522 337896 570528
rect 337658 568712 337714 568721
rect 337658 568647 337660 568656
rect 337712 568647 337714 568656
rect 337660 568618 337712 568624
rect 337384 561740 337436 561746
rect 337384 561682 337436 561688
rect 336924 560244 336976 560250
rect 336924 560186 336976 560192
rect 336936 559201 336964 560186
rect 336922 559192 336978 559201
rect 336922 559127 336978 559136
rect 337396 553761 337424 561682
rect 337658 561232 337714 561241
rect 337658 561167 337714 561176
rect 337672 560318 337700 561167
rect 337660 560312 337712 560318
rect 337660 560254 337712 560260
rect 337382 553752 337438 553761
rect 337382 553687 337438 553696
rect 337382 551032 337438 551041
rect 337382 550967 337438 550976
rect 337396 546553 337424 550967
rect 337658 548992 337714 549001
rect 337658 548927 337714 548936
rect 337672 547942 337700 548927
rect 337660 547936 337712 547942
rect 337660 547878 337712 547884
rect 337382 546544 337438 546553
rect 337382 546479 337438 546488
rect 337382 546272 337438 546281
rect 337382 546207 337438 546216
rect 337292 536784 337344 536790
rect 337292 536726 337344 536732
rect 337304 536081 337332 536726
rect 337290 536072 337346 536081
rect 337290 536007 337346 536016
rect 336832 532024 336884 532030
rect 336832 531966 336884 531972
rect 336844 531321 336872 531966
rect 336830 531312 336886 531321
rect 336830 531247 336886 531256
rect 336844 528970 336872 531247
rect 336832 528964 336884 528970
rect 336832 528906 336884 528912
rect 337396 525094 337424 546207
rect 337658 543552 337714 543561
rect 337658 543487 337714 543496
rect 337672 542434 337700 543487
rect 337660 542428 337712 542434
rect 337660 542370 337712 542376
rect 337474 541512 337530 541521
rect 337474 541447 337530 541456
rect 337488 541006 337516 541447
rect 337476 541000 337528 541006
rect 337476 540942 337528 540948
rect 337660 539572 337712 539578
rect 337660 539514 337712 539520
rect 337672 538801 337700 539514
rect 337658 538792 337714 538801
rect 337658 538727 337714 538736
rect 337658 533352 337714 533361
rect 337658 533287 337714 533296
rect 337672 532778 337700 533287
rect 337660 532772 337712 532778
rect 337660 532714 337712 532720
rect 337856 526454 337884 570522
rect 337948 556850 337976 630634
rect 338028 613420 338080 613426
rect 338028 613362 338080 613368
rect 337936 556844 337988 556850
rect 337936 556786 337988 556792
rect 337948 556481 337976 556786
rect 337934 556472 337990 556481
rect 337934 556407 337990 556416
rect 337844 526448 337896 526454
rect 337844 526390 337896 526396
rect 337856 525881 337884 526390
rect 337842 525872 337898 525881
rect 337842 525807 337898 525816
rect 337384 525088 337436 525094
rect 337384 525030 337436 525036
rect 337474 523832 337530 523841
rect 337474 523767 337530 523776
rect 337488 523054 337516 523767
rect 337476 523048 337528 523054
rect 337476 522990 337528 522996
rect 337474 521112 337530 521121
rect 337474 521047 337530 521056
rect 337488 520334 337516 521047
rect 337476 520328 337528 520334
rect 337476 520270 337528 520276
rect 337658 515672 337714 515681
rect 337658 515607 337714 515616
rect 337672 514826 337700 515607
rect 337660 514820 337712 514826
rect 337660 514762 337712 514768
rect 337658 513632 337714 513641
rect 337658 513567 337714 513576
rect 337672 513398 337700 513567
rect 337660 513392 337712 513398
rect 337660 513334 337712 513340
rect 337658 510912 337714 510921
rect 337658 510847 337714 510856
rect 337672 510678 337700 510847
rect 337660 510672 337712 510678
rect 337660 510614 337712 510620
rect 337106 506152 337162 506161
rect 337106 506087 337162 506096
rect 337120 505170 337148 506087
rect 337108 505164 337160 505170
rect 337108 505106 337160 505112
rect 337752 503736 337804 503742
rect 337752 503678 337804 503684
rect 337658 503432 337714 503441
rect 337658 503367 337714 503376
rect 337672 502382 337700 503367
rect 337660 502376 337712 502382
rect 337660 502318 337712 502324
rect 337764 500721 337792 503678
rect 337750 500712 337806 500721
rect 337750 500647 337806 500656
rect 337658 497992 337714 498001
rect 337658 497927 337714 497936
rect 337672 496874 337700 497927
rect 337660 496868 337712 496874
rect 337660 496810 337712 496816
rect 337474 495952 337530 495961
rect 337474 495887 337530 495896
rect 337488 495514 337516 495887
rect 337476 495508 337528 495514
rect 337476 495450 337528 495456
rect 337474 493232 337530 493241
rect 337474 493167 337530 493176
rect 337488 491366 337516 493167
rect 337476 491360 337528 491366
rect 337476 491302 337528 491308
rect 337658 490512 337714 490521
rect 337658 490447 337714 490456
rect 337672 489938 337700 490447
rect 337660 489932 337712 489938
rect 337660 489874 337712 489880
rect 337750 485752 337806 485761
rect 337750 485687 337806 485696
rect 337764 485110 337792 485687
rect 337752 485104 337804 485110
rect 337752 485046 337804 485052
rect 336738 480312 336794 480321
rect 336738 480247 336794 480256
rect 337764 480254 337792 485046
rect 337936 484356 337988 484362
rect 337936 484298 337988 484304
rect 337948 483041 337976 484298
rect 337934 483032 337990 483041
rect 337934 482967 337990 482976
rect 336752 479534 336780 480247
rect 337764 480226 337976 480254
rect 336740 479528 336792 479534
rect 336740 479470 336792 479476
rect 337750 478272 337806 478281
rect 337750 478207 337806 478216
rect 337658 475552 337714 475561
rect 337658 475487 337714 475496
rect 337672 474774 337700 475487
rect 337660 474768 337712 474774
rect 337660 474710 337712 474716
rect 337764 474162 337792 478207
rect 337752 474156 337804 474162
rect 337752 474098 337804 474104
rect 336830 472832 336886 472841
rect 336830 472767 336886 472776
rect 336738 470792 336794 470801
rect 336738 470727 336794 470736
rect 336752 469878 336780 470727
rect 336740 469872 336792 469878
rect 336740 469814 336792 469820
rect 336844 467498 336872 472767
rect 336832 467492 336884 467498
rect 336832 467434 336884 467440
rect 337658 465352 337714 465361
rect 337658 465287 337714 465296
rect 337672 461650 337700 465287
rect 337660 461644 337712 461650
rect 337660 461586 337712 461592
rect 337658 460592 337714 460601
rect 337658 460527 337714 460536
rect 337672 459610 337700 460527
rect 337660 459604 337712 459610
rect 337660 459546 337712 459552
rect 337658 457872 337714 457881
rect 337658 457807 337714 457816
rect 337672 456822 337700 457807
rect 337660 456816 337712 456822
rect 337660 456758 337712 456764
rect 337658 455152 337714 455161
rect 337658 455087 337714 455096
rect 337672 454102 337700 455087
rect 337660 454096 337712 454102
rect 337660 454038 337712 454044
rect 337566 453112 337622 453121
rect 337566 453047 337622 453056
rect 337580 451926 337608 453047
rect 337568 451920 337620 451926
rect 337568 451862 337620 451868
rect 337290 450392 337346 450401
rect 337290 450327 337346 450336
rect 337304 449954 337332 450327
rect 337292 449948 337344 449954
rect 337292 449890 337344 449896
rect 337106 447672 337162 447681
rect 337106 447607 337162 447616
rect 337120 446418 337148 447607
rect 337108 446412 337160 446418
rect 337108 446354 337160 446360
rect 337290 440192 337346 440201
rect 337290 440127 337346 440136
rect 337304 438938 337332 440127
rect 337292 438932 337344 438938
rect 337292 438874 337344 438880
rect 337290 437472 337346 437481
rect 337290 437407 337346 437416
rect 337304 436150 337332 437407
rect 337292 436144 337344 436150
rect 337292 436086 337344 436092
rect 337382 435432 337438 435441
rect 337382 435367 337438 435376
rect 337396 431254 337424 435367
rect 337658 432712 337714 432721
rect 337658 432647 337714 432656
rect 337672 432002 337700 432647
rect 337660 431996 337712 432002
rect 337660 431938 337712 431944
rect 337384 431248 337436 431254
rect 337384 431190 337436 431196
rect 336922 429992 336978 430001
rect 336922 429927 336978 429936
rect 336936 429214 336964 429927
rect 336924 429208 336976 429214
rect 336924 429150 336976 429156
rect 336922 427272 336978 427281
rect 336922 427207 336978 427216
rect 336936 426494 336964 427207
rect 336924 426488 336976 426494
rect 336924 426430 336976 426436
rect 337658 425232 337714 425241
rect 337658 425167 337714 425176
rect 337672 425134 337700 425167
rect 337660 425128 337712 425134
rect 337660 425070 337712 425076
rect 337658 422512 337714 422521
rect 337658 422447 337714 422456
rect 337672 422346 337700 422447
rect 337660 422340 337712 422346
rect 337660 422282 337712 422288
rect 337842 417752 337898 417761
rect 337842 417687 337898 417696
rect 336832 415404 336884 415410
rect 336832 415346 336884 415352
rect 336844 415041 336872 415346
rect 336830 415032 336886 415041
rect 336830 414967 336886 414976
rect 337382 412312 337438 412321
rect 337382 412247 337438 412256
rect 336922 409592 336978 409601
rect 336922 409527 336978 409536
rect 336936 408542 336964 409527
rect 336924 408536 336976 408542
rect 336924 408478 336976 408484
rect 337396 394058 337424 412247
rect 337476 409896 337528 409902
rect 337476 409838 337528 409844
rect 337488 401713 337516 409838
rect 337658 407552 337714 407561
rect 337658 407487 337714 407496
rect 337672 407182 337700 407487
rect 337660 407176 337712 407182
rect 337660 407118 337712 407124
rect 337750 404832 337806 404841
rect 337750 404767 337806 404776
rect 337764 404394 337792 404767
rect 337752 404388 337804 404394
rect 337752 404330 337804 404336
rect 337474 401704 337530 401713
rect 337474 401639 337530 401648
rect 337384 394052 337436 394058
rect 337384 393994 337436 394000
rect 337856 392630 337884 417687
rect 337948 394534 337976 480226
rect 338040 468518 338068 613362
rect 338776 570586 338804 643078
rect 351196 632738 351224 699654
rect 351184 632732 351236 632738
rect 351184 632674 351236 632680
rect 359476 616758 359504 700334
rect 358084 616752 358136 616758
rect 358084 616694 358136 616700
rect 359464 616752 359516 616758
rect 359464 616694 359516 616700
rect 358096 605198 358124 616694
rect 364352 613426 364380 702406
rect 397472 700398 397500 703520
rect 413664 702846 413692 703520
rect 412640 702840 412692 702846
rect 412640 702782 412692 702788
rect 413652 702840 413704 702846
rect 413652 702782 413704 702788
rect 412652 702506 412680 702782
rect 416780 702704 416832 702710
rect 416780 702646 416832 702652
rect 412640 702500 412692 702506
rect 412640 702442 412692 702448
rect 397460 700392 397512 700398
rect 397460 700334 397512 700340
rect 412652 618934 412680 702442
rect 412640 618928 412692 618934
rect 412640 618870 412692 618876
rect 391020 616888 391072 616894
rect 391020 616830 391072 616836
rect 364340 613420 364392 613426
rect 364340 613362 364392 613368
rect 391032 612882 391060 616830
rect 400864 616140 400916 616146
rect 400864 616082 400916 616088
rect 390560 612876 390612 612882
rect 390560 612818 390612 612824
rect 391020 612876 391072 612882
rect 391020 612818 391072 612824
rect 388536 610156 388588 610162
rect 388536 610098 388588 610104
rect 378876 606144 378928 606150
rect 378876 606086 378928 606092
rect 357440 605192 357492 605198
rect 357440 605134 357492 605140
rect 358084 605192 358136 605198
rect 358084 605134 358136 605140
rect 357452 604722 357480 605134
rect 357440 604716 357492 604722
rect 357440 604658 357492 604664
rect 339040 601928 339092 601934
rect 339040 601870 339092 601876
rect 338946 599040 339002 599049
rect 338946 598975 339002 598984
rect 338856 595060 338908 595066
rect 338856 595002 338908 595008
rect 338764 570580 338816 570586
rect 338764 570522 338816 570528
rect 338762 563952 338818 563961
rect 338762 563887 338818 563896
rect 338028 468512 338080 468518
rect 338028 468454 338080 468460
rect 338040 468081 338068 468454
rect 338026 468072 338082 468081
rect 338026 468007 338082 468016
rect 338026 444952 338082 444961
rect 338026 444887 338082 444896
rect 338040 443154 338068 444887
rect 338028 443148 338080 443154
rect 338028 443090 338080 443096
rect 338580 403640 338632 403646
rect 338580 403582 338632 403588
rect 338026 401704 338082 401713
rect 338026 401639 338082 401648
rect 337936 394528 337988 394534
rect 337936 394470 337988 394476
rect 337844 392624 337896 392630
rect 337844 392566 337896 392572
rect 336648 363724 336700 363730
rect 336648 363666 336700 363672
rect 336660 362982 336688 363666
rect 336648 362976 336700 362982
rect 336648 362918 336700 362924
rect 336740 362228 336792 362234
rect 336740 362170 336792 362176
rect 335452 211132 335504 211138
rect 335452 211074 335504 211080
rect 335464 209774 335492 211074
rect 335464 209746 335584 209774
rect 335452 202360 335504 202366
rect 335452 202302 335504 202308
rect 335464 197266 335492 202302
rect 335452 197260 335504 197266
rect 335452 197202 335504 197208
rect 335464 196081 335492 197202
rect 335450 196072 335506 196081
rect 335450 196007 335506 196016
rect 335452 180328 335504 180334
rect 335452 180270 335504 180276
rect 335464 135250 335492 180270
rect 335452 135244 335504 135250
rect 335452 135186 335504 135192
rect 335556 104854 335584 209746
rect 335634 185600 335690 185609
rect 335634 185535 335690 185544
rect 335648 161430 335676 185535
rect 335636 161424 335688 161430
rect 335636 161366 335688 161372
rect 335636 140072 335688 140078
rect 335636 140014 335688 140020
rect 335544 104848 335596 104854
rect 335544 104790 335596 104796
rect 335360 102060 335412 102066
rect 335360 102002 335412 102008
rect 334716 77308 334768 77314
rect 334716 77250 334768 77256
rect 333242 65512 333298 65521
rect 333242 65447 333298 65456
rect 333256 45529 333284 65447
rect 333242 45520 333298 45529
rect 333242 45455 333298 45464
rect 333256 44305 333284 45455
rect 332690 44296 332746 44305
rect 332690 44231 332746 44240
rect 333242 44296 333298 44305
rect 333242 44231 333298 44240
rect 332600 3528 332652 3534
rect 332600 3470 332652 3476
rect 332704 480 332732 44231
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 333900 480 333928 3470
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334728 354 334756 77250
rect 335648 16574 335676 140014
rect 336752 40730 336780 362170
rect 337384 331288 337436 331294
rect 337384 331230 337436 331236
rect 337396 233170 337424 331230
rect 337936 323604 337988 323610
rect 337936 323546 337988 323552
rect 337948 322998 337976 323546
rect 337936 322992 337988 322998
rect 337936 322934 337988 322940
rect 337384 233164 337436 233170
rect 337384 233106 337436 233112
rect 337384 216028 337436 216034
rect 337384 215970 337436 215976
rect 336832 179376 336884 179382
rect 336832 179318 336884 179324
rect 336844 178809 336872 179318
rect 336830 178800 336886 178809
rect 336830 178735 336886 178744
rect 337292 168224 337344 168230
rect 337292 168166 337344 168172
rect 337304 165578 337332 168166
rect 337292 165572 337344 165578
rect 337292 165514 337344 165520
rect 337396 115258 337424 215970
rect 337948 164898 337976 322934
rect 338040 316742 338068 401639
rect 338592 398614 338620 403582
rect 338580 398608 338632 398614
rect 338580 398550 338632 398556
rect 338776 365906 338804 563887
rect 338868 536110 338896 595002
rect 338960 552702 338988 598975
rect 339052 576162 339080 601870
rect 349896 600432 349948 600438
rect 349896 600374 349948 600380
rect 347964 599344 348016 599350
rect 347964 599286 348016 599292
rect 345480 597848 345532 597854
rect 340326 597816 340382 597825
rect 345480 597790 345532 597796
rect 340326 597751 340382 597760
rect 339684 597712 339736 597718
rect 339684 597654 339736 597660
rect 339500 594788 339552 594794
rect 339500 594730 339552 594736
rect 339512 594114 339540 594730
rect 339500 594108 339552 594114
rect 339500 594050 339552 594056
rect 339696 593366 339724 597654
rect 340340 595354 340368 597751
rect 345492 595354 345520 597790
rect 347976 595354 348004 599286
rect 349908 595354 349936 600374
rect 355138 596456 355194 596465
rect 355138 596391 355194 596400
rect 355152 595354 355180 596391
rect 357452 595354 357480 604658
rect 376760 602064 376812 602070
rect 376760 602006 376812 602012
rect 376772 600370 376800 602006
rect 374000 600364 374052 600370
rect 374000 600306 374052 600312
rect 376760 600364 376812 600370
rect 376760 600306 376812 600312
rect 371792 599276 371844 599282
rect 371792 599218 371844 599224
rect 364798 597952 364854 597961
rect 364798 597887 364854 597896
rect 340340 595326 340676 595354
rect 345492 595326 345828 595354
rect 347976 595326 348404 595354
rect 349908 595326 350336 595354
rect 355152 595326 355488 595354
rect 357420 595326 357480 595354
rect 364812 595354 364840 597887
rect 367100 597780 367152 597786
rect 367100 597722 367152 597728
rect 367112 595354 367140 597722
rect 369308 597644 369360 597650
rect 369308 597586 369360 597592
rect 364812 595326 365148 595354
rect 367080 595326 367140 595354
rect 369320 595354 369348 597586
rect 371804 595354 371832 599218
rect 374012 595354 374040 600306
rect 376772 595354 376800 600306
rect 369320 595326 369656 595354
rect 371804 595326 372232 595354
rect 374012 595326 374164 595354
rect 376740 595326 376800 595354
rect 378888 595354 378916 606086
rect 386420 604648 386472 604654
rect 386420 604590 386472 604596
rect 381452 603152 381504 603158
rect 381452 603094 381504 603100
rect 381464 595354 381492 603094
rect 383660 596352 383712 596358
rect 383660 596294 383712 596300
rect 383672 595354 383700 596294
rect 386432 595354 386460 604590
rect 378888 595326 379316 595354
rect 381464 595326 381892 595354
rect 383672 595326 383824 595354
rect 386400 595326 386460 595354
rect 388548 595354 388576 610098
rect 390572 595354 390600 612818
rect 400876 604790 400904 616082
rect 416792 615494 416820 702646
rect 429856 700330 429884 703520
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 456800 618316 456852 618322
rect 456800 618258 456852 618264
rect 456812 615494 456840 618258
rect 416792 615466 416912 615494
rect 456812 615466 457484 615494
rect 402980 611516 403032 611522
rect 402980 611458 403032 611464
rect 400220 604784 400272 604790
rect 400220 604726 400272 604732
rect 400864 604784 400916 604790
rect 400864 604726 400916 604732
rect 396080 604580 396132 604586
rect 396080 604522 396132 604528
rect 393320 600704 393372 600710
rect 393320 600646 393372 600652
rect 393332 595354 393360 600646
rect 396092 595354 396120 604522
rect 398196 601996 398248 602002
rect 398196 601938 398248 601944
rect 388548 595326 388976 595354
rect 390572 595326 390908 595354
rect 393332 595326 393484 595354
rect 396060 595326 396120 595354
rect 398208 595354 398236 601938
rect 400232 595354 400260 604726
rect 402992 595354 403020 611458
rect 412640 607368 412692 607374
rect 412640 607310 412692 607316
rect 409880 605940 409932 605946
rect 409880 605882 409932 605888
rect 407304 597916 407356 597922
rect 407304 597858 407356 597864
rect 405740 597712 405792 597718
rect 405740 597654 405792 597660
rect 405752 595354 405780 597654
rect 407028 597576 407080 597582
rect 407028 597518 407080 597524
rect 407040 596154 407068 597518
rect 407028 596148 407080 596154
rect 407028 596090 407080 596096
rect 398208 595326 398636 595354
rect 400232 595326 400568 595354
rect 402992 595326 403144 595354
rect 405720 595326 405780 595354
rect 407316 595354 407344 597858
rect 409892 595354 409920 605882
rect 412652 595354 412680 607310
rect 414388 603288 414440 603294
rect 414388 603230 414440 603236
rect 414400 598262 414428 603230
rect 415400 599208 415452 599214
rect 415400 599150 415452 599156
rect 414388 598256 414440 598262
rect 414388 598198 414440 598204
rect 415412 595354 415440 599150
rect 407316 595326 407652 595354
rect 409892 595326 410228 595354
rect 412652 595326 412804 595354
rect 415380 595326 415440 595354
rect 416884 595354 416912 615466
rect 420184 613420 420236 613426
rect 420184 613362 420236 613368
rect 420196 603265 420224 613362
rect 450360 611380 450412 611386
rect 450360 611322 450412 611328
rect 431960 608796 432012 608802
rect 431960 608738 432012 608744
rect 423956 603356 424008 603362
rect 423956 603298 424008 603304
rect 419538 603256 419594 603265
rect 419538 603191 419594 603200
rect 420182 603256 420238 603265
rect 420182 603191 420238 603200
rect 419552 595354 419580 603191
rect 422300 599140 422352 599146
rect 422300 599082 422352 599088
rect 422312 595354 422340 599082
rect 423968 595354 423996 603298
rect 429198 599176 429254 599185
rect 429198 599111 429254 599120
rect 429212 595354 429240 599111
rect 431972 595354 432000 608738
rect 436192 608728 436244 608734
rect 436192 608670 436244 608676
rect 433614 601896 433670 601905
rect 433614 601831 433670 601840
rect 433628 595354 433656 601831
rect 436204 595354 436232 608670
rect 443276 607232 443328 607238
rect 443276 607174 443328 607180
rect 440700 601724 440752 601730
rect 440700 601666 440752 601672
rect 438860 600500 438912 600506
rect 438860 600442 438912 600448
rect 438872 595354 438900 600442
rect 440712 595354 440740 601666
rect 443288 595354 443316 607174
rect 448520 606076 448572 606082
rect 448520 606018 448572 606024
rect 445850 601760 445906 601769
rect 445850 601695 445906 601704
rect 445864 595354 445892 601695
rect 448532 595354 448560 606018
rect 450372 595354 450400 611322
rect 452936 607436 452988 607442
rect 452936 607378 452988 607384
rect 452948 595354 452976 607378
rect 457456 595354 457484 615466
rect 462332 607918 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 613426 477540 702406
rect 494808 700330 494836 703520
rect 527192 702574 527220 703520
rect 538220 702636 538272 702642
rect 538220 702578 538272 702584
rect 527180 702568 527232 702574
rect 527180 702510 527232 702516
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 518164 700324 518216 700330
rect 518164 700266 518216 700272
rect 488540 632732 488592 632738
rect 488540 632674 488592 632680
rect 488552 615494 488580 632674
rect 510620 615528 510672 615534
rect 488552 615466 489040 615494
rect 510620 615470 510672 615476
rect 483848 614236 483900 614242
rect 483848 614178 483900 614184
rect 477500 613420 477552 613426
rect 477500 613362 477552 613368
rect 469680 610020 469732 610026
rect 469680 609962 469732 609968
rect 462320 607912 462372 607918
rect 462320 607854 462372 607860
rect 459560 605872 459612 605878
rect 459560 605814 459612 605820
rect 459572 595542 459600 605814
rect 462594 600536 462650 600545
rect 462594 600471 462650 600480
rect 459560 595536 459612 595542
rect 459560 595478 459612 595484
rect 460434 595536 460486 595542
rect 460434 595478 460486 595484
rect 460446 595354 460474 595478
rect 462608 595354 462636 600471
rect 467194 597816 467250 597825
rect 467194 597751 467250 597760
rect 465264 596556 465316 596562
rect 465264 596498 465316 596504
rect 465276 595354 465304 596498
rect 467208 595354 467236 597751
rect 469692 595354 469720 609962
rect 474188 600636 474240 600642
rect 474188 600578 474240 600584
rect 472992 597712 473044 597718
rect 472992 597654 473044 597660
rect 473004 595354 473032 597654
rect 416884 595326 417312 595354
rect 419552 595326 419888 595354
rect 422312 595326 422464 595354
rect 423968 595326 424396 595354
rect 429212 595326 429548 595354
rect 431972 595326 432124 595354
rect 433628 595326 434056 595354
rect 436204 595326 436632 595354
rect 438872 595326 439208 595354
rect 440712 595326 441140 595354
rect 443288 595326 443716 595354
rect 445864 595326 446292 595354
rect 448532 595326 448868 595354
rect 450372 595326 450800 595354
rect 452948 595326 453376 595354
rect 457456 595326 457884 595354
rect 460446 595340 460612 595354
rect 460460 595326 460612 595340
rect 462608 595326 463036 595354
rect 465276 595326 465612 595354
rect 467208 595326 467544 595354
rect 469692 595326 470120 595354
rect 472696 595326 473032 595354
rect 474200 595354 474228 600578
rect 479338 599040 479394 599049
rect 479338 598975 479394 598984
rect 477408 597780 477460 597786
rect 477408 597722 477460 597728
rect 477420 595354 477448 597722
rect 474200 595326 474628 595354
rect 477204 595326 477448 595354
rect 479352 595354 479380 598975
rect 482008 598256 482060 598262
rect 482008 598198 482060 598204
rect 482020 595354 482048 598198
rect 483860 595354 483888 614178
rect 486884 603220 486936 603226
rect 486884 603162 486936 603168
rect 486896 597650 486924 603162
rect 486884 597644 486936 597650
rect 486884 597586 486936 597592
rect 486896 595354 486924 597586
rect 479352 595326 479780 595354
rect 482020 595326 482356 595354
rect 483860 595326 484288 595354
rect 486864 595326 486924 595354
rect 489012 595354 489040 615466
rect 493508 612808 493560 612814
rect 493508 612750 493560 612756
rect 491300 610088 491352 610094
rect 491300 610030 491352 610036
rect 491312 595490 491340 610030
rect 491312 595462 491386 595490
rect 489012 595326 489440 595354
rect 491358 595340 491386 595462
rect 493520 595354 493548 612750
rect 498660 608660 498712 608666
rect 498660 608602 498712 608608
rect 496084 601928 496136 601934
rect 496084 601870 496136 601876
rect 496096 595354 496124 601870
rect 498672 595354 498700 608602
rect 507858 603120 507914 603129
rect 507858 603055 507914 603064
rect 500960 600568 501012 600574
rect 500960 600510 501012 600516
rect 500972 595490 501000 600510
rect 505742 599040 505798 599049
rect 505742 598975 505798 598984
rect 503628 597848 503680 597854
rect 503628 597790 503680 597796
rect 500972 595462 501046 595490
rect 493520 595326 493948 595354
rect 496096 595326 496524 595354
rect 498672 595326 499100 595354
rect 501018 595340 501046 595462
rect 503640 595354 503668 597790
rect 503608 595326 503668 595354
rect 505756 595354 505784 598975
rect 507872 595354 507900 603055
rect 510632 595490 510660 615470
rect 515402 604480 515458 604489
rect 515402 604415 515458 604424
rect 512828 599140 512880 599146
rect 512828 599082 512880 599088
rect 510632 595462 510706 595490
rect 505756 595326 506184 595354
rect 507872 595326 508116 595354
rect 510678 595340 510706 595462
rect 512840 595354 512868 599082
rect 515416 595354 515444 604415
rect 518176 597922 518204 700266
rect 534356 618928 534408 618934
rect 534356 618870 534408 618876
rect 534264 607912 534316 607918
rect 534264 607854 534316 607860
rect 520280 606008 520332 606014
rect 520280 605950 520332 605956
rect 518164 597916 518216 597922
rect 518164 597858 518216 597864
rect 518176 595354 518204 597858
rect 520292 595490 520320 605950
rect 524420 604512 524472 604518
rect 524420 604454 524472 604460
rect 522946 597816 523002 597825
rect 522946 597751 523002 597760
rect 520292 595462 520366 595490
rect 512840 595326 513268 595354
rect 515416 595326 515844 595354
rect 517776 595326 518204 595354
rect 520338 595340 520366 595462
rect 522960 595354 522988 597751
rect 522928 595326 522988 595354
rect 524432 595354 524460 604454
rect 534080 599004 534132 599010
rect 534080 598946 534132 598952
rect 527180 597576 527232 597582
rect 527180 597518 527232 597524
rect 532608 597576 532660 597582
rect 532608 597518 532660 597524
rect 527192 595354 527220 597518
rect 529940 596216 529992 596222
rect 529940 596158 529992 596164
rect 529952 595490 529980 596158
rect 529952 595462 530026 595490
rect 524432 595326 524860 595354
rect 527192 595326 527436 595354
rect 529998 595340 530026 595462
rect 532620 595354 532648 597518
rect 532588 595326 532648 595354
rect 460584 595134 460612 595326
rect 352564 595128 352616 595134
rect 460572 595128 460624 595134
rect 359646 595096 359702 595105
rect 352616 595076 352912 595082
rect 352564 595070 352912 595076
rect 352576 595054 352912 595070
rect 359702 595054 359996 595082
rect 426636 595066 426972 595082
rect 426624 595060 426972 595066
rect 359646 595031 359702 595040
rect 426676 595054 426972 595060
rect 455952 595066 456288 595082
rect 460572 595070 460624 595076
rect 455952 595060 456300 595066
rect 455952 595054 456248 595060
rect 426624 595002 426676 595008
rect 456248 595002 456300 595008
rect 362222 594960 362278 594969
rect 362278 594918 362572 594946
rect 362222 594895 362278 594904
rect 342916 594794 343252 594810
rect 342904 594788 343252 594794
rect 342956 594782 343252 594788
rect 342904 594730 342956 594736
rect 339684 593360 339736 593366
rect 339684 593302 339736 593308
rect 339040 576156 339092 576162
rect 339040 576098 339092 576104
rect 338948 552696 339000 552702
rect 338948 552638 339000 552644
rect 338856 536104 338908 536110
rect 338856 536046 338908 536052
rect 534092 531321 534120 598946
rect 534170 566672 534226 566681
rect 534170 566607 534226 566616
rect 534078 531312 534134 531321
rect 534078 531247 534134 531256
rect 534078 490512 534134 490521
rect 534078 490447 534134 490456
rect 339314 488472 339370 488481
rect 339314 488407 339370 488416
rect 339328 487218 339356 488407
rect 339316 487212 339368 487218
rect 339316 487154 339368 487160
rect 339132 403708 339184 403714
rect 339132 403650 339184 403656
rect 339144 399634 339172 403650
rect 339132 399628 339184 399634
rect 339132 399570 339184 399576
rect 339328 388482 339356 487154
rect 533434 409592 533490 409601
rect 533356 409550 533434 409578
rect 339868 400920 339920 400926
rect 339868 400862 339920 400868
rect 339500 399832 339552 399838
rect 339500 399774 339552 399780
rect 339512 398886 339540 399774
rect 339500 398880 339552 398886
rect 339406 398848 339462 398857
rect 339500 398822 339552 398828
rect 339406 398783 339462 398792
rect 339316 388476 339368 388482
rect 339316 388418 339368 388424
rect 338764 365900 338816 365906
rect 338764 365842 338816 365848
rect 338028 316736 338080 316742
rect 338028 316678 338080 316684
rect 338120 193860 338172 193866
rect 338120 193802 338172 193808
rect 337936 164892 337988 164898
rect 337936 164834 337988 164840
rect 337474 158808 337530 158817
rect 337474 158743 337530 158752
rect 337488 140758 337516 158743
rect 337476 140752 337528 140758
rect 337476 140694 337528 140700
rect 337476 131776 337528 131782
rect 337476 131718 337528 131724
rect 337384 115252 337436 115258
rect 337384 115194 337436 115200
rect 336832 80708 336884 80714
rect 336832 80650 336884 80656
rect 336844 77314 336872 80650
rect 336832 77308 336884 77314
rect 336832 77250 336884 77256
rect 337488 49026 337516 131718
rect 338132 121378 338160 193802
rect 338304 185700 338356 185706
rect 338304 185642 338356 185648
rect 338212 183048 338264 183054
rect 338212 182990 338264 182996
rect 338224 146946 338252 182990
rect 338316 160750 338344 185642
rect 338304 160744 338356 160750
rect 338304 160686 338356 160692
rect 338776 152522 338804 365842
rect 339420 187066 339448 398783
rect 339408 187060 339460 187066
rect 339408 187002 339460 187008
rect 339512 168230 339540 398822
rect 339880 398478 339908 400862
rect 340018 399838 340046 400044
rect 340006 399832 340058 399838
rect 341950 399786 341978 400044
rect 344526 399786 344554 400044
rect 347102 399786 347130 400044
rect 349034 399838 349062 400044
rect 340006 399774 340058 399780
rect 340984 399758 341978 399786
rect 343744 399758 344554 399786
rect 346412 399758 347130 399786
rect 347872 399832 347924 399838
rect 347872 399774 347924 399780
rect 349022 399832 349074 399838
rect 351610 399786 351638 400044
rect 354186 399922 354214 400044
rect 349022 399774 349074 399780
rect 339868 398472 339920 398478
rect 339868 398414 339920 398420
rect 340984 382974 341012 399758
rect 343638 396808 343694 396817
rect 341524 396772 341576 396778
rect 343638 396743 343694 396752
rect 341524 396714 341576 396720
rect 340972 382968 341024 382974
rect 340972 382910 341024 382916
rect 340880 362976 340932 362982
rect 340880 362918 340932 362924
rect 340142 362808 340198 362817
rect 340142 362743 340198 362752
rect 340156 362273 340184 362743
rect 340142 362264 340198 362273
rect 340142 362199 340198 362208
rect 340156 361758 340184 362199
rect 340144 361752 340196 361758
rect 340144 361694 340196 361700
rect 339684 182912 339736 182918
rect 339684 182854 339736 182860
rect 339592 182232 339644 182238
rect 339592 182174 339644 182180
rect 339500 168224 339552 168230
rect 339500 168166 339552 168172
rect 338764 152516 338816 152522
rect 338764 152458 338816 152464
rect 339408 147620 339460 147626
rect 339408 147562 339460 147568
rect 339420 146946 339448 147562
rect 338212 146940 338264 146946
rect 338212 146882 338264 146888
rect 339408 146940 339460 146946
rect 339408 146882 339460 146888
rect 339604 131034 339632 182174
rect 339696 153202 339724 182854
rect 340144 173188 340196 173194
rect 340144 173130 340196 173136
rect 339684 153196 339736 153202
rect 339684 153138 339736 153144
rect 339592 131028 339644 131034
rect 339592 130970 339644 130976
rect 338212 123480 338264 123486
rect 338212 123422 338264 123428
rect 338120 121372 338172 121378
rect 338120 121314 338172 121320
rect 337476 49020 337528 49026
rect 337476 48962 337528 48968
rect 337476 42220 337528 42226
rect 337476 42162 337528 42168
rect 336740 40724 336792 40730
rect 336740 40666 336792 40672
rect 337488 33114 337516 42162
rect 338028 41336 338080 41342
rect 338028 41278 338080 41284
rect 338040 40730 338068 41278
rect 338028 40724 338080 40730
rect 338028 40666 338080 40672
rect 337476 33108 337528 33114
rect 337476 33050 337528 33056
rect 337488 31822 337516 33050
rect 336740 31816 336792 31822
rect 336740 31758 336792 31764
rect 337476 31816 337528 31822
rect 337476 31758 337528 31764
rect 336004 31204 336056 31210
rect 336004 31146 336056 31152
rect 335648 16546 335952 16574
rect 335924 3482 335952 16546
rect 336016 3602 336044 31146
rect 336752 16574 336780 31758
rect 336832 26240 336884 26246
rect 336830 26208 336832 26217
rect 336884 26208 336886 26217
rect 336830 26143 336886 26152
rect 336844 25537 336872 26143
rect 336830 25528 336886 25537
rect 336830 25463 336886 25472
rect 338224 16574 338252 123422
rect 340156 108934 340184 173130
rect 340144 108928 340196 108934
rect 340144 108870 340196 108876
rect 340892 90982 340920 362918
rect 340984 163538 341012 382910
rect 341536 238610 341564 396714
rect 342996 378820 343048 378826
rect 342996 378762 343048 378768
rect 342260 361684 342312 361690
rect 342260 361626 342312 361632
rect 341524 238604 341576 238610
rect 341524 238546 341576 238552
rect 341524 225616 341576 225622
rect 341524 225558 341576 225564
rect 341064 184272 341116 184278
rect 341064 184214 341116 184220
rect 340972 163532 341024 163538
rect 340972 163474 341024 163480
rect 341076 151774 341104 184214
rect 341064 151768 341116 151774
rect 341064 151710 341116 151716
rect 340972 144220 341024 144226
rect 340972 144162 341024 144168
rect 340880 90976 340932 90982
rect 340880 90918 340932 90924
rect 340892 90370 340920 90918
rect 340880 90364 340932 90370
rect 340880 90306 340932 90312
rect 340142 28928 340198 28937
rect 340142 28863 340198 28872
rect 340156 28257 340184 28863
rect 340142 28248 340198 28257
rect 340142 28183 340198 28192
rect 336752 16546 337056 16574
rect 338224 16546 338712 16574
rect 336004 3596 336056 3602
rect 336004 3538 336056 3544
rect 335924 3454 336320 3482
rect 336292 480 336320 3454
rect 335054 354 335166 480
rect 334728 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 340156 6914 340184 28183
rect 339880 6886 340184 6914
rect 339880 480 339908 6886
rect 340984 3670 341012 144162
rect 341536 58002 341564 225558
rect 341524 57996 341576 58002
rect 341524 57938 341576 57944
rect 340972 3664 341024 3670
rect 340972 3606 341024 3612
rect 341536 3534 341564 57938
rect 342272 41410 342300 361626
rect 342904 287088 342956 287094
rect 342904 287030 342956 287036
rect 342442 187096 342498 187105
rect 342442 187031 342498 187040
rect 342352 177336 342404 177342
rect 342352 177278 342404 177284
rect 342364 115938 342392 177278
rect 342456 136542 342484 187031
rect 342444 136536 342496 136542
rect 342444 136478 342496 136484
rect 342352 115932 342404 115938
rect 342352 115874 342404 115880
rect 342916 95266 342944 287030
rect 343008 224806 343036 378762
rect 342996 224800 343048 224806
rect 342996 224742 343048 224748
rect 343008 224505 343036 224742
rect 342994 224496 343050 224505
rect 342994 224431 343050 224440
rect 343652 126954 343680 396743
rect 343744 389842 343772 399758
rect 343824 392760 343876 392766
rect 343824 392702 343876 392708
rect 343732 389836 343784 389842
rect 343732 389778 343784 389784
rect 343836 296714 343864 392702
rect 345754 382936 345810 382945
rect 345754 382871 345810 382880
rect 345664 352504 345716 352510
rect 345664 352446 345716 352452
rect 344284 340196 344336 340202
rect 344284 340138 344336 340144
rect 343744 296686 343864 296714
rect 343744 291174 343772 296686
rect 343732 291168 343784 291174
rect 343732 291110 343784 291116
rect 343744 290494 343772 291110
rect 343732 290488 343784 290494
rect 343732 290430 343784 290436
rect 343824 188624 343876 188630
rect 343824 188566 343876 188572
rect 343730 178664 343786 178673
rect 343730 178599 343786 178608
rect 343744 129742 343772 178599
rect 343836 151774 343864 188566
rect 344296 176798 344324 340138
rect 345572 227044 345624 227050
rect 345572 226986 345624 226992
rect 345584 226234 345612 226986
rect 345572 226228 345624 226234
rect 345572 226170 345624 226176
rect 345020 210452 345072 210458
rect 345020 210394 345072 210400
rect 344284 176792 344336 176798
rect 344284 176734 344336 176740
rect 343824 151768 343876 151774
rect 343824 151710 343876 151716
rect 343836 151065 343864 151710
rect 343822 151056 343878 151065
rect 343822 150991 343878 151000
rect 343824 140820 343876 140826
rect 343824 140762 343876 140768
rect 343836 136610 343864 140762
rect 343824 136604 343876 136610
rect 343824 136546 343876 136552
rect 343732 129736 343784 129742
rect 343732 129678 343784 129684
rect 342996 126948 343048 126954
rect 342996 126890 343048 126896
rect 343640 126948 343692 126954
rect 343640 126890 343692 126896
rect 342904 95260 342956 95266
rect 342904 95202 342956 95208
rect 343008 50454 343036 126890
rect 344296 94518 344324 176734
rect 345032 122806 345060 210394
rect 345112 182980 345164 182986
rect 345112 182922 345164 182928
rect 345124 147558 345152 182922
rect 345112 147552 345164 147558
rect 345112 147494 345164 147500
rect 345020 122800 345072 122806
rect 345020 122742 345072 122748
rect 345676 111110 345704 352446
rect 345768 263566 345796 382871
rect 346308 353320 346360 353326
rect 346308 353262 346360 353268
rect 346320 352578 346348 353262
rect 346308 352572 346360 352578
rect 346308 352514 346360 352520
rect 345848 316872 345900 316878
rect 345848 316814 345900 316820
rect 345756 263560 345808 263566
rect 345756 263502 345808 263508
rect 345756 226228 345808 226234
rect 345756 226170 345808 226176
rect 345664 111104 345716 111110
rect 345664 111046 345716 111052
rect 345768 100706 345796 226170
rect 345860 223378 345888 316814
rect 345848 223372 345900 223378
rect 345848 223314 345900 223320
rect 346412 140826 346440 399758
rect 347780 396908 347832 396914
rect 347780 396850 347832 396856
rect 346492 392828 346544 392834
rect 346492 392770 346544 392776
rect 346504 206922 346532 392770
rect 347044 363792 347096 363798
rect 347044 363734 347096 363740
rect 347056 235754 347084 363734
rect 347044 235748 347096 235754
rect 347044 235690 347096 235696
rect 347792 227118 347820 396850
rect 347884 386238 347912 399774
rect 350644 399758 351638 399786
rect 354140 399894 354214 399922
rect 350540 392012 350592 392018
rect 350540 391954 350592 391960
rect 347872 386232 347924 386238
rect 347872 386174 347924 386180
rect 349436 360392 349488 360398
rect 349436 360334 349488 360340
rect 348424 326460 348476 326466
rect 348424 326402 348476 326408
rect 347780 227112 347832 227118
rect 347780 227054 347832 227060
rect 346584 211812 346636 211818
rect 346584 211754 346636 211760
rect 346492 206916 346544 206922
rect 346492 206858 346544 206864
rect 346492 186992 346544 186998
rect 346492 186934 346544 186940
rect 346400 140820 346452 140826
rect 346400 140762 346452 140768
rect 346504 120086 346532 186934
rect 346596 121378 346624 211754
rect 347688 206916 347740 206922
rect 347688 206858 347740 206864
rect 347700 206310 347728 206858
rect 347688 206304 347740 206310
rect 347688 206246 347740 206252
rect 347778 196616 347834 196625
rect 347778 196551 347834 196560
rect 346676 180396 346728 180402
rect 346676 180338 346728 180344
rect 346688 146266 346716 180338
rect 346676 146260 346728 146266
rect 346676 146202 346728 146208
rect 346584 121372 346636 121378
rect 346584 121314 346636 121320
rect 346492 120080 346544 120086
rect 346492 120022 346544 120028
rect 347226 117328 347282 117337
rect 347226 117263 347228 117272
rect 347280 117263 347282 117272
rect 347228 117234 347280 117240
rect 347240 116618 347268 117234
rect 347228 116612 347280 116618
rect 347228 116554 347280 116560
rect 347792 110430 347820 196551
rect 347870 180024 347926 180033
rect 347870 179959 347926 179968
rect 347884 125594 347912 179959
rect 348436 178702 348464 326402
rect 349250 202192 349306 202201
rect 349250 202127 349306 202136
rect 349264 201521 349292 202127
rect 349250 201512 349306 201521
rect 349250 201447 349306 201456
rect 348424 178696 348476 178702
rect 348424 178638 348476 178644
rect 347964 175976 348016 175982
rect 347964 175918 348016 175924
rect 347976 137970 348004 175918
rect 347964 137964 348016 137970
rect 347964 137906 348016 137912
rect 347872 125588 347924 125594
rect 347872 125530 347924 125536
rect 347780 110424 347832 110430
rect 347780 110366 347832 110372
rect 345756 100700 345808 100706
rect 345756 100642 345808 100648
rect 344284 94512 344336 94518
rect 344284 94454 344336 94460
rect 347044 73976 347096 73982
rect 347044 73918 347096 73924
rect 346400 73840 346452 73846
rect 346400 73782 346452 73788
rect 345020 61396 345072 61402
rect 345020 61338 345072 61344
rect 345032 58002 345060 61338
rect 345020 57996 345072 58002
rect 345020 57938 345072 57944
rect 342996 50448 343048 50454
rect 342996 50390 343048 50396
rect 342352 50380 342404 50386
rect 342352 50322 342404 50328
rect 342260 41404 342312 41410
rect 342260 41346 342312 41352
rect 342272 40798 342300 41346
rect 342260 40792 342312 40798
rect 342260 40734 342312 40740
rect 342364 16574 342392 50322
rect 342904 49020 342956 49026
rect 342904 48962 342956 48968
rect 342916 28937 342944 48962
rect 345756 35284 345808 35290
rect 345756 35226 345808 35232
rect 342902 28928 342958 28937
rect 342902 28863 342958 28872
rect 342364 16546 342944 16574
rect 342168 3664 342220 3670
rect 342168 3606 342220 3612
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 341524 3528 341576 3534
rect 341524 3470 341576 3476
rect 340984 480 341012 3470
rect 342180 480 342208 3606
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 345768 10946 345796 35226
rect 346412 16574 346440 73782
rect 346412 16546 346992 16574
rect 345296 10940 345348 10946
rect 345296 10882 345348 10888
rect 345756 10940 345808 10946
rect 345756 10882 345808 10888
rect 344560 3596 344612 3602
rect 344560 3538 344612 3544
rect 344572 480 344600 3538
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 10882
rect 346964 480 346992 16546
rect 347056 6798 347084 73918
rect 348424 13116 348476 13122
rect 348424 13058 348476 13064
rect 348436 6798 348464 13058
rect 349160 11008 349212 11014
rect 349160 10950 349212 10956
rect 347044 6792 347096 6798
rect 347044 6734 347096 6740
rect 348424 6792 348476 6798
rect 348424 6734 348476 6740
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 354 348138 480
rect 348436 354 348464 6734
rect 349172 3346 349200 10950
rect 349264 3534 349292 201447
rect 349344 180192 349396 180198
rect 349344 180134 349396 180140
rect 349356 128314 349384 180134
rect 349344 128308 349396 128314
rect 349344 128250 349396 128256
rect 349448 8294 349476 360334
rect 349804 358964 349856 358970
rect 349804 358906 349856 358912
rect 349816 233918 349844 358906
rect 349896 281580 349948 281586
rect 349896 281522 349948 281528
rect 349908 242185 349936 281522
rect 349894 242176 349950 242185
rect 349894 242111 349950 242120
rect 349896 234660 349948 234666
rect 349896 234602 349948 234608
rect 349804 233912 349856 233918
rect 349804 233854 349856 233860
rect 349908 171086 349936 234602
rect 349896 171080 349948 171086
rect 349896 171022 349948 171028
rect 350552 59362 350580 391954
rect 350644 192506 350672 399758
rect 354140 398478 354168 399894
rect 356762 399786 356790 400044
rect 358694 399838 358722 400044
rect 356716 399758 356790 399786
rect 357440 399832 357492 399838
rect 357440 399774 357492 399780
rect 358682 399832 358734 399838
rect 361270 399786 361298 400044
rect 363846 399786 363874 400044
rect 365778 399786 365806 400044
rect 368354 399838 368382 400044
rect 358682 399774 358734 399780
rect 353392 398472 353444 398478
rect 353392 398414 353444 398420
rect 354128 398472 354180 398478
rect 354128 398414 354180 398420
rect 351920 392692 351972 392698
rect 351920 392634 351972 392640
rect 351184 356312 351236 356318
rect 351184 356254 351236 356260
rect 351196 240825 351224 356254
rect 351276 279472 351328 279478
rect 351276 279414 351328 279420
rect 351182 240816 351238 240825
rect 351182 240751 351238 240760
rect 351184 228540 351236 228546
rect 351184 228482 351236 228488
rect 350632 192500 350684 192506
rect 350632 192442 350684 192448
rect 350540 59356 350592 59362
rect 350540 59298 350592 59304
rect 350552 58818 350580 59298
rect 350540 58812 350592 58818
rect 350540 58754 350592 58760
rect 349804 33788 349856 33794
rect 349804 33730 349856 33736
rect 349816 11014 349844 33730
rect 349804 11008 349856 11014
rect 349804 10950 349856 10956
rect 349436 8288 349488 8294
rect 349436 8230 349488 8236
rect 349712 8288 349764 8294
rect 349712 8230 349764 8236
rect 349724 7614 349752 8230
rect 349712 7608 349764 7614
rect 349712 7550 349764 7556
rect 351196 4146 351224 228482
rect 351288 155242 351316 279414
rect 351932 210458 351960 392634
rect 352564 370524 352616 370530
rect 352564 370466 352616 370472
rect 352576 235686 352604 370466
rect 353298 357504 353354 357513
rect 353298 357439 353354 357448
rect 352564 235680 352616 235686
rect 352564 235622 352616 235628
rect 351920 210452 351972 210458
rect 351920 210394 351972 210400
rect 351920 203856 351972 203862
rect 351920 203798 351972 203804
rect 351368 180260 351420 180266
rect 351368 180202 351420 180208
rect 351380 171086 351408 180202
rect 351368 171080 351420 171086
rect 351368 171022 351420 171028
rect 351276 155236 351328 155242
rect 351276 155178 351328 155184
rect 351380 102134 351408 171022
rect 351932 114442 351960 203798
rect 352012 203584 352064 203590
rect 352012 203526 352064 203532
rect 352024 149054 352052 203526
rect 352012 149048 352064 149054
rect 352012 148990 352064 148996
rect 351920 114436 351972 114442
rect 351920 114378 351972 114384
rect 351368 102128 351420 102134
rect 351368 102070 351420 102076
rect 353312 93838 353340 357439
rect 353404 234666 353432 398414
rect 356716 397526 356744 399758
rect 356796 398132 356848 398138
rect 356796 398074 356848 398080
rect 355232 397520 355284 397526
rect 355232 397462 355284 397468
rect 356704 397520 356756 397526
rect 356704 397462 356756 397468
rect 355244 396778 355272 397462
rect 355232 396772 355284 396778
rect 355232 396714 355284 396720
rect 354678 396672 354734 396681
rect 354678 396607 354734 396616
rect 353944 333328 353996 333334
rect 353944 333270 353996 333276
rect 353956 263566 353984 333270
rect 354588 281648 354640 281654
rect 354588 281590 354640 281596
rect 353944 263560 353996 263566
rect 353944 263502 353996 263508
rect 353392 234660 353444 234666
rect 353392 234602 353444 234608
rect 353944 233980 353996 233986
rect 353944 233922 353996 233928
rect 353956 125594 353984 233922
rect 354036 139392 354088 139398
rect 354036 139334 354088 139340
rect 353944 125588 353996 125594
rect 353944 125530 353996 125536
rect 353300 93832 353352 93838
rect 353300 93774 353352 93780
rect 353312 93158 353340 93774
rect 353300 93152 353352 93158
rect 353300 93094 353352 93100
rect 354048 61538 354076 139334
rect 354600 115938 354628 281590
rect 354692 139398 354720 396607
rect 355508 393984 355560 393990
rect 355508 393926 355560 393932
rect 355324 347064 355376 347070
rect 355324 347006 355376 347012
rect 355336 197334 355364 347006
rect 355416 331900 355468 331906
rect 355416 331842 355468 331848
rect 354772 197328 354824 197334
rect 354772 197270 354824 197276
rect 355324 197328 355376 197334
rect 355324 197270 355376 197276
rect 354680 139392 354732 139398
rect 354680 139334 354732 139340
rect 354784 118658 354812 197270
rect 355428 195974 355456 331842
rect 355520 276690 355548 393926
rect 356808 393314 356836 398074
rect 357348 395480 357400 395486
rect 357348 395422 357400 395428
rect 357360 395350 357388 395422
rect 357348 395344 357400 395350
rect 357348 395286 357400 395292
rect 356716 393286 356836 393314
rect 356716 376106 356744 393286
rect 356060 376100 356112 376106
rect 356060 376042 356112 376048
rect 356704 376100 356756 376106
rect 356704 376042 356756 376048
rect 355508 276684 355560 276690
rect 355508 276626 355560 276632
rect 354864 195968 354916 195974
rect 354864 195910 354916 195916
rect 355416 195968 355468 195974
rect 355416 195910 355468 195916
rect 354876 139330 354904 195910
rect 356072 155922 356100 376042
rect 356796 303000 356848 303006
rect 356796 302942 356848 302948
rect 356704 268388 356756 268394
rect 356704 268330 356756 268336
rect 356244 198008 356296 198014
rect 356244 197950 356296 197956
rect 356152 195288 356204 195294
rect 356152 195230 356204 195236
rect 356060 155916 356112 155922
rect 356060 155858 356112 155864
rect 355324 149116 355376 149122
rect 355324 149058 355376 149064
rect 354864 139324 354916 139330
rect 354864 139266 354916 139272
rect 354772 118652 354824 118658
rect 354772 118594 354824 118600
rect 354588 115932 354640 115938
rect 354588 115874 354640 115880
rect 355336 87650 355364 149058
rect 356164 106282 356192 195230
rect 356256 131102 356284 197950
rect 356244 131096 356296 131102
rect 356244 131038 356296 131044
rect 356152 106276 356204 106282
rect 356152 106218 356204 106224
rect 356716 95198 356744 268330
rect 356808 233034 356836 302942
rect 357360 237318 357388 395286
rect 357348 237312 357400 237318
rect 357348 237254 357400 237260
rect 356796 233028 356848 233034
rect 356796 232970 356848 232976
rect 357452 133210 357480 399774
rect 360212 399758 361298 399786
rect 363616 399758 363874 399786
rect 365732 399758 365806 399786
rect 367100 399832 367152 399838
rect 367100 399774 367152 399780
rect 368342 399832 368394 399838
rect 370930 399786 370958 400044
rect 373506 399786 373534 400044
rect 375438 399786 375466 400044
rect 378014 399786 378042 400044
rect 380590 399786 380618 400044
rect 382522 399786 382550 400044
rect 385098 399922 385126 400044
rect 385098 399894 385172 399922
rect 368342 399774 368394 399780
rect 359280 399628 359332 399634
rect 359280 399570 359332 399576
rect 359292 398886 359320 399570
rect 358820 398880 358872 398886
rect 358820 398822 358872 398828
rect 359280 398880 359332 398886
rect 359280 398822 359332 398828
rect 358084 299600 358136 299606
rect 358084 299542 358136 299548
rect 357532 242956 357584 242962
rect 357532 242898 357584 242904
rect 357544 133890 357572 242898
rect 358096 235890 358124 299542
rect 358832 242962 358860 398822
rect 359464 361616 359516 361622
rect 359464 361558 359516 361564
rect 359476 342242 359504 361558
rect 359464 342236 359516 342242
rect 359464 342178 359516 342184
rect 359476 341630 359504 342178
rect 359464 341624 359516 341630
rect 359464 341566 359516 341572
rect 360016 341624 360068 341630
rect 360016 341566 360068 341572
rect 359464 320884 359516 320890
rect 359464 320826 359516 320832
rect 358820 242956 358872 242962
rect 358820 242898 358872 242904
rect 358084 235884 358136 235890
rect 358084 235826 358136 235832
rect 359476 215286 359504 320826
rect 360028 280906 360056 341566
rect 360108 302388 360160 302394
rect 360108 302330 360160 302336
rect 360016 280900 360068 280906
rect 360016 280842 360068 280848
rect 359648 273964 359700 273970
rect 359648 273906 359700 273912
rect 359660 273290 359688 273906
rect 359648 273284 359700 273290
rect 359648 273226 359700 273232
rect 360016 273284 360068 273290
rect 360016 273226 360068 273232
rect 358820 215280 358872 215286
rect 358820 215222 358872 215228
rect 359464 215280 359516 215286
rect 359464 215222 359516 215228
rect 357532 133884 357584 133890
rect 357532 133826 357584 133832
rect 357440 133204 357492 133210
rect 357440 133146 357492 133152
rect 358832 114510 358860 215222
rect 360028 148374 360056 273226
rect 360016 148368 360068 148374
rect 360016 148310 360068 148316
rect 359464 145104 359516 145110
rect 359464 145046 359516 145052
rect 358820 114504 358872 114510
rect 358820 114446 358872 114452
rect 356796 96688 356848 96694
rect 356796 96630 356848 96636
rect 356704 95192 356756 95198
rect 356704 95134 356756 95140
rect 355324 87644 355376 87650
rect 355324 87586 355376 87592
rect 354036 61532 354088 61538
rect 354036 61474 354088 61480
rect 355324 60036 355376 60042
rect 355324 59978 355376 59984
rect 351184 4140 351236 4146
rect 351184 4082 351236 4088
rect 351644 4140 351696 4146
rect 351644 4082 351696 4088
rect 349252 3528 349304 3534
rect 349252 3470 349304 3476
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 349172 3318 349292 3346
rect 349264 480 349292 3318
rect 350460 480 350488 3470
rect 351656 480 351684 4082
rect 355336 3466 355364 59978
rect 356808 8226 356836 96630
rect 359476 41342 359504 145046
rect 360120 137970 360148 302330
rect 360108 137964 360160 137970
rect 360108 137906 360160 137912
rect 360212 113830 360240 399758
rect 363616 395826 363644 399758
rect 365076 396772 365128 396778
rect 365076 396714 365128 396720
rect 363604 395820 363656 395826
rect 363604 395762 363656 395768
rect 363616 365090 363644 395762
rect 364984 374672 365036 374678
rect 364984 374614 365036 374620
rect 364996 374134 365024 374614
rect 364984 374128 365036 374134
rect 364984 374070 365036 374076
rect 363604 365084 363656 365090
rect 363604 365026 363656 365032
rect 362224 340196 362276 340202
rect 362224 340138 362276 340144
rect 360844 312588 360896 312594
rect 360844 312530 360896 312536
rect 360292 309868 360344 309874
rect 360292 309810 360344 309816
rect 360304 309194 360332 309810
rect 360292 309188 360344 309194
rect 360292 309130 360344 309136
rect 360856 131102 360884 312530
rect 361488 309188 361540 309194
rect 361488 309130 361540 309136
rect 361500 218822 361528 309130
rect 361488 218816 361540 218822
rect 361488 218758 361540 218764
rect 360844 131096 360896 131102
rect 360844 131038 360896 131044
rect 360936 129804 360988 129810
rect 360936 129746 360988 129752
rect 360200 113824 360252 113830
rect 360200 113766 360252 113772
rect 359464 41336 359516 41342
rect 359464 41278 359516 41284
rect 360948 13802 360976 129746
rect 362236 129742 362264 340138
rect 363602 336016 363658 336025
rect 363602 335951 363658 335960
rect 362960 316804 363012 316810
rect 362960 316746 363012 316752
rect 362972 316062 363000 316746
rect 362960 316056 363012 316062
rect 362960 315998 363012 316004
rect 362868 303680 362920 303686
rect 362868 303622 362920 303628
rect 362224 129736 362276 129742
rect 362224 129678 362276 129684
rect 362880 114510 362908 303622
rect 362960 247104 363012 247110
rect 362960 247046 363012 247052
rect 362972 246362 363000 247046
rect 362960 246356 363012 246362
rect 362960 246298 363012 246304
rect 362958 231840 363014 231849
rect 362958 231775 363014 231784
rect 362972 231742 363000 231775
rect 362960 231736 363012 231742
rect 362960 231678 363012 231684
rect 362868 114504 362920 114510
rect 362868 114446 362920 114452
rect 363616 114442 363644 335951
rect 364248 316056 364300 316062
rect 364248 315998 364300 316004
rect 364156 264988 364208 264994
rect 364156 264930 364208 264936
rect 363696 246356 363748 246362
rect 363696 246298 363748 246304
rect 363708 151094 363736 246298
rect 364168 231849 364196 264930
rect 364154 231840 364210 231849
rect 364154 231775 364210 231784
rect 364260 218754 364288 315998
rect 364706 246256 364762 246265
rect 364706 246191 364762 246200
rect 364720 245682 364748 246191
rect 364708 245676 364760 245682
rect 364708 245618 364760 245624
rect 364248 218748 364300 218754
rect 364248 218690 364300 218696
rect 363788 188352 363840 188358
rect 363788 188294 363840 188300
rect 363696 151088 363748 151094
rect 363696 151030 363748 151036
rect 363604 114436 363656 114442
rect 363604 114378 363656 114384
rect 363604 107704 363656 107710
rect 363604 107646 363656 107652
rect 363616 60110 363644 107646
rect 363800 106282 363828 188294
rect 363788 106276 363840 106282
rect 363788 106218 363840 106224
rect 363604 60104 363656 60110
rect 363604 60046 363656 60052
rect 364996 38622 365024 374070
rect 365088 230450 365116 396714
rect 365732 387190 365760 399758
rect 367008 387864 367060 387870
rect 367008 387806 367060 387812
rect 367020 387190 367048 387806
rect 365720 387184 365772 387190
rect 365720 387126 365772 387132
rect 367008 387184 367060 387190
rect 367008 387126 367060 387132
rect 366364 367804 366416 367810
rect 366364 367746 366416 367752
rect 365260 334620 365312 334626
rect 365260 334562 365312 334568
rect 365168 290488 365220 290494
rect 365168 290430 365220 290436
rect 365076 230444 365128 230450
rect 365076 230386 365128 230392
rect 365076 185632 365128 185638
rect 365076 185574 365128 185580
rect 365088 117298 365116 185574
rect 365180 142118 365208 290430
rect 365272 259418 365300 334562
rect 365260 259412 365312 259418
rect 365260 259354 365312 259360
rect 365628 245676 365680 245682
rect 365628 245618 365680 245624
rect 365640 151162 365668 245618
rect 365628 151156 365680 151162
rect 365628 151098 365680 151104
rect 365168 142112 365220 142118
rect 365168 142054 365220 142060
rect 365076 117292 365128 117298
rect 365076 117234 365128 117240
rect 366376 109002 366404 367746
rect 367008 289128 367060 289134
rect 367008 289070 367060 289076
rect 367020 288454 367048 289070
rect 367008 288448 367060 288454
rect 367008 288390 367060 288396
rect 367020 121446 367048 288390
rect 367112 212498 367140 399774
rect 369872 399758 370958 399786
rect 372632 399758 373534 399786
rect 375392 399758 375466 399786
rect 377968 399758 378042 399786
rect 380544 399758 380618 399786
rect 382476 399758 382550 399786
rect 368388 399560 368440 399566
rect 368388 399502 368440 399508
rect 368400 399022 368428 399502
rect 368388 399016 368440 399022
rect 368388 398958 368440 398964
rect 367744 319524 367796 319530
rect 367744 319466 367796 319472
rect 367100 212492 367152 212498
rect 367100 212434 367152 212440
rect 367112 134570 367140 212434
rect 367100 134564 367152 134570
rect 367100 134506 367152 134512
rect 367008 121440 367060 121446
rect 367008 121382 367060 121388
rect 366364 108996 366416 109002
rect 366364 108938 366416 108944
rect 367756 107642 367784 319466
rect 368296 251864 368348 251870
rect 368296 251806 368348 251812
rect 368308 251258 368336 251806
rect 368296 251252 368348 251258
rect 368296 251194 368348 251200
rect 367744 107636 367796 107642
rect 367744 107578 367796 107584
rect 365076 105596 365128 105602
rect 365076 105538 365128 105544
rect 364984 38616 365036 38622
rect 364984 38558 365036 38564
rect 365088 38010 365116 105538
rect 368308 95130 368336 251194
rect 368400 235890 368428 398958
rect 369676 395344 369728 395350
rect 369676 395286 369728 395292
rect 368480 392624 368532 392630
rect 368480 392566 368532 392572
rect 368388 235884 368440 235890
rect 368388 235826 368440 235832
rect 368492 191826 368520 392566
rect 369124 369164 369176 369170
rect 369124 369106 369176 369112
rect 368480 191820 368532 191826
rect 368480 191762 368532 191768
rect 368940 191820 368992 191826
rect 368940 191762 368992 191768
rect 368952 191146 368980 191762
rect 368940 191140 368992 191146
rect 368940 191082 368992 191088
rect 369136 169726 369164 369106
rect 369688 232558 369716 395286
rect 369872 322250 369900 399758
rect 371976 395412 372028 395418
rect 371976 395354 372028 395360
rect 371884 334688 371936 334694
rect 371884 334630 371936 334636
rect 369860 322244 369912 322250
rect 369860 322186 369912 322192
rect 370504 322244 370556 322250
rect 370504 322186 370556 322192
rect 369768 297424 369820 297430
rect 369768 297366 369820 297372
rect 369780 296750 369808 297366
rect 369768 296744 369820 296750
rect 369768 296686 369820 296692
rect 369676 232552 369728 232558
rect 369676 232494 369728 232500
rect 369124 169720 369176 169726
rect 369124 169662 369176 169668
rect 369124 145580 369176 145586
rect 369124 145522 369176 145528
rect 368296 95124 368348 95130
rect 368296 95066 368348 95072
rect 365628 38616 365680 38622
rect 365628 38558 365680 38564
rect 365076 38004 365128 38010
rect 365076 37946 365128 37952
rect 365640 37942 365668 38558
rect 365628 37936 365680 37942
rect 365628 37878 365680 37884
rect 369136 24818 369164 145522
rect 369780 91050 369808 296686
rect 369860 286340 369912 286346
rect 369860 286282 369912 286288
rect 369872 285734 369900 286282
rect 369860 285728 369912 285734
rect 369860 285670 369912 285676
rect 370516 121378 370544 322186
rect 371148 285728 371200 285734
rect 371148 285670 371200 285676
rect 371056 259412 371108 259418
rect 371056 259354 371108 259360
rect 371068 258126 371096 259354
rect 371056 258120 371108 258126
rect 371056 258062 371108 258068
rect 371068 209098 371096 258062
rect 371160 229906 371188 285670
rect 371240 280900 371292 280906
rect 371240 280842 371292 280848
rect 371252 280226 371280 280842
rect 371240 280220 371292 280226
rect 371240 280162 371292 280168
rect 371148 229900 371200 229906
rect 371148 229842 371200 229848
rect 371056 209092 371108 209098
rect 371056 209034 371108 209040
rect 371896 149054 371924 334630
rect 371988 278050 372016 395354
rect 372632 365158 372660 399758
rect 375392 395486 375420 399758
rect 377968 398449 377996 399758
rect 380544 398682 380572 399758
rect 380624 399492 380676 399498
rect 380624 399434 380676 399440
rect 380636 398682 380664 399434
rect 380532 398676 380584 398682
rect 380532 398618 380584 398624
rect 380624 398676 380676 398682
rect 380624 398618 380676 398624
rect 376758 398440 376814 398449
rect 376758 398375 376814 398384
rect 377954 398440 378010 398449
rect 377954 398375 378010 398384
rect 375380 395480 375432 395486
rect 375380 395422 375432 395428
rect 373908 393304 373960 393310
rect 373908 393246 373960 393252
rect 372620 365152 372672 365158
rect 372620 365094 372672 365100
rect 373264 315308 373316 315314
rect 373264 315250 373316 315256
rect 372620 311908 372672 311914
rect 372620 311850 372672 311856
rect 372632 309874 372660 311850
rect 372620 309868 372672 309874
rect 372620 309810 372672 309816
rect 373276 290494 373304 315250
rect 373724 303748 373776 303754
rect 373724 303690 373776 303696
rect 373264 290488 373316 290494
rect 373264 290430 373316 290436
rect 372528 280220 372580 280226
rect 372528 280162 372580 280168
rect 371976 278044 372028 278050
rect 371976 277986 372028 277992
rect 371976 276072 372028 276078
rect 371976 276014 372028 276020
rect 371988 223514 372016 276014
rect 372540 240854 372568 280162
rect 373264 253224 373316 253230
rect 373264 253166 373316 253172
rect 372528 240848 372580 240854
rect 372528 240790 372580 240796
rect 371976 223508 372028 223514
rect 371976 223450 372028 223456
rect 371884 149048 371936 149054
rect 371884 148990 371936 148996
rect 370504 121372 370556 121378
rect 370504 121314 370556 121320
rect 371988 95062 372016 223450
rect 373276 144294 373304 253166
rect 373356 247716 373408 247722
rect 373356 247658 373408 247664
rect 373368 235958 373396 247658
rect 373736 241913 373764 303690
rect 373816 290488 373868 290494
rect 373816 290430 373868 290436
rect 373722 241904 373778 241913
rect 373722 241839 373778 241848
rect 373356 235952 373408 235958
rect 373356 235894 373408 235900
rect 373828 205018 373856 290430
rect 373920 277438 373948 393246
rect 374644 392760 374696 392766
rect 374644 392702 374696 392708
rect 373908 277432 373960 277438
rect 373908 277374 373960 277380
rect 373816 205012 373868 205018
rect 373816 204954 373868 204960
rect 373356 147688 373408 147694
rect 373356 147630 373408 147636
rect 373264 144288 373316 144294
rect 373264 144230 373316 144236
rect 371976 95056 372028 95062
rect 371976 94998 372028 95004
rect 369768 91044 369820 91050
rect 369768 90986 369820 90992
rect 373368 47734 373396 147630
rect 374656 103494 374684 392702
rect 376772 369170 376800 398375
rect 382476 395418 382504 399758
rect 385144 398546 385172 399894
rect 387674 399838 387702 400044
rect 386420 399832 386472 399838
rect 386420 399774 386472 399780
rect 387662 399832 387714 399838
rect 390250 399786 390278 400044
rect 392182 399786 392210 400044
rect 394758 399786 394786 400044
rect 397334 399838 397362 400044
rect 387662 399774 387714 399780
rect 385132 398540 385184 398546
rect 385132 398482 385184 398488
rect 385144 397526 385172 398482
rect 385132 397520 385184 397526
rect 385132 397462 385184 397468
rect 385684 397520 385736 397526
rect 385684 397462 385736 397468
rect 382464 395412 382516 395418
rect 382464 395354 382516 395360
rect 377404 392692 377456 392698
rect 377404 392634 377456 392640
rect 376760 369164 376812 369170
rect 376760 369106 376812 369112
rect 375104 359508 375156 359514
rect 375104 359450 375156 359456
rect 374736 302932 374788 302938
rect 374736 302874 374788 302880
rect 374748 302258 374776 302874
rect 374736 302252 374788 302258
rect 374736 302194 374788 302200
rect 375116 237182 375144 359450
rect 377416 316878 377444 392634
rect 379428 392624 379480 392630
rect 379428 392566 379480 392572
rect 379336 369164 379388 369170
rect 379336 369106 379388 369112
rect 379244 334620 379296 334626
rect 379244 334562 379296 334568
rect 379152 318096 379204 318102
rect 379152 318038 379204 318044
rect 377404 316872 377456 316878
rect 377404 316814 377456 316820
rect 377496 307148 377548 307154
rect 377496 307090 377548 307096
rect 376208 302320 376260 302326
rect 376208 302262 376260 302268
rect 375288 302252 375340 302258
rect 375288 302194 375340 302200
rect 375196 277636 375248 277642
rect 375196 277578 375248 277584
rect 375208 277438 375236 277578
rect 375196 277432 375248 277438
rect 375196 277374 375248 277380
rect 375104 237176 375156 237182
rect 375104 237118 375156 237124
rect 375208 152590 375236 277374
rect 375196 152584 375248 152590
rect 375196 152526 375248 152532
rect 374644 103488 374696 103494
rect 374644 103430 374696 103436
rect 374642 102776 374698 102785
rect 374642 102711 374698 102720
rect 374656 100026 374684 102711
rect 374644 100020 374696 100026
rect 374644 99962 374696 99968
rect 374656 86358 374684 99962
rect 375300 92342 375328 302194
rect 376116 300960 376168 300966
rect 376116 300902 376168 300908
rect 376024 282940 376076 282946
rect 376024 282882 376076 282888
rect 376036 239018 376064 282882
rect 376128 275330 376156 300902
rect 376220 280838 376248 302262
rect 376942 297120 376998 297129
rect 376942 297055 376998 297064
rect 376956 296750 376984 297055
rect 376944 296744 376996 296750
rect 376944 296686 376996 296692
rect 377402 293040 377458 293049
rect 377402 292975 377458 292984
rect 376942 291000 376998 291009
rect 376942 290935 376998 290944
rect 376956 290494 376984 290935
rect 376944 290488 376996 290494
rect 376944 290430 376996 290436
rect 376942 288960 376998 288969
rect 376942 288895 376998 288904
rect 376956 288454 376984 288895
rect 376944 288448 376996 288454
rect 376944 288390 376996 288396
rect 376942 286920 376998 286929
rect 376942 286855 376998 286864
rect 376956 285734 376984 286855
rect 376944 285728 376996 285734
rect 376944 285670 376996 285676
rect 377310 284200 377366 284209
rect 377310 284135 377366 284144
rect 377324 283626 377352 284135
rect 377312 283620 377364 283626
rect 377312 283562 377364 283568
rect 376942 282160 376998 282169
rect 376942 282095 376998 282104
rect 376956 281586 376984 282095
rect 376944 281580 376996 281586
rect 376944 281522 376996 281528
rect 376208 280832 376260 280838
rect 376208 280774 376260 280780
rect 376942 280256 376998 280265
rect 376942 280191 376944 280200
rect 376996 280191 376998 280200
rect 376944 280162 376996 280168
rect 376758 278080 376814 278089
rect 376758 278015 376814 278024
rect 376772 277642 376800 278015
rect 376760 277636 376812 277642
rect 376760 277578 376812 277584
rect 376116 275324 376168 275330
rect 376116 275266 376168 275272
rect 376942 265160 376998 265169
rect 376942 265095 376998 265104
rect 376956 264994 376984 265095
rect 376944 264988 376996 264994
rect 376944 264930 376996 264936
rect 376576 263628 376628 263634
rect 376576 263570 376628 263576
rect 376114 250200 376170 250209
rect 376114 250135 376170 250144
rect 376024 239012 376076 239018
rect 376024 238954 376076 238960
rect 376128 234598 376156 250135
rect 376588 238746 376616 263570
rect 377312 263560 377364 263566
rect 377312 263502 377364 263508
rect 377324 263265 377352 263502
rect 377310 263256 377366 263265
rect 377310 263191 377366 263200
rect 376942 259040 376998 259049
rect 376942 258975 376998 258984
rect 376956 258126 376984 258975
rect 376944 258120 376996 258126
rect 376944 258062 376996 258068
rect 377312 256012 377364 256018
rect 377312 255954 377364 255960
rect 377324 254425 377352 255954
rect 377310 254416 377366 254425
rect 377310 254351 377366 254360
rect 376942 252240 376998 252249
rect 376942 252175 376998 252184
rect 376956 251258 376984 252175
rect 376944 251252 376996 251258
rect 376944 251194 376996 251200
rect 376942 248160 376998 248169
rect 376942 248095 376998 248104
rect 376956 247110 376984 248095
rect 376944 247104 376996 247110
rect 376944 247046 376996 247052
rect 376942 246120 376998 246129
rect 376942 246055 376998 246064
rect 376956 245682 376984 246055
rect 376944 245676 376996 245682
rect 376944 245618 376996 245624
rect 376666 242040 376722 242049
rect 376666 241975 376722 241984
rect 376576 238740 376628 238746
rect 376576 238682 376628 238688
rect 376116 234592 376168 234598
rect 376116 234534 376168 234540
rect 376024 193928 376076 193934
rect 376024 193870 376076 193876
rect 376036 106962 376064 193870
rect 376128 159390 376156 234534
rect 376680 212430 376708 241975
rect 377416 235822 377444 292975
rect 377508 263634 377536 307090
rect 377954 299296 378010 299305
rect 377954 299231 378010 299240
rect 377968 289814 377996 299231
rect 379164 295322 379192 318038
rect 379152 295316 379204 295322
rect 379152 295258 379204 295264
rect 379164 295225 379192 295258
rect 379150 295216 379206 295225
rect 379150 295151 379206 295160
rect 377956 289808 378008 289814
rect 377956 289750 378008 289756
rect 378784 289808 378836 289814
rect 378784 289750 378836 289756
rect 377864 283620 377916 283626
rect 377864 283562 377916 283568
rect 377772 276072 377824 276078
rect 377770 276040 377772 276049
rect 377824 276040 377826 276049
rect 377770 275975 377826 275984
rect 377770 274000 377826 274009
rect 377770 273935 377826 273944
rect 377784 273290 377812 273935
rect 377772 273284 377824 273290
rect 377772 273226 377824 273232
rect 377496 263628 377548 263634
rect 377496 263570 377548 263576
rect 377404 235816 377456 235822
rect 377404 235758 377456 235764
rect 377416 233986 377444 235758
rect 377404 233980 377456 233986
rect 377404 233922 377456 233928
rect 376668 212424 376720 212430
rect 376668 212366 376720 212372
rect 377876 210458 377904 283562
rect 378046 254416 378102 254425
rect 378046 254351 378102 254360
rect 377954 244080 378010 244089
rect 377954 244015 378010 244024
rect 377968 237153 377996 244015
rect 377954 237144 378010 237153
rect 377954 237079 378010 237088
rect 377968 236201 377996 237079
rect 378060 236706 378088 254351
rect 378048 236700 378100 236706
rect 378048 236642 378100 236648
rect 377954 236192 378010 236201
rect 377954 236127 378010 236136
rect 377956 228404 378008 228410
rect 377956 228346 378008 228352
rect 377864 210452 377916 210458
rect 377864 210394 377916 210400
rect 376116 159384 376168 159390
rect 376116 159326 376168 159332
rect 377404 147756 377456 147762
rect 377404 147698 377456 147704
rect 376668 144288 376720 144294
rect 376668 144230 376720 144236
rect 376680 140078 376708 144230
rect 376668 140072 376720 140078
rect 376668 140014 376720 140020
rect 376024 106956 376076 106962
rect 376024 106898 376076 106904
rect 375288 92336 375340 92342
rect 375288 92278 375340 92284
rect 374644 86352 374696 86358
rect 374644 86294 374696 86300
rect 373356 47728 373408 47734
rect 373356 47670 373408 47676
rect 369124 24812 369176 24818
rect 369124 24754 369176 24760
rect 377416 17338 377444 147698
rect 377968 126886 377996 228346
rect 378046 228304 378102 228313
rect 378046 228239 378102 228248
rect 378060 227769 378088 228239
rect 378046 227760 378102 227769
rect 378046 227695 378102 227704
rect 377956 126880 378008 126886
rect 377956 126822 378008 126828
rect 378060 95334 378088 227695
rect 378796 110430 378824 289750
rect 379256 272105 379284 334562
rect 378874 272096 378930 272105
rect 378874 272031 378930 272040
rect 379242 272096 379298 272105
rect 379242 272031 379298 272040
rect 378888 229094 378916 272031
rect 379244 267708 379296 267714
rect 379244 267650 379296 267656
rect 379256 267209 379284 267650
rect 379242 267200 379298 267209
rect 379242 267135 379298 267144
rect 378888 229066 379008 229094
rect 378980 216646 379008 229066
rect 379256 228478 379284 267135
rect 379348 261225 379376 369106
rect 379440 274009 379468 392566
rect 381544 387116 381596 387122
rect 381544 387058 381596 387064
rect 381556 378894 381584 387058
rect 380900 378888 380952 378894
rect 380900 378830 380952 378836
rect 381544 378888 381596 378894
rect 381544 378830 381596 378836
rect 379520 319456 379572 319462
rect 379520 319398 379572 319404
rect 379532 276049 379560 319398
rect 379612 307216 379664 307222
rect 379612 307158 379664 307164
rect 379624 299305 379652 307158
rect 380912 303754 380940 378830
rect 384304 373312 384356 373318
rect 384304 373254 384356 373260
rect 384316 309194 384344 373254
rect 385040 354748 385092 354754
rect 385040 354690 385092 354696
rect 384304 309188 384356 309194
rect 384304 309130 384356 309136
rect 380900 303748 380952 303754
rect 380900 303690 380952 303696
rect 380912 299962 380940 303690
rect 384316 299962 384344 309130
rect 385052 302394 385080 354690
rect 385696 313478 385724 397462
rect 386432 373998 386460 399774
rect 389192 399758 390278 399786
rect 391952 399758 392210 399786
rect 394712 399758 394786 399786
rect 396080 399832 396132 399838
rect 396080 399774 396132 399780
rect 397322 399832 397374 399838
rect 399266 399786 399294 400044
rect 401842 399786 401870 400044
rect 404418 399786 404446 400044
rect 406994 399838 407022 400044
rect 397322 399774 397374 399780
rect 389192 379642 389220 399758
rect 391204 395412 391256 395418
rect 391204 395354 391256 395360
rect 389180 379636 389232 379642
rect 389180 379578 389232 379584
rect 389824 379636 389876 379642
rect 389824 379578 389876 379584
rect 386420 373992 386472 373998
rect 386420 373934 386472 373940
rect 386328 313948 386380 313954
rect 386328 313890 386380 313896
rect 385684 313472 385736 313478
rect 385684 313414 385736 313420
rect 386340 309942 386368 313890
rect 386328 309936 386380 309942
rect 386328 309878 386380 309884
rect 386432 307222 386460 373934
rect 389836 363662 389864 379578
rect 389824 363656 389876 363662
rect 389824 363598 389876 363604
rect 391216 324970 391244 395354
rect 391952 359514 391980 399758
rect 391940 359508 391992 359514
rect 391940 359450 391992 359456
rect 393964 359508 394016 359514
rect 393964 359450 394016 359456
rect 391204 324964 391256 324970
rect 391204 324906 391256 324912
rect 393976 321570 394004 359450
rect 393964 321564 394016 321570
rect 393964 321506 394016 321512
rect 386512 314628 386564 314634
rect 386512 314570 386564 314576
rect 386420 307216 386472 307222
rect 386420 307158 386472 307164
rect 385040 302388 385092 302394
rect 385040 302330 385092 302336
rect 385776 302388 385828 302394
rect 385776 302330 385828 302336
rect 380912 299934 381294 299962
rect 383962 299934 384344 299962
rect 385788 299948 385816 302330
rect 386524 299962 386552 314570
rect 389180 313472 389232 313478
rect 389180 313414 389232 313420
rect 389192 303686 389220 313414
rect 391204 309868 391256 309874
rect 391204 309810 391256 309816
rect 391216 306406 391244 309810
rect 391204 306400 391256 306406
rect 391204 306342 391256 306348
rect 389180 303680 389232 303686
rect 389180 303622 389232 303628
rect 389192 299962 389220 303622
rect 391216 299962 391244 306342
rect 393976 301034 394004 321506
rect 394712 319530 394740 399758
rect 396092 334694 396120 399774
rect 398852 399758 399294 399786
rect 401796 399758 401870 399786
rect 404372 399758 404446 399786
rect 405740 399832 405792 399838
rect 405740 399774 405792 399780
rect 406982 399832 407034 399838
rect 408926 399786 408954 400044
rect 411502 399786 411530 400044
rect 414078 399786 414106 400044
rect 406982 399774 407034 399780
rect 396080 334688 396132 334694
rect 396080 334630 396132 334636
rect 394700 319524 394752 319530
rect 394700 319466 394752 319472
rect 395344 309936 395396 309942
rect 395344 309878 395396 309884
rect 395356 303686 395384 309878
rect 398852 307154 398880 399758
rect 401796 395350 401824 399758
rect 401784 395344 401836 395350
rect 401784 395286 401836 395292
rect 399484 381540 399536 381546
rect 399484 381482 399536 381488
rect 399496 307834 399524 381482
rect 404372 377534 404400 399758
rect 405752 392766 405780 399774
rect 408880 399758 408954 399786
rect 411456 399758 411530 399786
rect 414032 399758 414106 399786
rect 416010 399786 416038 400044
rect 418586 399786 418614 400044
rect 421162 399786 421190 400044
rect 423738 399786 423766 400044
rect 425670 399786 425698 400044
rect 428246 399786 428274 400044
rect 430822 399786 430850 400044
rect 432754 399786 432782 400044
rect 435330 399786 435358 400044
rect 437906 399786 437934 400044
rect 440482 399786 440510 400044
rect 442414 399786 442442 400044
rect 444990 399786 445018 400044
rect 447566 399786 447594 400044
rect 449498 399786 449526 400044
rect 452074 399786 452102 400044
rect 454650 399786 454678 400044
rect 416010 399758 416084 399786
rect 408880 396778 408908 399758
rect 411456 398818 411484 399758
rect 411444 398812 411496 398818
rect 411444 398754 411496 398760
rect 408868 396772 408920 396778
rect 408868 396714 408920 396720
rect 414032 395418 414060 399758
rect 414112 396772 414164 396778
rect 414112 396714 414164 396720
rect 414020 395412 414072 395418
rect 414020 395354 414072 395360
rect 405740 392760 405792 392766
rect 405740 392702 405792 392708
rect 409788 389836 409840 389842
rect 409788 389778 409840 389784
rect 406384 388476 406436 388482
rect 406384 388418 406436 388424
rect 404360 377528 404412 377534
rect 404360 377470 404412 377476
rect 405004 377528 405056 377534
rect 405004 377470 405056 377476
rect 403624 367192 403676 367198
rect 403624 367134 403676 367140
rect 401600 336048 401652 336054
rect 401600 335990 401652 335996
rect 401612 334014 401640 335990
rect 401600 334008 401652 334014
rect 401600 333950 401652 333956
rect 399484 307828 399536 307834
rect 399484 307770 399536 307776
rect 398840 307148 398892 307154
rect 398840 307090 398892 307096
rect 399496 303754 399524 307770
rect 399484 303748 399536 303754
rect 399484 303690 399536 303696
rect 395344 303680 395396 303686
rect 395344 303622 395396 303628
rect 393596 301028 393648 301034
rect 393596 300970 393648 300976
rect 393964 301028 394016 301034
rect 393964 300970 394016 300976
rect 386524 299934 387734 299962
rect 389192 299934 389666 299962
rect 391216 299934 391598 299962
rect 393608 299948 393636 300970
rect 395356 299962 395384 303622
rect 398104 303612 398156 303618
rect 398104 303554 398156 303560
rect 395356 299934 395462 299962
rect 398116 299948 398144 303554
rect 399496 299962 399524 303690
rect 401612 299962 401640 333950
rect 403636 302598 403664 367134
rect 405016 305114 405044 377470
rect 405004 305108 405056 305114
rect 405004 305050 405056 305056
rect 405016 303618 405044 305050
rect 406396 303890 406424 388418
rect 409800 306374 409828 389778
rect 413284 361752 413336 361758
rect 413284 361694 413336 361700
rect 410522 353424 410578 353433
rect 410522 353359 410578 353368
rect 409616 306346 409828 306374
rect 409616 305046 409644 306346
rect 410536 305658 410564 353359
rect 413296 321706 413324 361694
rect 413284 321700 413336 321706
rect 413284 321642 413336 321648
rect 410524 305652 410576 305658
rect 410524 305594 410576 305600
rect 409604 305040 409656 305046
rect 409604 304982 409656 304988
rect 406384 303884 406436 303890
rect 406384 303826 406436 303832
rect 405004 303612 405056 303618
rect 405004 303554 405056 303560
rect 403624 302592 403676 302598
rect 403624 302534 403676 302540
rect 403636 299962 403664 302534
rect 406396 299962 406424 303826
rect 407672 302252 407724 302258
rect 407672 302194 407724 302200
rect 399496 299934 399970 299962
rect 401612 299934 401902 299962
rect 403636 299934 403834 299962
rect 405858 299934 406424 299962
rect 407684 299948 407712 302194
rect 409616 300966 409644 304982
rect 409604 300960 409656 300966
rect 409604 300902 409656 300908
rect 412364 300960 412416 300966
rect 412364 300902 412416 300908
rect 409616 299948 409644 300902
rect 412376 299554 412404 300902
rect 414124 299962 414152 396714
rect 416056 395350 416084 399758
rect 418172 399758 418614 399786
rect 421116 399758 421190 399786
rect 423692 399758 423766 399786
rect 425624 399758 425698 399786
rect 428200 399758 428274 399786
rect 430592 399758 430850 399786
rect 432064 399758 432782 399786
rect 434732 399758 435358 399786
rect 437492 399758 437934 399786
rect 440252 399758 440510 399786
rect 441632 399758 442442 399786
rect 444392 399758 445018 399786
rect 447152 399758 447594 399786
rect 448532 399758 449526 399786
rect 452028 399758 452102 399786
rect 454604 399758 454678 399786
rect 457226 399786 457254 400044
rect 459158 399786 459186 400044
rect 461734 399786 461762 400044
rect 464310 399786 464338 400044
rect 466242 399786 466270 400044
rect 468818 399786 468846 400044
rect 471394 399786 471422 400044
rect 473970 399786 473998 400044
rect 475902 399838 475930 400044
rect 457226 399758 457300 399786
rect 416044 395344 416096 395350
rect 416044 395286 416096 395292
rect 418172 392698 418200 399758
rect 421010 395448 421066 395457
rect 421010 395383 421066 395392
rect 418160 392692 418212 392698
rect 418160 392634 418212 392640
rect 417424 366376 417476 366382
rect 417424 366318 417476 366324
rect 417436 356046 417464 366318
rect 418804 365016 418856 365022
rect 418804 364958 418856 364964
rect 417424 356040 417476 356046
rect 417424 355982 417476 355988
rect 417436 325694 417464 355982
rect 417436 325666 417648 325694
rect 415584 316056 415636 316062
rect 415584 315998 415636 316004
rect 414032 299948 414152 299962
rect 415596 299962 415624 315998
rect 417620 303822 417648 325666
rect 417608 303816 417660 303822
rect 417608 303758 417660 303764
rect 417620 299962 417648 303758
rect 418816 301510 418844 364958
rect 420184 321700 420236 321706
rect 420184 321642 420236 321648
rect 420196 312662 420224 321642
rect 420184 312656 420236 312662
rect 420184 312598 420236 312604
rect 419540 309800 419592 309806
rect 419540 309742 419592 309748
rect 419552 309126 419580 309742
rect 419540 309120 419592 309126
rect 419540 309062 419592 309068
rect 420184 309120 420236 309126
rect 420184 309062 420236 309068
rect 418804 301504 418856 301510
rect 418804 301446 418856 301452
rect 420196 299962 420224 309062
rect 421024 300830 421052 395383
rect 421116 393990 421144 399758
rect 421104 393984 421156 393990
rect 421104 393926 421156 393932
rect 423692 365974 423720 399758
rect 425624 396778 425652 399758
rect 428200 399022 428228 399758
rect 428188 399016 428240 399022
rect 428188 398958 428240 398964
rect 425612 396772 425664 396778
rect 425612 396714 425664 396720
rect 423680 365968 423732 365974
rect 423680 365910 423732 365916
rect 424324 365968 424376 365974
rect 424324 365910 424376 365916
rect 424336 355366 424364 365910
rect 429844 356720 429896 356726
rect 429844 356662 429896 356668
rect 425704 355428 425756 355434
rect 425704 355370 425756 355376
rect 424324 355360 424376 355366
rect 424324 355302 424376 355308
rect 425716 325694 425744 355370
rect 429108 348424 429160 348430
rect 429108 348366 429160 348372
rect 425716 325666 425928 325694
rect 425900 302530 425928 325666
rect 425888 302524 425940 302530
rect 425888 302466 425940 302472
rect 423864 302320 423916 302326
rect 423864 302262 423916 302268
rect 421012 300824 421064 300830
rect 421012 300766 421064 300772
rect 421840 300824 421892 300830
rect 421840 300766 421892 300772
rect 414032 299934 414138 299948
rect 415596 299934 416544 299962
rect 417620 299934 418002 299962
rect 420026 299934 420224 299962
rect 421852 299962 421880 300766
rect 421852 299948 422064 299962
rect 423876 299948 423904 302262
rect 425900 299962 425928 302466
rect 429120 302462 429148 348366
rect 429856 303958 429884 356662
rect 430592 312594 430620 399758
rect 432064 363662 432092 399758
rect 431960 363656 432012 363662
rect 431960 363598 432012 363604
rect 432052 363656 432104 363662
rect 432052 363598 432104 363604
rect 430580 312588 430632 312594
rect 430580 312530 430632 312536
rect 429844 303952 429896 303958
rect 429844 303894 429896 303900
rect 430304 303952 430356 303958
rect 430304 303894 430356 303900
rect 428372 302456 428424 302462
rect 428372 302398 428424 302404
rect 429108 302456 429160 302462
rect 429108 302398 429160 302404
rect 421866 299934 422064 299948
rect 425900 299934 426374 299962
rect 428384 299948 428412 302398
rect 430316 299948 430344 303894
rect 431972 299962 432000 363598
rect 434732 322250 434760 399758
rect 434812 394528 434864 394534
rect 434812 394470 434864 394476
rect 434824 387705 434852 394470
rect 434810 387696 434866 387705
rect 434810 387631 434866 387640
rect 437388 351960 437440 351966
rect 437388 351902 437440 351908
rect 434720 322244 434772 322250
rect 434720 322186 434772 322192
rect 437400 309126 437428 351902
rect 437492 347070 437520 399758
rect 440252 386306 440280 399758
rect 440332 398948 440384 398954
rect 440332 398890 440384 398896
rect 440344 398546 440372 398890
rect 440332 398540 440384 398546
rect 440332 398482 440384 398488
rect 440516 387864 440568 387870
rect 440516 387806 440568 387812
rect 440240 386300 440292 386306
rect 440240 386242 440292 386248
rect 440332 365084 440384 365090
rect 440332 365026 440384 365032
rect 438860 351212 438912 351218
rect 438860 351154 438912 351160
rect 438872 350538 438900 351154
rect 438860 350532 438912 350538
rect 438860 350474 438912 350480
rect 440148 350532 440200 350538
rect 440148 350474 440200 350480
rect 437480 347064 437532 347070
rect 437480 347006 437532 347012
rect 438768 322244 438820 322250
rect 438768 322186 438820 322192
rect 436928 309120 436980 309126
rect 436928 309062 436980 309068
rect 437388 309120 437440 309126
rect 437388 309062 437440 309068
rect 436940 308514 436968 309062
rect 436928 308508 436980 308514
rect 436928 308450 436980 308456
rect 434168 307828 434220 307834
rect 434168 307770 434220 307776
rect 431972 299934 432170 299962
rect 434180 299948 434208 307770
rect 438780 306374 438808 322186
rect 438504 306346 438808 306374
rect 438504 300898 438532 306346
rect 440160 302394 440188 350474
rect 440240 329112 440292 329118
rect 440240 329054 440292 329060
rect 440252 328438 440280 329054
rect 440240 328432 440292 328438
rect 440240 328374 440292 328380
rect 440148 302388 440200 302394
rect 440148 302330 440200 302336
rect 436008 300892 436060 300898
rect 436008 300834 436060 300840
rect 438492 300892 438544 300898
rect 438492 300834 438544 300840
rect 436020 299948 436048 300834
rect 438504 299962 438532 300834
rect 440160 299962 440188 302330
rect 438058 299934 438532 299962
rect 439990 299934 440188 299962
rect 414032 299606 414060 299934
rect 416516 299674 416544 299934
rect 416504 299668 416556 299674
rect 416504 299610 416556 299616
rect 422036 299606 422064 299934
rect 438860 299668 438912 299674
rect 438860 299610 438912 299616
rect 411824 299538 412404 299554
rect 414020 299600 414072 299606
rect 422024 299600 422076 299606
rect 414072 299548 414520 299554
rect 414020 299542 414520 299548
rect 422024 299542 422076 299548
rect 411812 299532 412404 299538
rect 411864 299526 412404 299532
rect 414032 299538 414520 299542
rect 414032 299532 414532 299538
rect 414032 299526 414480 299532
rect 411812 299474 411864 299480
rect 414480 299474 414532 299480
rect 438872 299470 438900 299610
rect 438860 299464 438912 299470
rect 438860 299406 438912 299412
rect 379610 299296 379666 299305
rect 379610 299231 379666 299240
rect 440344 291145 440372 365026
rect 440330 291136 440386 291145
rect 440330 291071 440386 291080
rect 440344 289882 440372 291071
rect 440332 289876 440384 289882
rect 440332 289818 440384 289824
rect 440422 288824 440478 288833
rect 440422 288759 440478 288768
rect 379518 276040 379574 276049
rect 379518 275975 379574 275984
rect 440330 276040 440386 276049
rect 440330 275975 440386 275984
rect 379426 274000 379482 274009
rect 379426 273935 379482 273944
rect 379334 261216 379390 261225
rect 379334 261151 379390 261160
rect 379348 260914 379376 261151
rect 379336 260908 379388 260914
rect 379336 260850 379388 260856
rect 379348 258074 379376 260850
rect 440240 259412 440292 259418
rect 440240 259354 440292 259360
rect 440252 259185 440280 259354
rect 440238 259176 440294 259185
rect 440238 259111 440294 259120
rect 379348 258046 379468 258074
rect 379244 228472 379296 228478
rect 379244 228414 379296 228420
rect 378968 216640 379020 216646
rect 378968 216582 379020 216588
rect 378876 145036 378928 145042
rect 378876 144978 378928 144984
rect 378784 110424 378836 110430
rect 378784 110366 378836 110372
rect 378048 95328 378100 95334
rect 378048 95270 378100 95276
rect 378888 25566 378916 144978
rect 378980 104854 379008 216582
rect 379440 149802 379468 258046
rect 379888 256760 379940 256766
rect 379888 256702 379940 256708
rect 379900 248414 379928 256702
rect 379624 248386 379928 248414
rect 379624 238814 379652 248386
rect 379702 242312 379758 242321
rect 379702 242247 379758 242256
rect 379716 240530 379744 242247
rect 381544 240712 381596 240718
rect 381544 240654 381596 240660
rect 381634 240680 381690 240689
rect 379716 240502 380848 240530
rect 379612 238808 379664 238814
rect 379612 238750 379664 238756
rect 380820 218754 380848 240502
rect 380164 218748 380216 218754
rect 380164 218690 380216 218696
rect 380808 218748 380860 218754
rect 380808 218690 380860 218696
rect 379428 149796 379480 149802
rect 379428 149738 379480 149744
rect 380176 117298 380204 218690
rect 381556 203590 381584 240654
rect 381690 240638 381938 240666
rect 381634 240615 381690 240624
rect 381832 240122 381860 240638
rect 382278 240272 382334 240281
rect 382278 240207 382334 240216
rect 381832 240108 382030 240122
rect 381832 240094 382044 240108
rect 382016 232626 382044 240094
rect 382188 239488 382240 239494
rect 382188 239430 382240 239436
rect 382096 239420 382148 239426
rect 382096 239362 382148 239368
rect 382108 238950 382136 239362
rect 382200 239154 382228 239430
rect 382188 239148 382240 239154
rect 382188 239090 382240 239096
rect 382096 238944 382148 238950
rect 382096 238886 382148 238892
rect 382004 232620 382056 232626
rect 382004 232562 382056 232568
rect 381544 203584 381596 203590
rect 381544 203526 381596 203532
rect 381544 146464 381596 146470
rect 381544 146406 381596 146412
rect 380164 117292 380216 117298
rect 380164 117234 380216 117240
rect 378968 104848 379020 104854
rect 378968 104790 379020 104796
rect 381556 54602 381584 146406
rect 382108 103494 382136 238886
rect 382096 103488 382148 103494
rect 382096 103430 382148 103436
rect 382200 92478 382228 239090
rect 382292 233102 382320 240207
rect 383962 240094 384344 240122
rect 384316 238474 384344 240094
rect 384304 238468 384356 238474
rect 384304 238410 384356 238416
rect 383014 236056 383070 236065
rect 383014 235991 383070 236000
rect 382280 233096 382332 233102
rect 382280 233038 382332 233044
rect 382924 212424 382976 212430
rect 382924 212366 382976 212372
rect 382936 93566 382964 212366
rect 383028 120086 383056 235991
rect 384316 171834 384344 238410
rect 385880 233306 385908 240108
rect 387260 240094 387734 240122
rect 389758 240094 389864 240122
rect 387260 238678 387288 240094
rect 387248 238672 387300 238678
rect 387248 238614 387300 238620
rect 387064 233980 387116 233986
rect 387064 233922 387116 233928
rect 385868 233300 385920 233306
rect 385868 233242 385920 233248
rect 385880 219434 385908 233242
rect 386328 229832 386380 229838
rect 386328 229774 386380 229780
rect 385696 219406 385908 219434
rect 385696 218006 385724 219406
rect 385684 218000 385736 218006
rect 385684 217942 385736 217948
rect 384304 171828 384356 171834
rect 384304 171770 384356 171776
rect 385696 129742 385724 217942
rect 385684 129736 385736 129742
rect 385684 129678 385736 129684
rect 385684 127628 385736 127634
rect 385684 127570 385736 127576
rect 383016 120080 383068 120086
rect 383016 120022 383068 120028
rect 382924 93560 382976 93566
rect 382924 93502 382976 93508
rect 382188 92472 382240 92478
rect 382188 92414 382240 92420
rect 381544 54596 381596 54602
rect 381544 54538 381596 54544
rect 378876 25560 378928 25566
rect 378876 25502 378928 25508
rect 377404 17332 377456 17338
rect 377404 17274 377456 17280
rect 385696 15162 385724 127570
rect 386340 92274 386368 229774
rect 387076 111790 387104 233922
rect 387156 232552 387208 232558
rect 387156 232494 387208 232500
rect 387168 134570 387196 232494
rect 387260 149734 387288 238614
rect 389836 237969 389864 240094
rect 391308 240094 391598 240122
rect 390468 239080 390520 239086
rect 390468 239022 390520 239028
rect 390480 238950 390508 239022
rect 390468 238944 390520 238950
rect 390468 238886 390520 238892
rect 389822 237960 389878 237969
rect 389822 237895 389878 237904
rect 388444 232620 388496 232626
rect 388444 232562 388496 232568
rect 387248 149728 387300 149734
rect 387248 149670 387300 149676
rect 387248 148436 387300 148442
rect 387248 148378 387300 148384
rect 387156 134564 387208 134570
rect 387156 134506 387208 134512
rect 387156 113824 387208 113830
rect 387156 113766 387208 113772
rect 387064 111784 387116 111790
rect 387064 111726 387116 111732
rect 387168 93770 387196 113766
rect 387260 93838 387288 148378
rect 388456 102134 388484 232562
rect 388628 218816 388680 218822
rect 388628 218758 388680 218764
rect 388640 218074 388668 218758
rect 388628 218068 388680 218074
rect 388628 218010 388680 218016
rect 389088 218068 389140 218074
rect 389088 218010 389140 218016
rect 389100 170406 389128 218010
rect 389836 182850 389864 237895
rect 390376 193860 390428 193866
rect 390376 193802 390428 193808
rect 389824 182844 389876 182850
rect 389824 182786 389876 182792
rect 389088 170400 389140 170406
rect 389088 170342 389140 170348
rect 390388 142154 390416 193802
rect 390204 142126 390416 142154
rect 390204 136649 390232 142126
rect 390190 136640 390246 136649
rect 390190 136575 390246 136584
rect 390204 135318 390232 136575
rect 390192 135312 390244 135318
rect 390192 135254 390244 135260
rect 390480 111722 390508 238886
rect 391308 235686 391336 240094
rect 393608 238542 393636 240108
rect 395988 239556 396040 239562
rect 395988 239498 396040 239504
rect 396000 238882 396028 239498
rect 395988 238876 396040 238882
rect 395988 238818 396040 238824
rect 393596 238536 393648 238542
rect 393596 238478 393648 238484
rect 392584 236700 392636 236706
rect 392584 236642 392636 236648
rect 391296 235680 391348 235686
rect 391296 235622 391348 235628
rect 391204 231260 391256 231266
rect 391204 231202 391256 231208
rect 390468 111716 390520 111722
rect 390468 111658 390520 111664
rect 388444 102128 388496 102134
rect 388444 102070 388496 102076
rect 387248 93832 387300 93838
rect 387248 93774 387300 93780
rect 387156 93764 387208 93770
rect 387156 93706 387208 93712
rect 391216 93702 391244 231202
rect 391308 193934 391336 235622
rect 391848 213240 391900 213246
rect 391848 213182 391900 213188
rect 391296 193928 391348 193934
rect 391296 193870 391348 193876
rect 391860 137902 391888 213182
rect 392596 147014 392624 236642
rect 393608 236026 393636 238478
rect 394608 236768 394660 236774
rect 394608 236710 394660 236716
rect 393596 236020 393648 236026
rect 393596 235962 393648 235968
rect 393228 220108 393280 220114
rect 393228 220050 393280 220056
rect 392676 181484 392728 181490
rect 392676 181426 392728 181432
rect 392584 147008 392636 147014
rect 392584 146950 392636 146956
rect 391848 137896 391900 137902
rect 391848 137838 391900 137844
rect 391940 135312 391992 135318
rect 391940 135254 391992 135260
rect 391296 132592 391348 132598
rect 391296 132534 391348 132540
rect 391204 93696 391256 93702
rect 391204 93638 391256 93644
rect 386328 92268 386380 92274
rect 386328 92210 386380 92216
rect 391308 28966 391336 132534
rect 391952 98666 391980 135254
rect 392584 132524 392636 132530
rect 392584 132466 392636 132472
rect 391940 98660 391992 98666
rect 391940 98602 391992 98608
rect 391296 28960 391348 28966
rect 391296 28902 391348 28908
rect 392596 22098 392624 132466
rect 392688 128314 392716 181426
rect 392676 128308 392728 128314
rect 392676 128250 392728 128256
rect 393240 102066 393268 220050
rect 393964 179444 394016 179450
rect 393964 179386 394016 179392
rect 393228 102060 393280 102066
rect 393228 102002 393280 102008
rect 393976 93634 394004 179386
rect 394056 134700 394108 134706
rect 394056 134642 394108 134648
rect 394068 101454 394096 134642
rect 394620 132598 394648 236710
rect 395344 236020 395396 236026
rect 395344 235962 395396 235968
rect 394608 132592 394660 132598
rect 394608 132534 394660 132540
rect 395356 122330 395384 235962
rect 395896 202156 395948 202162
rect 395896 202098 395948 202104
rect 395804 146940 395856 146946
rect 395804 146882 395856 146888
rect 395436 123276 395488 123282
rect 395436 123218 395488 123224
rect 395344 122324 395396 122330
rect 395344 122266 395396 122272
rect 395344 109064 395396 109070
rect 395344 109006 395396 109012
rect 394056 101448 394108 101454
rect 394056 101390 394108 101396
rect 393964 93628 394016 93634
rect 393964 93570 394016 93576
rect 392584 22092 392636 22098
rect 392584 22034 392636 22040
rect 385684 15156 385736 15162
rect 385684 15098 385736 15104
rect 360936 13796 360988 13802
rect 360936 13738 360988 13744
rect 356796 8220 356848 8226
rect 356796 8162 356848 8168
rect 395356 4826 395384 109006
rect 395448 53786 395476 123218
rect 395816 94858 395844 146882
rect 395908 129878 395936 202098
rect 395896 129872 395948 129878
rect 395896 129814 395948 129820
rect 396000 113150 396028 238818
rect 396092 230450 396120 240108
rect 398116 235890 398144 240108
rect 399956 238814 399984 240108
rect 401994 240094 402284 240122
rect 398932 238808 398984 238814
rect 398932 238750 398984 238756
rect 399944 238808 399996 238814
rect 399944 238750 399996 238756
rect 398104 235884 398156 235890
rect 398104 235826 398156 235832
rect 397368 235272 397420 235278
rect 397368 235214 397420 235220
rect 396080 230444 396132 230450
rect 396080 230386 396132 230392
rect 396092 230042 396120 230386
rect 396080 230036 396132 230042
rect 396080 229978 396132 229984
rect 396724 230036 396776 230042
rect 396724 229978 396776 229984
rect 396080 191140 396132 191146
rect 396080 191082 396132 191088
rect 396092 134706 396120 191082
rect 396736 176118 396764 229978
rect 396724 176112 396776 176118
rect 396724 176054 396776 176060
rect 396816 147824 396868 147830
rect 396816 147766 396868 147772
rect 396080 134700 396132 134706
rect 396080 134642 396132 134648
rect 396722 119096 396778 119105
rect 396722 119031 396778 119040
rect 395988 113144 396040 113150
rect 395988 113086 396040 113092
rect 395804 94852 395856 94858
rect 395804 94794 395856 94800
rect 395436 53780 395488 53786
rect 395436 53722 395488 53728
rect 396736 19310 396764 119031
rect 396828 71126 396856 147766
rect 397380 140321 397408 235214
rect 398116 191826 398144 235826
rect 398944 209166 398972 238750
rect 402256 235754 402284 240094
rect 403820 237182 403848 240108
rect 405752 238754 405780 240108
rect 405660 238726 405780 238754
rect 405660 238066 405688 238726
rect 407776 238610 407804 240108
rect 410366 240094 410564 240122
rect 407764 238604 407816 238610
rect 407764 238546 407816 238552
rect 405648 238060 405700 238066
rect 405648 238002 405700 238008
rect 402980 237176 403032 237182
rect 402980 237118 403032 237124
rect 403808 237176 403860 237182
rect 403808 237118 403860 237124
rect 402244 235748 402296 235754
rect 402244 235690 402296 235696
rect 399116 227044 399168 227050
rect 399116 226986 399168 226992
rect 398932 209160 398984 209166
rect 398932 209102 398984 209108
rect 398104 191820 398156 191826
rect 398104 191762 398156 191768
rect 398746 180024 398802 180033
rect 398746 179959 398802 179968
rect 398102 174584 398158 174593
rect 398102 174519 398158 174528
rect 398116 151814 398144 174519
rect 398656 160744 398708 160750
rect 398656 160686 398708 160692
rect 398116 151786 398236 151814
rect 397552 149796 397604 149802
rect 397552 149738 397604 149744
rect 397458 145616 397514 145625
rect 397458 145551 397514 145560
rect 397472 145110 397500 145551
rect 397460 145104 397512 145110
rect 397460 145046 397512 145052
rect 397460 144288 397512 144294
rect 397458 144256 397460 144265
rect 397512 144256 397514 144265
rect 397458 144191 397514 144200
rect 397564 143721 397592 149738
rect 397550 143712 397606 143721
rect 397550 143647 397606 143656
rect 397550 142216 397606 142225
rect 397550 142151 397552 142160
rect 397604 142151 397606 142160
rect 397552 142122 397604 142128
rect 397460 142112 397512 142118
rect 397460 142054 397512 142060
rect 397472 141681 397500 142054
rect 397458 141672 397514 141681
rect 397458 141607 397514 141616
rect 397366 140312 397422 140321
rect 397366 140247 397422 140256
rect 397460 139392 397512 139398
rect 397460 139334 397512 139340
rect 397472 138961 397500 139334
rect 397458 138952 397514 138961
rect 397458 138887 397514 138896
rect 397552 137964 397604 137970
rect 397552 137906 397604 137912
rect 397460 137896 397512 137902
rect 397460 137838 397512 137844
rect 397472 137601 397500 137838
rect 397458 137592 397514 137601
rect 397458 137527 397514 137536
rect 397564 136921 397592 137906
rect 397550 136912 397606 136921
rect 397550 136847 397606 136856
rect 397458 135416 397514 135425
rect 397458 135351 397514 135360
rect 397472 135318 397500 135351
rect 397460 135312 397512 135318
rect 397460 135254 397512 135260
rect 397458 134736 397514 134745
rect 397458 134671 397460 134680
rect 397512 134671 397514 134680
rect 397460 134642 397512 134648
rect 397458 133376 397514 133385
rect 397458 133311 397514 133320
rect 397472 132530 397500 133311
rect 397550 132696 397606 132705
rect 397550 132631 397606 132640
rect 397564 132598 397592 132631
rect 397552 132592 397604 132598
rect 397552 132534 397604 132540
rect 397460 132524 397512 132530
rect 397460 132466 397512 132472
rect 397550 130656 397606 130665
rect 397550 130591 397606 130600
rect 397458 129976 397514 129985
rect 397380 129934 397458 129962
rect 397380 123486 397408 129934
rect 397458 129911 397514 129920
rect 397564 129810 397592 130591
rect 398208 129985 398236 151786
rect 398194 129976 398250 129985
rect 398194 129911 398250 129920
rect 398288 129872 398340 129878
rect 398288 129814 398340 129820
rect 397552 129804 397604 129810
rect 397552 129746 397604 129752
rect 397460 129736 397512 129742
rect 397460 129678 397512 129684
rect 397472 128761 397500 129678
rect 397458 128752 397514 128761
rect 397458 128687 397514 128696
rect 397458 127936 397514 127945
rect 397458 127871 397514 127880
rect 397472 127634 397500 127871
rect 397460 127628 397512 127634
rect 397460 127570 397512 127576
rect 397552 126948 397604 126954
rect 397552 126890 397604 126896
rect 397460 126880 397512 126886
rect 397460 126822 397512 126828
rect 397472 126721 397500 126822
rect 397458 126712 397514 126721
rect 397458 126647 397514 126656
rect 397564 126041 397592 126890
rect 397550 126032 397606 126041
rect 397550 125967 397606 125976
rect 397460 125588 397512 125594
rect 397460 125530 397512 125536
rect 397472 125361 397500 125530
rect 397458 125352 397514 125361
rect 397458 125287 397514 125296
rect 397458 123856 397514 123865
rect 397458 123791 397514 123800
rect 397368 123480 397420 123486
rect 397368 123422 397420 123428
rect 397472 123282 397500 123791
rect 397460 123276 397512 123282
rect 397460 123218 397512 123224
rect 398194 123176 398250 123185
rect 398194 123111 398250 123120
rect 397460 122324 397512 122330
rect 397460 122266 397512 122272
rect 397472 121961 397500 122266
rect 397458 121952 397514 121961
rect 397458 121887 397514 121896
rect 397460 121440 397512 121446
rect 397460 121382 397512 121388
rect 397472 121281 397500 121382
rect 397458 121272 397514 121281
rect 397458 121207 397514 121216
rect 397460 120080 397512 120086
rect 397460 120022 397512 120028
rect 397472 119921 397500 120022
rect 397458 119912 397514 119921
rect 397458 119847 397514 119856
rect 397460 117292 397512 117298
rect 397460 117234 397512 117240
rect 397472 117201 397500 117234
rect 397458 117192 397514 117201
rect 397458 117127 397514 117136
rect 397460 115932 397512 115938
rect 397460 115874 397512 115880
rect 397472 115161 397500 115874
rect 397458 115152 397514 115161
rect 397458 115087 397514 115096
rect 397460 114504 397512 114510
rect 397458 114472 397460 114481
rect 397512 114472 397514 114481
rect 397458 114407 397514 114416
rect 397460 113144 397512 113150
rect 397458 113112 397460 113121
rect 397512 113112 397514 113121
rect 397458 113047 397514 113056
rect 397460 111784 397512 111790
rect 397460 111726 397512 111732
rect 397472 111081 397500 111726
rect 397552 111104 397604 111110
rect 397458 111072 397514 111081
rect 397552 111046 397604 111052
rect 397458 111007 397514 111016
rect 397460 110424 397512 110430
rect 397458 110392 397460 110401
rect 397512 110392 397514 110401
rect 397458 110327 397514 110336
rect 397458 108216 397514 108225
rect 397458 108151 397514 108160
rect 397472 107710 397500 108151
rect 397460 107704 397512 107710
rect 397460 107646 397512 107652
rect 397458 105632 397514 105641
rect 397564 105618 397592 111046
rect 397734 109576 397790 109585
rect 397734 109511 397790 109520
rect 397748 109070 397776 109511
rect 397736 109064 397788 109070
rect 397736 109006 397788 109012
rect 397644 106956 397696 106962
rect 397644 106898 397696 106904
rect 397656 106321 397684 106898
rect 397642 106312 397698 106321
rect 397642 106247 397698 106256
rect 397514 105590 397592 105618
rect 397458 105567 397460 105576
rect 397512 105567 397514 105576
rect 397460 105538 397512 105544
rect 397656 105482 397684 106247
rect 397472 105454 397684 105482
rect 396906 96656 396962 96665
rect 396906 96591 396962 96600
rect 396816 71120 396868 71126
rect 396816 71062 396868 71068
rect 396920 31754 396948 96591
rect 397472 89010 397500 105454
rect 397552 104848 397604 104854
rect 397552 104790 397604 104796
rect 397564 103601 397592 104790
rect 398010 104136 398066 104145
rect 398010 104071 398066 104080
rect 397550 103592 397606 103601
rect 397550 103527 397606 103536
rect 397552 103488 397604 103494
rect 397552 103430 397604 103436
rect 397564 102921 397592 103430
rect 397550 102912 397606 102921
rect 397550 102847 397606 102856
rect 397552 102128 397604 102134
rect 397552 102070 397604 102076
rect 397564 101561 397592 102070
rect 397644 102060 397696 102066
rect 397644 102002 397696 102008
rect 397550 101552 397606 101561
rect 397550 101487 397606 101496
rect 397656 100881 397684 102002
rect 397642 100872 397698 100881
rect 397642 100807 397698 100816
rect 397552 100020 397604 100026
rect 397552 99962 397604 99968
rect 397564 99521 397592 99962
rect 397550 99512 397606 99521
rect 397550 99447 397606 99456
rect 397550 97336 397606 97345
rect 397550 97271 397606 97280
rect 397564 96694 397592 97271
rect 397552 96688 397604 96694
rect 397552 96630 397604 96636
rect 398024 93854 398052 104071
rect 398024 93826 398144 93854
rect 397460 89004 397512 89010
rect 397460 88946 397512 88952
rect 398116 46918 398144 93826
rect 398208 90982 398236 123111
rect 398300 117881 398328 129814
rect 398668 127945 398696 160686
rect 398760 132161 398788 179959
rect 398932 152652 398984 152658
rect 398932 152594 398984 152600
rect 398746 132152 398802 132161
rect 398746 132087 398802 132096
rect 398760 131782 398788 132087
rect 398748 131776 398800 131782
rect 398748 131718 398800 131724
rect 398654 127936 398710 127945
rect 398654 127871 398710 127880
rect 398286 117872 398342 117881
rect 398286 117807 398342 117816
rect 398944 116521 398972 152594
rect 399024 134564 399076 134570
rect 399024 134506 399076 134512
rect 398930 116512 398986 116521
rect 398930 116447 398986 116456
rect 399036 97850 399064 134506
rect 399128 98841 399156 226986
rect 402256 192574 402284 235690
rect 402244 192568 402296 192574
rect 402244 192510 402296 192516
rect 399484 191820 399536 191826
rect 399484 191762 399536 191768
rect 399114 98832 399170 98841
rect 399114 98767 399170 98776
rect 399024 97844 399076 97850
rect 399024 97786 399076 97792
rect 398196 90976 398248 90982
rect 398196 90918 398248 90924
rect 399036 84194 399064 97786
rect 399496 93838 399524 191762
rect 401600 169108 401652 169114
rect 401600 169050 401652 169056
rect 400220 152516 400272 152522
rect 400220 152458 400272 152464
rect 400232 151814 400260 152458
rect 400232 151786 400536 151814
rect 400036 148368 400088 148374
rect 400036 148310 400088 148316
rect 400048 145860 400076 148310
rect 400128 147008 400180 147014
rect 400128 146950 400180 146956
rect 400140 146334 400168 146950
rect 400128 146328 400180 146334
rect 400128 146270 400180 146276
rect 399852 145444 399904 145450
rect 399852 145386 399904 145392
rect 399864 144974 399892 145386
rect 399852 144968 399904 144974
rect 399852 144910 399904 144916
rect 400140 140049 400168 146270
rect 400508 145466 400536 151786
rect 401612 145874 401640 169050
rect 402612 148028 402664 148034
rect 402612 147970 402664 147976
rect 401612 145846 401994 145874
rect 402624 145860 402652 147970
rect 402992 146946 403020 237118
rect 404360 213308 404412 213314
rect 404360 213250 404412 213256
rect 403624 180124 403676 180130
rect 403624 180066 403676 180072
rect 403636 148034 403664 180066
rect 403624 148028 403676 148034
rect 403624 147970 403676 147976
rect 402980 146940 403032 146946
rect 402980 146882 403032 146888
rect 404372 145874 404400 213250
rect 405660 152522 405688 238002
rect 405740 204944 405792 204950
rect 405740 204886 405792 204892
rect 405648 152516 405700 152522
rect 405648 152458 405700 152464
rect 405752 151814 405780 204886
rect 407776 191146 407804 238546
rect 408500 233912 408552 233918
rect 408500 233854 408552 233860
rect 407764 191140 407816 191146
rect 407764 191082 407816 191088
rect 408512 171134 408540 233854
rect 410536 233034 410564 240094
rect 411916 240094 412206 240122
rect 411916 237318 411944 240094
rect 411904 237312 411956 237318
rect 411904 237254 411956 237260
rect 410524 233028 410576 233034
rect 410524 232970 410576 232976
rect 409880 228472 409932 228478
rect 409880 228414 409932 228420
rect 408512 171106 408632 171134
rect 407764 169040 407816 169046
rect 407764 168982 407816 168988
rect 405752 151786 405872 151814
rect 405844 147830 405872 151786
rect 406476 151156 406528 151162
rect 406476 151098 406528 151104
rect 405832 147824 405884 147830
rect 405832 147766 405884 147772
rect 404372 145846 404570 145874
rect 405844 145860 405872 147766
rect 406488 145860 406516 151098
rect 407776 146470 407804 168982
rect 408408 153876 408460 153882
rect 408408 153818 408460 153824
rect 407764 146464 407816 146470
rect 407764 146406 407816 146412
rect 407776 145860 407804 146406
rect 408420 145860 408448 153818
rect 408604 145874 408632 171106
rect 409892 148578 409920 228414
rect 409972 176112 410024 176118
rect 409972 176054 410024 176060
rect 409880 148572 409932 148578
rect 409880 148514 409932 148520
rect 409984 145874 410012 176054
rect 410536 163538 410564 232970
rect 410524 163532 410576 163538
rect 410524 163474 410576 163480
rect 411916 156670 411944 237254
rect 414020 236836 414072 236842
rect 414020 236778 414072 236784
rect 412640 166320 412692 166326
rect 412640 166262 412692 166268
rect 411904 156664 411956 156670
rect 411904 156606 411956 156612
rect 412272 151088 412324 151094
rect 412272 151030 412324 151036
rect 410708 148572 410760 148578
rect 410708 148514 410760 148520
rect 410720 145874 410748 148514
rect 408604 145846 409078 145874
rect 409984 145846 410366 145874
rect 410720 145846 411010 145874
rect 412284 145860 412312 151030
rect 412652 145874 412680 166262
rect 414032 145874 414060 236778
rect 414216 220114 414244 240108
rect 415412 240094 416070 240122
rect 417436 240094 418002 240122
rect 420026 240094 420224 240122
rect 414294 226944 414350 226953
rect 414294 226879 414350 226888
rect 414204 220108 414256 220114
rect 414204 220050 414256 220056
rect 414308 171134 414336 226879
rect 415412 226302 415440 240094
rect 417436 238377 417464 240094
rect 420196 238678 420224 240094
rect 420932 240094 421866 240122
rect 424336 240094 424442 240122
rect 420184 238672 420236 238678
rect 420184 238614 420236 238620
rect 417422 238368 417478 238377
rect 417422 238303 417478 238312
rect 415400 226296 415452 226302
rect 415400 226238 415452 226244
rect 416964 192500 417016 192506
rect 416964 192442 417016 192448
rect 416872 187060 416924 187066
rect 416872 187002 416924 187008
rect 414308 171106 414520 171134
rect 414492 145874 414520 171106
rect 415400 167680 415452 167686
rect 415400 167622 415452 167628
rect 415412 151814 415440 167622
rect 415412 151786 415532 151814
rect 412652 145846 412942 145874
rect 414032 145846 414230 145874
rect 414492 145846 414874 145874
rect 415504 145860 415532 151786
rect 416884 147694 416912 187002
rect 416976 171134 417004 192442
rect 417436 186998 417464 238303
rect 418804 229764 418856 229770
rect 418804 229706 418856 229712
rect 417424 186992 417476 186998
rect 417424 186934 417476 186940
rect 418816 171134 418844 229706
rect 419448 217320 419500 217326
rect 419448 217262 419500 217268
rect 416976 171106 417096 171134
rect 418816 171106 418936 171134
rect 416872 147688 416924 147694
rect 416872 147630 416924 147636
rect 416884 145874 416912 147630
rect 416806 145846 416912 145874
rect 417068 145874 417096 171106
rect 418712 152584 418764 152590
rect 418712 152526 418764 152532
rect 417068 145846 417450 145874
rect 418724 145860 418752 152526
rect 418908 147762 418936 171106
rect 419460 148510 419488 217262
rect 420196 152658 420224 238614
rect 420932 219366 420960 240094
rect 424336 238746 424364 240094
rect 424324 238740 424376 238746
rect 424324 238682 424376 238688
rect 422300 237720 422352 237726
rect 422300 237662 422352 237668
rect 422312 237250 422340 237662
rect 422300 237244 422352 237250
rect 422300 237186 422352 237192
rect 420920 219360 420972 219366
rect 420920 219302 420972 219308
rect 420932 218142 420960 219302
rect 420920 218136 420972 218142
rect 420920 218078 420972 218084
rect 421656 218136 421708 218142
rect 421656 218078 421708 218084
rect 421564 204944 421616 204950
rect 421564 204886 421616 204892
rect 420276 189848 420328 189854
rect 420276 189790 420328 189796
rect 420184 152652 420236 152658
rect 420184 152594 420236 152600
rect 420288 149122 420316 189790
rect 420276 149116 420328 149122
rect 420276 149058 420328 149064
rect 419448 148504 419500 148510
rect 419448 148446 419500 148452
rect 418896 147756 418948 147762
rect 418896 147698 418948 147704
rect 418908 145874 418936 147698
rect 420288 145874 420316 149058
rect 421288 148504 421340 148510
rect 421288 148446 421340 148452
rect 418908 145846 419382 145874
rect 420288 145846 420670 145874
rect 421300 145860 421328 148446
rect 421576 147626 421604 204886
rect 421668 201550 421696 218078
rect 421656 201544 421708 201550
rect 421656 201486 421708 201492
rect 422208 201544 422260 201550
rect 422208 201486 422260 201492
rect 421564 147620 421616 147626
rect 421564 147562 421616 147568
rect 421932 147620 421984 147626
rect 421932 147562 421984 147568
rect 421944 145860 421972 147562
rect 422220 146985 422248 201486
rect 422312 169114 422340 237186
rect 423588 215960 423640 215966
rect 423588 215902 423640 215908
rect 422760 170400 422812 170406
rect 422760 170342 422812 170348
rect 422300 169108 422352 169114
rect 422300 169050 422352 169056
rect 422206 146976 422262 146985
rect 422206 146911 422262 146920
rect 422772 145874 422800 170342
rect 423600 145874 423628 215902
rect 424336 159458 424364 238682
rect 426360 237726 426388 240108
rect 427924 240094 428306 240122
rect 429212 240094 430238 240122
rect 427924 238785 427952 240094
rect 427910 238776 427966 238785
rect 427910 238711 427966 238720
rect 426348 237720 426400 237726
rect 426348 237662 426400 237668
rect 426440 236904 426492 236910
rect 426440 236846 426492 236852
rect 424324 159452 424376 159458
rect 424324 159394 424376 159400
rect 425796 152584 425848 152590
rect 425796 152526 425848 152532
rect 425152 148368 425204 148374
rect 425152 148310 425204 148316
rect 422772 145846 423246 145874
rect 423600 145846 423890 145874
rect 425164 145860 425192 148310
rect 425808 145860 425836 152526
rect 426452 148578 426480 236846
rect 426624 231124 426676 231130
rect 426624 231066 426676 231072
rect 426532 164892 426584 164898
rect 426532 164834 426584 164840
rect 426544 151814 426572 164834
rect 426636 153882 426664 231066
rect 427924 219434 427952 238711
rect 429108 236972 429160 236978
rect 429108 236914 429160 236920
rect 427832 219406 427952 219434
rect 427084 201544 427136 201550
rect 427084 201486 427136 201492
rect 427096 193186 427124 201486
rect 427084 193180 427136 193186
rect 427084 193122 427136 193128
rect 427832 180130 427860 219406
rect 427820 180124 427872 180130
rect 427820 180066 427872 180072
rect 428464 176044 428516 176050
rect 428464 175986 428516 175992
rect 426624 153876 426676 153882
rect 426624 153818 426676 153824
rect 426544 151786 426664 151814
rect 426440 148572 426492 148578
rect 426440 148514 426492 148520
rect 426636 145874 426664 151786
rect 427452 148572 427504 148578
rect 427452 148514 427504 148520
rect 427464 145874 427492 148514
rect 428476 148442 428504 175986
rect 428464 148436 428516 148442
rect 428464 148378 428516 148384
rect 429120 147694 429148 236914
rect 429212 213246 429240 240094
rect 432248 238066 432276 240108
rect 432236 238060 432288 238066
rect 432236 238002 432288 238008
rect 434088 237454 434116 240108
rect 434732 240094 436034 240122
rect 432696 237448 432748 237454
rect 432696 237390 432748 237396
rect 434076 237448 434128 237454
rect 434076 237390 434128 237396
rect 432604 236700 432656 236706
rect 432604 236642 432656 236648
rect 431960 233164 432012 233170
rect 431960 233106 432012 233112
rect 429200 213240 429252 213246
rect 429200 213182 429252 213188
rect 431224 209092 431276 209098
rect 431224 209034 431276 209040
rect 429200 176792 429252 176798
rect 429200 176734 429252 176740
rect 429212 171134 429240 176734
rect 429212 171106 429976 171134
rect 429660 153264 429712 153270
rect 429660 153206 429712 153212
rect 429108 147688 429160 147694
rect 429108 147630 429160 147636
rect 429120 145874 429148 147630
rect 426636 145846 427110 145874
rect 427464 145846 427754 145874
rect 429042 145846 429148 145874
rect 429672 145860 429700 153206
rect 429948 145874 429976 171106
rect 431236 146946 431264 209034
rect 431316 180872 431368 180878
rect 431316 180814 431368 180820
rect 431328 148782 431356 180814
rect 431592 153332 431644 153338
rect 431592 153274 431644 153280
rect 431316 148776 431368 148782
rect 431316 148718 431368 148724
rect 431224 146940 431276 146946
rect 431224 146882 431276 146888
rect 429948 145846 430330 145874
rect 431604 145860 431632 153274
rect 431972 153270 432000 233106
rect 431960 153264 432012 153270
rect 431960 153206 432012 153212
rect 432616 146402 432644 236642
rect 432708 233170 432736 237390
rect 432696 233164 432748 233170
rect 432696 233106 432748 233112
rect 434732 222154 434760 240094
rect 438596 239018 438624 240108
rect 439504 239692 439556 239698
rect 439504 239634 439556 239640
rect 438858 239456 438914 239465
rect 438858 239391 438914 239400
rect 435364 239012 435416 239018
rect 435364 238954 435416 238960
rect 438584 239012 438636 239018
rect 438584 238954 438636 238960
rect 434720 222148 434772 222154
rect 434720 222090 434772 222096
rect 433984 218748 434036 218754
rect 433984 218690 434036 218696
rect 433996 146402 434024 218690
rect 435376 166326 435404 238954
rect 436744 238808 436796 238814
rect 436744 238750 436796 238756
rect 436008 222148 436060 222154
rect 436008 222090 436060 222096
rect 436020 221474 436048 222090
rect 436008 221468 436060 221474
rect 436008 221410 436060 221416
rect 435456 205012 435508 205018
rect 435456 204954 435508 204960
rect 435364 166320 435416 166326
rect 435364 166262 435416 166268
rect 435468 149054 435496 204954
rect 435548 192568 435600 192574
rect 435548 192510 435600 192516
rect 435456 149048 435508 149054
rect 435456 148990 435508 148996
rect 434168 148776 434220 148782
rect 434168 148718 434220 148724
rect 432604 146396 432656 146402
rect 432604 146338 432656 146344
rect 433524 146396 433576 146402
rect 433524 146338 433576 146344
rect 433984 146396 434036 146402
rect 433984 146338 434036 146344
rect 432616 145874 432644 146338
rect 432262 145846 432644 145874
rect 433536 145860 433564 146338
rect 434180 145860 434208 148718
rect 435456 148436 435508 148442
rect 435456 148378 435508 148384
rect 435468 145860 435496 148378
rect 435560 148306 435588 192510
rect 436284 182844 436336 182850
rect 436284 182786 436336 182792
rect 436296 171134 436324 182786
rect 436296 171106 436416 171134
rect 435548 148300 435600 148306
rect 435548 148242 435600 148248
rect 436100 148232 436152 148238
rect 436100 148174 436152 148180
rect 436112 145860 436140 148174
rect 436388 145874 436416 171106
rect 436756 148374 436784 238750
rect 438596 238746 438624 238954
rect 438872 238950 438900 239391
rect 438860 238944 438912 238950
rect 438860 238886 438912 238892
rect 438584 238740 438636 238746
rect 438584 238682 438636 238688
rect 439516 216034 439544 239634
rect 440252 236978 440280 259111
rect 440240 236972 440292 236978
rect 440240 236914 440292 236920
rect 439504 216028 439556 216034
rect 439504 215970 439556 215976
rect 439504 198008 439556 198014
rect 439504 197950 439556 197956
rect 436744 148368 436796 148374
rect 436744 148310 436796 148316
rect 438032 148300 438084 148306
rect 438032 148242 438084 148248
rect 436388 145846 436770 145874
rect 438044 145860 438072 148242
rect 438676 148164 438728 148170
rect 438676 148106 438728 148112
rect 438688 145860 438716 148106
rect 439516 147801 439544 197950
rect 440240 186992 440292 186998
rect 440240 186934 440292 186940
rect 439596 162172 439648 162178
rect 439596 162114 439648 162120
rect 439608 148170 439636 162114
rect 439596 148164 439648 148170
rect 439596 148106 439648 148112
rect 439502 147792 439558 147801
rect 439502 147727 439558 147736
rect 439962 147792 440018 147801
rect 439962 147727 440018 147736
rect 439976 145860 440004 147727
rect 440252 145874 440280 186934
rect 440344 167686 440372 275975
rect 440436 239562 440464 288759
rect 440528 257145 440556 387806
rect 441632 331906 441660 399758
rect 444392 383654 444420 399758
rect 444392 383626 444512 383654
rect 444484 371890 444512 383626
rect 444472 371884 444524 371890
rect 444472 371826 444524 371832
rect 442172 352572 442224 352578
rect 442172 352514 442224 352520
rect 442184 351898 442212 352514
rect 442172 351892 442224 351898
rect 442172 351834 442224 351840
rect 442908 351892 442960 351898
rect 442908 351834 442960 351840
rect 441620 331900 441672 331906
rect 441620 331842 441672 331848
rect 440884 328432 440936 328438
rect 440884 328374 440936 328380
rect 440896 276049 440924 328374
rect 440976 312656 441028 312662
rect 440976 312598 441028 312604
rect 440988 287065 441016 312598
rect 441712 307080 441764 307086
rect 441712 307022 441764 307028
rect 441620 304292 441672 304298
rect 441620 304234 441672 304240
rect 441528 287088 441580 287094
rect 440974 287056 441030 287065
rect 440974 286991 441030 287000
rect 441526 287056 441528 287065
rect 441580 287056 441582 287065
rect 441526 286991 441582 287000
rect 440882 276040 440938 276049
rect 440882 275975 440938 275984
rect 440514 257136 440570 257145
rect 440514 257071 440570 257080
rect 440528 256766 440556 257071
rect 440516 256760 440568 256766
rect 440516 256702 440568 256708
rect 441632 248169 441660 304234
rect 441724 295089 441752 307022
rect 442814 297120 442870 297129
rect 442814 297055 442870 297064
rect 442828 296954 442856 297055
rect 442816 296948 442868 296954
rect 442816 296890 442868 296896
rect 441710 295080 441766 295089
rect 441710 295015 441766 295024
rect 442814 295080 442870 295089
rect 442814 295015 442870 295024
rect 442828 294642 442856 295015
rect 442816 294636 442868 294642
rect 442816 294578 442868 294584
rect 442172 285660 442224 285666
rect 442172 285602 442224 285608
rect 442184 285025 442212 285602
rect 442170 285016 442226 285025
rect 442170 284951 442226 284960
rect 442722 282160 442778 282169
rect 442722 282095 442778 282104
rect 442736 281858 442764 282095
rect 442724 281852 442776 281858
rect 442724 281794 442776 281800
rect 442814 280256 442870 280265
rect 442814 280191 442816 280200
rect 442868 280191 442870 280200
rect 442816 280162 442868 280168
rect 442630 278080 442686 278089
rect 442630 278015 442686 278024
rect 442644 277438 442672 278015
rect 442632 277432 442684 277438
rect 442632 277374 442684 277380
rect 442722 274000 442778 274009
rect 442722 273935 442778 273944
rect 442736 273290 442764 273935
rect 442724 273284 442776 273290
rect 442724 273226 442776 273232
rect 442816 272128 442868 272134
rect 442814 272096 442816 272105
rect 442868 272096 442870 272105
rect 442814 272031 442870 272040
rect 442262 269920 442318 269929
rect 442262 269855 442318 269864
rect 442276 269142 442304 269855
rect 442264 269136 442316 269142
rect 442264 269078 442316 269084
rect 442814 267200 442870 267209
rect 442814 267135 442870 267144
rect 442828 266422 442856 267135
rect 442816 266416 442868 266422
rect 442816 266358 442868 266364
rect 442354 265160 442410 265169
rect 442354 265095 442356 265104
rect 442408 265095 442410 265104
rect 442356 265066 442408 265072
rect 442722 263120 442778 263129
rect 442722 263055 442778 263064
rect 442736 262274 442764 263055
rect 442724 262268 442776 262274
rect 442724 262210 442776 262216
rect 442816 261520 442868 261526
rect 442816 261462 442868 261468
rect 442828 261225 442856 261462
rect 441710 261216 441766 261225
rect 441710 261151 441766 261160
rect 442814 261216 442870 261225
rect 442814 261151 442870 261160
rect 441618 248160 441674 248169
rect 441618 248095 441674 248104
rect 441632 247081 441660 248095
rect 441618 247072 441674 247081
rect 441618 247007 441674 247016
rect 441618 246256 441674 246265
rect 441618 246191 441674 246200
rect 440424 239556 440476 239562
rect 440424 239498 440476 239504
rect 441632 239426 441660 246191
rect 441724 239494 441752 261151
rect 442920 258074 442948 351834
rect 443092 316736 443144 316742
rect 443092 316678 443144 316684
rect 443000 303884 443052 303890
rect 443000 303826 443052 303832
rect 442736 258046 442948 258074
rect 442736 251258 442764 258046
rect 442906 252376 442962 252385
rect 442906 252311 442962 252320
rect 442920 251870 442948 252311
rect 442908 251864 442960 251870
rect 442908 251806 442960 251812
rect 442724 251252 442776 251258
rect 442724 251194 442776 251200
rect 442736 250345 442764 251194
rect 442722 250336 442778 250345
rect 442722 250271 442778 250280
rect 441802 247072 441858 247081
rect 441802 247007 441858 247016
rect 441712 239488 441764 239494
rect 441712 239430 441764 239436
rect 441620 239420 441672 239426
rect 441620 239362 441672 239368
rect 441816 238754 441844 247007
rect 442908 246356 442960 246362
rect 442908 246298 442960 246304
rect 442920 246265 442948 246298
rect 442906 246256 442962 246265
rect 442906 246191 442962 246200
rect 442170 244080 442226 244089
rect 442170 244015 442226 244024
rect 442184 242962 442212 244015
rect 442172 242956 442224 242962
rect 442172 242898 442224 242904
rect 442908 242208 442960 242214
rect 442906 242176 442908 242185
rect 442960 242176 442962 242185
rect 442906 242111 442962 242120
rect 441632 238726 441844 238754
rect 441632 227050 441660 238726
rect 441620 227044 441672 227050
rect 441620 226986 441672 226992
rect 441620 198076 441672 198082
rect 441620 198018 441672 198024
rect 441632 171134 441660 198018
rect 441632 171106 442120 171134
rect 440332 167680 440384 167686
rect 440332 167622 440384 167628
rect 441896 147824 441948 147830
rect 441896 147766 441948 147772
rect 440252 145846 440634 145874
rect 441908 145860 441936 147766
rect 442092 145874 442120 171106
rect 442724 149048 442776 149054
rect 442724 148990 442776 148996
rect 442736 147830 442764 148990
rect 443012 148238 443040 303826
rect 443104 255105 443132 316678
rect 444380 303748 444432 303754
rect 444380 303690 444432 303696
rect 443182 293040 443238 293049
rect 443182 292975 443238 292984
rect 443090 255096 443146 255105
rect 443090 255031 443146 255040
rect 443104 238814 443132 255031
rect 443092 238808 443144 238814
rect 443092 238750 443144 238756
rect 443196 237017 443224 292975
rect 443276 242956 443328 242962
rect 443276 242898 443328 242904
rect 443182 237008 443238 237017
rect 443182 236943 443184 236952
rect 443236 236943 443238 236952
rect 443184 236914 443236 236920
rect 443196 236883 443224 236914
rect 443288 209774 443316 242898
rect 443736 239420 443788 239426
rect 443736 239362 443788 239368
rect 443748 238746 443776 239362
rect 443736 238740 443788 238746
rect 443736 238682 443788 238688
rect 443104 209746 443316 209774
rect 443104 206990 443132 209746
rect 443092 206984 443144 206990
rect 443092 206926 443144 206932
rect 443104 151814 443132 206926
rect 443644 163532 443696 163538
rect 443644 163474 443696 163480
rect 443104 151786 443224 151814
rect 443000 148232 443052 148238
rect 443000 148174 443052 148180
rect 442724 147824 442776 147830
rect 442724 147766 442776 147772
rect 442092 145846 442566 145874
rect 443196 145860 443224 151786
rect 443656 148034 443684 163474
rect 444392 151814 444420 303690
rect 444484 242214 444512 371826
rect 445024 358828 445076 358834
rect 445024 358770 445076 358776
rect 444564 296948 444616 296954
rect 444564 296890 444616 296896
rect 444472 242208 444524 242214
rect 444472 242150 444524 242156
rect 444484 202162 444512 242150
rect 444576 239698 444604 296890
rect 445036 285734 445064 358770
rect 447152 318850 447180 399758
rect 448532 320890 448560 399758
rect 452028 398138 452056 399758
rect 454604 398750 454632 399758
rect 457272 398818 457300 399758
rect 458192 399758 459186 399786
rect 460952 399758 461762 399786
rect 464264 399758 464338 399786
rect 466196 399758 466270 399786
rect 467852 399758 468846 399786
rect 470612 399758 471422 399786
rect 473372 399758 473998 399786
rect 474740 399832 474792 399838
rect 474740 399774 474792 399780
rect 475890 399832 475942 399838
rect 478478 399786 478506 400044
rect 481054 399786 481082 400044
rect 475890 399774 475942 399780
rect 457260 398812 457312 398818
rect 457260 398754 457312 398760
rect 454592 398744 454644 398750
rect 454592 398686 454644 398692
rect 452016 398132 452068 398138
rect 452016 398074 452068 398080
rect 452844 395344 452896 395350
rect 452844 395286 452896 395292
rect 452660 363656 452712 363662
rect 452660 363598 452712 363604
rect 450544 355360 450596 355366
rect 450544 355302 450596 355308
rect 448520 320884 448572 320890
rect 448520 320826 448572 320832
rect 447140 318844 447192 318850
rect 447140 318786 447192 318792
rect 447152 318102 447180 318786
rect 447140 318096 447192 318102
rect 447140 318038 447192 318044
rect 450556 312594 450584 355302
rect 452568 315308 452620 315314
rect 452568 315250 452620 315256
rect 452580 314702 452608 315250
rect 451280 314696 451332 314702
rect 451280 314638 451332 314644
rect 452568 314696 452620 314702
rect 452568 314638 452620 314644
rect 450544 312588 450596 312594
rect 450544 312530 450596 312536
rect 448612 305652 448664 305658
rect 448612 305594 448664 305600
rect 447140 303952 447192 303958
rect 447140 303894 447192 303900
rect 446404 302524 446456 302530
rect 446404 302466 446456 302472
rect 445024 285728 445076 285734
rect 445024 285670 445076 285676
rect 444656 265124 444708 265130
rect 444656 265066 444708 265072
rect 444564 239692 444616 239698
rect 444564 239634 444616 239640
rect 444668 233918 444696 265066
rect 444656 233912 444708 233918
rect 444656 233854 444708 233860
rect 444472 202156 444524 202162
rect 444472 202098 444524 202104
rect 445852 178696 445904 178702
rect 445852 178638 445904 178644
rect 444564 176724 444616 176730
rect 444564 176666 444616 176672
rect 444576 171134 444604 176666
rect 445864 171134 445892 178638
rect 444576 171106 444696 171134
rect 445864 171106 446352 171134
rect 444392 151786 444512 151814
rect 443644 148028 443696 148034
rect 443644 147970 443696 147976
rect 444484 145860 444512 151786
rect 444668 145874 444696 171106
rect 446036 148028 446088 148034
rect 446036 147970 446088 147976
rect 446048 145874 446076 147970
rect 446324 147370 446352 171106
rect 446416 147626 446444 302466
rect 446496 301028 446548 301034
rect 446496 300970 446548 300976
rect 446508 259350 446536 300970
rect 446496 259344 446548 259350
rect 446496 259286 446548 259292
rect 446496 256760 446548 256766
rect 446496 256702 446548 256708
rect 446508 148578 446536 256702
rect 446586 201512 446642 201521
rect 446586 201447 446642 201456
rect 446600 151814 446628 201447
rect 447152 162178 447180 303894
rect 448520 301504 448572 301510
rect 448520 301446 448572 301452
rect 447784 287088 447836 287094
rect 447784 287030 447836 287036
rect 447140 162172 447192 162178
rect 447140 162114 447192 162120
rect 446600 151786 446812 151814
rect 446496 148572 446548 148578
rect 446496 148514 446548 148520
rect 446404 147620 446456 147626
rect 446404 147562 446456 147568
rect 446324 147342 446720 147370
rect 446692 145874 446720 147342
rect 446784 145994 446812 151786
rect 447796 147014 447824 287030
rect 448532 251870 448560 301446
rect 448624 272134 448652 305594
rect 449900 300892 449952 300898
rect 449900 300834 449952 300840
rect 448612 272128 448664 272134
rect 448612 272070 448664 272076
rect 448624 267734 448652 272070
rect 448796 269136 448848 269142
rect 448796 269078 448848 269084
rect 448624 267706 448744 267734
rect 448612 259344 448664 259350
rect 448612 259286 448664 259292
rect 448624 258126 448652 259286
rect 448612 258120 448664 258126
rect 448612 258062 448664 258068
rect 448520 251864 448572 251870
rect 448520 251806 448572 251812
rect 448624 151814 448652 258062
rect 448716 227730 448744 267706
rect 448808 235278 448836 269078
rect 448796 235272 448848 235278
rect 448796 235214 448848 235220
rect 449912 234530 449940 300834
rect 449992 289876 450044 289882
rect 449992 289818 450044 289824
rect 450004 236842 450032 289818
rect 450084 281852 450136 281858
rect 450084 281794 450136 281800
rect 449992 236836 450044 236842
rect 449992 236778 450044 236784
rect 449900 234524 449952 234530
rect 449900 234466 449952 234472
rect 448704 227724 448756 227730
rect 448704 227666 448756 227672
rect 448716 226438 448744 227666
rect 448704 226432 448756 226438
rect 448704 226374 448756 226380
rect 449164 226432 449216 226438
rect 449164 226374 449216 226380
rect 449176 166326 449204 226374
rect 449164 166320 449216 166326
rect 449164 166262 449216 166268
rect 449072 159452 449124 159458
rect 449072 159394 449124 159400
rect 448440 151786 448652 151814
rect 447784 147008 447836 147014
rect 447784 146950 447836 146956
rect 446772 145988 446824 145994
rect 446772 145930 446824 145936
rect 448440 145874 448468 151786
rect 448980 147756 449032 147762
rect 448980 147698 449032 147704
rect 444668 145846 445142 145874
rect 446048 145846 446430 145874
rect 446692 145846 447074 145874
rect 448362 145846 448468 145874
rect 448992 145860 449020 147698
rect 400508 145438 401350 145466
rect 403544 145450 403926 145466
rect 417068 145450 417096 145846
rect 423600 145586 423628 145846
rect 423588 145580 423640 145586
rect 423588 145522 423640 145528
rect 403532 145444 403926 145450
rect 400508 144226 400536 145438
rect 403584 145438 403926 145444
rect 417056 145444 417108 145450
rect 403532 145386 403584 145392
rect 417056 145386 417108 145392
rect 400496 144220 400548 144226
rect 400496 144162 400548 144168
rect 449084 143478 449112 159394
rect 449256 156664 449308 156670
rect 449256 156606 449308 156612
rect 449268 151814 449296 156606
rect 449268 151786 449480 151814
rect 449256 145988 449308 145994
rect 449256 145930 449308 145936
rect 449268 145625 449296 145930
rect 449254 145616 449310 145625
rect 449254 145551 449310 145560
rect 449072 143472 449124 143478
rect 449072 143414 449124 143420
rect 449346 143440 449402 143449
rect 449346 143375 449402 143384
rect 400126 140040 400182 140049
rect 400126 139975 400182 139984
rect 449164 130076 449216 130082
rect 449164 130018 449216 130024
rect 449176 122834 449204 130018
rect 449084 122806 449204 122834
rect 399574 111888 399630 111897
rect 399574 111823 399630 111832
rect 399588 111722 399616 111823
rect 399576 111716 399628 111722
rect 399576 111658 399628 111664
rect 399484 93832 399536 93838
rect 399484 93774 399536 93780
rect 398852 84166 399064 84194
rect 398104 46912 398156 46918
rect 398104 46854 398156 46860
rect 398852 35222 398880 84166
rect 399588 46918 399616 111658
rect 399668 97844 399720 97850
rect 399668 97786 399720 97792
rect 399680 96778 399708 97786
rect 399680 96750 400062 96778
rect 400692 95266 400720 96084
rect 400680 95260 400732 95266
rect 400680 95202 400732 95208
rect 401336 88194 401364 96084
rect 402624 88330 402652 96084
rect 403268 93634 403296 96084
rect 403256 93628 403308 93634
rect 403256 93570 403308 93576
rect 404556 92410 404584 96084
rect 405200 93838 405228 96084
rect 405188 93832 405240 93838
rect 405188 93774 405240 93780
rect 404544 92404 404596 92410
rect 404544 92346 404596 92352
rect 405740 92268 405792 92274
rect 405740 92210 405792 92216
rect 405752 91798 405780 92210
rect 406488 91798 406516 96084
rect 407132 93702 407160 96084
rect 407120 93696 407172 93702
rect 407120 93638 407172 93644
rect 407132 92274 407160 93638
rect 407120 92268 407172 92274
rect 407120 92210 407172 92216
rect 405740 91792 405792 91798
rect 405740 91734 405792 91740
rect 406476 91792 406528 91798
rect 406476 91734 406528 91740
rect 403624 90364 403676 90370
rect 403624 90306 403676 90312
rect 401600 88324 401652 88330
rect 401600 88266 401652 88272
rect 402612 88324 402664 88330
rect 402612 88266 402664 88272
rect 400864 88188 400916 88194
rect 400864 88130 400916 88136
rect 401324 88188 401376 88194
rect 401324 88130 401376 88136
rect 399576 46912 399628 46918
rect 399576 46854 399628 46860
rect 398840 35216 398892 35222
rect 398840 35158 398892 35164
rect 396908 31748 396960 31754
rect 396908 31690 396960 31696
rect 396724 19304 396776 19310
rect 396724 19246 396776 19252
rect 400876 10946 400904 88130
rect 401612 86290 401640 88266
rect 401600 86284 401652 86290
rect 401600 86226 401652 86232
rect 400864 10940 400916 10946
rect 400864 10882 400916 10888
rect 395344 4820 395396 4826
rect 395344 4762 395396 4768
rect 403636 4146 403664 90306
rect 405752 50386 405780 91734
rect 407776 84194 407804 96084
rect 409064 93854 409092 96084
rect 409064 93826 409184 93854
rect 409156 89690 409184 93826
rect 409144 89684 409196 89690
rect 409144 89626 409196 89632
rect 408500 89004 408552 89010
rect 408500 88946 408552 88952
rect 407224 84166 407804 84194
rect 405740 50380 405792 50386
rect 405740 50322 405792 50328
rect 407224 36718 407252 84166
rect 408512 61402 408540 88946
rect 408500 61396 408552 61402
rect 408500 61338 408552 61344
rect 409156 51882 409184 89626
rect 409708 89010 409736 96084
rect 410996 92478 411024 96084
rect 410984 92472 411036 92478
rect 410984 92414 411036 92420
rect 409696 89004 409748 89010
rect 409696 88946 409748 88952
rect 411640 84194 411668 96084
rect 412928 84194 412956 96084
rect 413572 89622 413600 96084
rect 413560 89616 413612 89622
rect 413560 89558 413612 89564
rect 414216 84194 414244 96084
rect 415504 90982 415532 96084
rect 416148 92342 416176 96084
rect 417436 93770 417464 96084
rect 416780 93764 416832 93770
rect 416780 93706 416832 93712
rect 417424 93764 417476 93770
rect 417424 93706 417476 93712
rect 416792 92886 416820 93706
rect 418080 92886 418108 96084
rect 419368 95334 419396 96084
rect 419356 95328 419408 95334
rect 419356 95270 419408 95276
rect 416780 92880 416832 92886
rect 416780 92822 416832 92828
rect 418068 92880 418120 92886
rect 418068 92822 418120 92828
rect 416136 92336 416188 92342
rect 416136 92278 416188 92284
rect 416148 91118 416176 92278
rect 416136 91112 416188 91118
rect 416136 91054 416188 91060
rect 415492 90976 415544 90982
rect 415492 90918 415544 90924
rect 416688 90976 416740 90982
rect 416688 90918 416740 90924
rect 416700 86970 416728 90918
rect 416688 86964 416740 86970
rect 416688 86906 416740 86912
rect 411272 84166 411668 84194
rect 412652 84166 412956 84194
rect 414032 84166 414244 84194
rect 411272 78674 411300 84166
rect 411260 78668 411312 78674
rect 411260 78610 411312 78616
rect 409144 51876 409196 51882
rect 409144 51818 409196 51824
rect 407212 36712 407264 36718
rect 407212 36654 407264 36660
rect 412652 8294 412680 84166
rect 412640 8288 412692 8294
rect 412640 8230 412692 8236
rect 414032 6866 414060 84166
rect 416792 60042 416820 92822
rect 418896 92540 418948 92546
rect 418896 92482 418948 92488
rect 418804 86964 418856 86970
rect 418804 86906 418856 86912
rect 416780 60036 416832 60042
rect 416780 59978 416832 59984
rect 418816 6866 418844 86906
rect 418908 72486 418936 92482
rect 418988 91112 419040 91118
rect 418988 91054 419040 91060
rect 419000 86970 419028 91054
rect 418988 86964 419040 86970
rect 418988 86906 419040 86912
rect 420012 84194 420040 96084
rect 420656 92546 420684 96084
rect 420644 92540 420696 92546
rect 420644 92482 420696 92488
rect 421944 84194 421972 96084
rect 422588 95198 422616 96084
rect 422576 95192 422628 95198
rect 422576 95134 422628 95140
rect 423876 93702 423904 96084
rect 423864 93696 423916 93702
rect 423864 93638 423916 93644
rect 424520 92546 424548 96084
rect 425808 94926 425836 96084
rect 425796 94920 425848 94926
rect 425796 94862 425848 94868
rect 422944 92540 422996 92546
rect 422944 92482 422996 92488
rect 424508 92540 424560 92546
rect 424508 92482 424560 92488
rect 419644 84166 420040 84194
rect 420932 84166 421972 84194
rect 419644 80034 419672 84166
rect 419632 80028 419684 80034
rect 419632 79970 419684 79976
rect 418896 72480 418948 72486
rect 418896 72422 418948 72428
rect 420932 20670 420960 84166
rect 422956 41410 422984 92482
rect 426452 90914 426480 96084
rect 427740 91089 427768 96084
rect 427726 91080 427782 91089
rect 427726 91015 427782 91024
rect 426440 90908 426492 90914
rect 426440 90850 426492 90856
rect 427728 90908 427780 90914
rect 427728 90850 427780 90856
rect 422944 41404 422996 41410
rect 422944 41346 422996 41352
rect 427740 35222 427768 90850
rect 428384 90370 428412 96084
rect 428372 90364 428424 90370
rect 428372 90306 428424 90312
rect 429028 89010 429056 96084
rect 430316 93786 430344 96084
rect 430960 95062 430988 96084
rect 430948 95056 431000 95062
rect 430948 94998 431000 95004
rect 432248 94858 432276 96084
rect 432236 94852 432288 94858
rect 432236 94794 432288 94800
rect 430394 93800 430450 93809
rect 430316 93758 430394 93786
rect 427820 89004 427872 89010
rect 427820 88946 427872 88952
rect 429016 89004 429068 89010
rect 429016 88946 429068 88952
rect 427832 80714 427860 88946
rect 430316 84194 430344 93758
rect 430394 93735 430450 93744
rect 432892 92342 432920 96084
rect 432880 92336 432932 92342
rect 432880 92278 432932 92284
rect 434180 84194 434208 96084
rect 434824 84194 434852 96084
rect 435468 93854 435496 96084
rect 436756 94994 436784 96084
rect 436744 94988 436796 94994
rect 436744 94930 436796 94936
rect 435376 93826 435496 93854
rect 435376 93634 435404 93826
rect 435364 93628 435416 93634
rect 435364 93570 435416 93576
rect 429856 84166 430344 84194
rect 433352 84166 434208 84194
rect 434732 84166 434852 84194
rect 427820 80708 427872 80714
rect 427820 80650 427872 80656
rect 427728 35216 427780 35222
rect 427728 35158 427780 35164
rect 420920 20664 420972 20670
rect 420920 20606 420972 20612
rect 429856 9654 429884 84166
rect 433352 77246 433380 84166
rect 433340 77240 433392 77246
rect 433340 77182 433392 77188
rect 434732 59362 434760 84166
rect 434720 59356 434772 59362
rect 434720 59298 434772 59304
rect 435376 57254 435404 93570
rect 437400 91050 437428 96084
rect 438688 95198 438716 96084
rect 438676 95192 438728 95198
rect 438676 95134 438728 95140
rect 438688 95062 438716 95134
rect 438124 95056 438176 95062
rect 438124 94998 438176 95004
rect 438676 95056 438728 95062
rect 438676 94998 438728 95004
rect 438768 95056 438820 95062
rect 438768 94998 438820 95004
rect 437388 91044 437440 91050
rect 437388 90986 437440 90992
rect 435364 57248 435416 57254
rect 435364 57190 435416 57196
rect 438136 33794 438164 94998
rect 438780 94858 438808 94998
rect 438768 94852 438820 94858
rect 438768 94794 438820 94800
rect 439332 84194 439360 96084
rect 440620 93566 440648 96084
rect 441264 94790 441292 96084
rect 441908 95334 441936 96084
rect 441896 95328 441948 95334
rect 441896 95270 441948 95276
rect 442998 95296 443054 95305
rect 442998 95231 443054 95240
rect 441252 94784 441304 94790
rect 441252 94726 441304 94732
rect 440608 93560 440660 93566
rect 440608 93502 440660 93508
rect 438872 84166 439360 84194
rect 438872 73166 438900 84166
rect 438860 73160 438912 73166
rect 438860 73102 438912 73108
rect 438124 33788 438176 33794
rect 438124 33730 438176 33736
rect 443012 26246 443040 95231
rect 443196 93566 443224 96084
rect 443840 95305 443868 96084
rect 443826 95296 443882 95305
rect 443826 95231 443882 95240
rect 443184 93560 443236 93566
rect 443184 93502 443236 93508
rect 445128 84194 445156 96084
rect 445772 93854 445800 96084
rect 447060 95130 447088 96084
rect 447048 95124 447100 95130
rect 447048 95066 447100 95072
rect 445772 93826 445892 93854
rect 447704 93838 447732 96084
rect 448992 95266 449020 96084
rect 448980 95260 449032 95266
rect 448980 95202 449032 95208
rect 444392 84166 445156 84194
rect 444392 49026 444420 84166
rect 444380 49020 444432 49026
rect 444380 48962 444432 48968
rect 445864 39438 445892 93826
rect 447692 93832 447744 93838
rect 447692 93774 447744 93780
rect 447784 92540 447836 92546
rect 447784 92482 447836 92488
rect 447796 64870 447824 92482
rect 447784 64864 447836 64870
rect 447784 64806 447836 64812
rect 445852 39432 445904 39438
rect 445852 39374 445904 39380
rect 443000 26240 443052 26246
rect 443000 26182 443052 26188
rect 449084 13122 449112 122806
rect 449360 117298 449388 143375
rect 449452 141545 449480 151786
rect 449624 148572 449676 148578
rect 449624 148514 449676 148520
rect 449636 145860 449664 148514
rect 449532 143472 449584 143478
rect 449532 143414 449584 143420
rect 449544 143313 449572 143414
rect 449530 143304 449586 143313
rect 449530 143239 449586 143248
rect 449438 141536 449494 141545
rect 449438 141471 449494 141480
rect 449438 130112 449494 130121
rect 449438 130047 449440 130056
rect 449492 130047 449494 130056
rect 449440 130018 449492 130024
rect 449912 129169 449940 234466
rect 450096 233102 450124 281794
rect 451292 236910 451320 314638
rect 451372 302456 451424 302462
rect 451372 302398 451424 302404
rect 451280 236904 451332 236910
rect 451280 236846 451332 236852
rect 450084 233096 450136 233102
rect 450084 233038 450136 233044
rect 450096 232354 450124 233038
rect 450084 232348 450136 232354
rect 450084 232290 450136 232296
rect 450544 232348 450596 232354
rect 450544 232290 450596 232296
rect 449992 209160 450044 209166
rect 449992 209102 450044 209108
rect 450004 138009 450032 209102
rect 450084 171828 450136 171834
rect 450084 171770 450136 171776
rect 449990 138000 450046 138009
rect 449990 137935 450046 137944
rect 450096 135561 450124 171770
rect 450556 136649 450584 232290
rect 451384 231130 451412 302398
rect 451372 231124 451424 231130
rect 451372 231066 451424 231072
rect 451648 210452 451700 210458
rect 451648 210394 451700 210400
rect 451372 200184 451424 200190
rect 451372 200126 451424 200132
rect 451384 142154 451412 200126
rect 451464 198756 451516 198762
rect 451464 198698 451516 198704
rect 451476 142361 451504 198698
rect 451556 155236 451608 155242
rect 451556 155178 451608 155184
rect 451568 147801 451596 155178
rect 451554 147792 451610 147801
rect 451554 147727 451610 147736
rect 451556 147620 451608 147626
rect 451556 147562 451608 147568
rect 451462 142352 451518 142361
rect 451462 142287 451518 142296
rect 451292 142126 451412 142154
rect 451292 138961 451320 142126
rect 451278 138952 451334 138961
rect 451278 138887 451334 138896
rect 450542 136640 450598 136649
rect 450542 136575 450598 136584
rect 450082 135552 450138 135561
rect 450082 135487 450138 135496
rect 449992 132456 450044 132462
rect 449992 132398 450044 132404
rect 450004 131209 450032 132398
rect 449990 131200 450046 131209
rect 449990 131135 450046 131144
rect 449898 129160 449954 129169
rect 449898 129095 449954 129104
rect 449348 117292 449400 117298
rect 449348 117234 449400 117240
rect 449360 117065 449388 117234
rect 449346 117056 449402 117065
rect 449346 116991 449402 117000
rect 449898 101960 449954 101969
rect 449898 101895 449954 101904
rect 449636 92546 449664 96084
rect 449624 92540 449676 92546
rect 449624 92482 449676 92488
rect 449912 15978 449940 101895
rect 450004 33114 450032 131135
rect 451568 125361 451596 147562
rect 451554 125352 451610 125361
rect 451554 125287 451610 125296
rect 451280 124772 451332 124778
rect 451280 124714 451332 124720
rect 451292 124681 451320 124714
rect 451278 124672 451334 124681
rect 451278 124607 451334 124616
rect 451660 124001 451688 210394
rect 452568 144900 452620 144906
rect 452568 144842 452620 144848
rect 452580 144401 452608 144842
rect 452566 144392 452622 144401
rect 452566 144327 452622 144336
rect 452474 142896 452530 142905
rect 452474 142831 452530 142840
rect 452488 142186 452516 142831
rect 452476 142180 452528 142186
rect 452476 142122 452528 142128
rect 451924 140480 451976 140486
rect 451924 140422 451976 140428
rect 451936 140321 451964 140422
rect 451922 140312 451978 140321
rect 451922 140247 451978 140256
rect 452108 138916 452160 138922
rect 452108 138858 452160 138864
rect 452120 138281 452148 138858
rect 452106 138272 452162 138281
rect 452106 138207 452162 138216
rect 451924 135244 451976 135250
rect 451924 135186 451976 135192
rect 451936 134201 451964 135186
rect 451922 134192 451978 134201
rect 451922 134127 451978 134136
rect 452200 133884 452252 133890
rect 452200 133826 452252 133832
rect 452212 133521 452240 133826
rect 452198 133512 452254 133521
rect 452198 133447 452254 133456
rect 452566 130792 452622 130801
rect 452672 130778 452700 363598
rect 452752 294636 452804 294642
rect 452752 294578 452804 294584
rect 452622 130750 452700 130778
rect 452566 130727 452622 130736
rect 452568 129736 452620 129742
rect 452568 129678 452620 129684
rect 452580 129441 452608 129678
rect 452566 129432 452622 129441
rect 452566 129367 452622 129376
rect 452108 128308 452160 128314
rect 452108 128250 452160 128256
rect 452120 127401 452148 128250
rect 452106 127392 452162 127401
rect 452106 127327 452162 127336
rect 452568 126948 452620 126954
rect 452568 126890 452620 126896
rect 452580 126721 452608 126890
rect 452566 126712 452622 126721
rect 452566 126647 452622 126656
rect 452568 125588 452620 125594
rect 452568 125530 452620 125536
rect 452580 125361 452608 125530
rect 452566 125352 452622 125361
rect 452566 125287 452622 125296
rect 451646 123992 451702 124001
rect 451646 123927 451702 123936
rect 452568 122664 452620 122670
rect 452566 122632 452568 122641
rect 452620 122632 452622 122641
rect 452566 122567 452622 122576
rect 450082 120456 450138 120465
rect 450082 120391 450138 120400
rect 449992 33108 450044 33114
rect 449992 33050 450044 33056
rect 449900 15972 449952 15978
rect 449900 15914 449952 15920
rect 449072 13116 449124 13122
rect 449072 13058 449124 13064
rect 450096 12442 450124 120391
rect 452476 118652 452528 118658
rect 452476 118594 452528 118600
rect 452488 117881 452516 118594
rect 452474 117872 452530 117881
rect 452474 117807 452530 117816
rect 451556 115864 451608 115870
rect 451554 115832 451556 115841
rect 451608 115832 451610 115841
rect 451554 115767 451610 115776
rect 451370 115016 451426 115025
rect 451370 114951 451426 114960
rect 451278 106312 451334 106321
rect 451278 106247 451334 106256
rect 450174 104136 450230 104145
rect 450174 104071 450230 104080
rect 450188 82754 450216 104071
rect 450176 82748 450228 82754
rect 450176 82690 450228 82696
rect 451292 38622 451320 106247
rect 451384 66910 451412 114951
rect 452476 114504 452528 114510
rect 452476 114446 452528 114452
rect 452488 113801 452516 114446
rect 452474 113792 452530 113801
rect 452474 113727 452530 113736
rect 452764 113174 452792 294578
rect 452856 236774 452884 395286
rect 457272 393314 457300 398754
rect 457272 393310 457484 393314
rect 457272 393304 457496 393310
rect 457272 393286 457444 393304
rect 457444 393246 457496 393252
rect 456800 380180 456852 380186
rect 456800 380122 456852 380128
rect 456812 379574 456840 380122
rect 456800 379568 456852 379574
rect 456800 379510 456852 379516
rect 456812 373994 456840 379510
rect 456812 373966 456932 373994
rect 454040 358896 454092 358902
rect 454040 358838 454092 358844
rect 454052 259418 454080 358838
rect 455420 305108 455472 305114
rect 455420 305050 455472 305056
rect 454132 299600 454184 299606
rect 454132 299542 454184 299548
rect 454040 259412 454092 259418
rect 454040 259354 454092 259360
rect 454040 238060 454092 238066
rect 454040 238002 454092 238008
rect 452844 236768 452896 236774
rect 452844 236710 452896 236716
rect 452844 206304 452896 206310
rect 452844 206246 452896 206252
rect 452672 113146 452792 113174
rect 452476 111784 452528 111790
rect 452476 111726 452528 111732
rect 452566 111752 452622 111761
rect 452488 111081 452516 111726
rect 452566 111687 452568 111696
rect 452620 111687 452622 111696
rect 452568 111658 452620 111664
rect 452474 111072 452530 111081
rect 452474 111007 452530 111016
rect 452108 110356 452160 110362
rect 452108 110298 452160 110304
rect 452120 109721 452148 110298
rect 452106 109712 452162 109721
rect 452106 109647 452162 109656
rect 451554 109032 451610 109041
rect 451554 108967 451610 108976
rect 451568 73846 451596 108967
rect 451738 108216 451794 108225
rect 451738 108151 451794 108160
rect 451556 73840 451608 73846
rect 451556 73782 451608 73788
rect 451752 69834 451780 108151
rect 452566 106992 452622 107001
rect 452672 106978 452700 113146
rect 452856 109041 452884 206246
rect 452936 191140 452988 191146
rect 452936 191082 452988 191088
rect 452842 109032 452898 109041
rect 452842 108967 452898 108976
rect 452622 106950 452700 106978
rect 452566 106927 452622 106936
rect 452566 104952 452622 104961
rect 452566 104887 452568 104896
rect 452620 104887 452622 104896
rect 452568 104858 452620 104864
rect 452948 103514 452976 191082
rect 452672 103486 452976 103514
rect 452568 103080 452620 103086
rect 452568 103022 452620 103028
rect 452580 102921 452608 103022
rect 452566 102912 452622 102921
rect 452566 102847 452622 102856
rect 452568 100700 452620 100706
rect 452568 100642 452620 100648
rect 452580 100201 452608 100642
rect 452566 100192 452622 100201
rect 452566 100127 452622 100136
rect 452292 98932 452344 98938
rect 452292 98874 452344 98880
rect 452304 98161 452332 98874
rect 452290 98152 452346 98161
rect 452290 98087 452346 98096
rect 452566 97472 452622 97481
rect 452672 97458 452700 103486
rect 454052 98938 454080 238002
rect 454144 224913 454172 299542
rect 454130 224904 454186 224913
rect 454130 224839 454186 224848
rect 454132 193928 454184 193934
rect 454132 193870 454184 193876
rect 454144 103086 454172 193870
rect 455432 152590 455460 305050
rect 456800 302320 456852 302326
rect 456800 302262 456852 302268
rect 455512 226364 455564 226370
rect 455512 226306 455564 226312
rect 455420 152584 455472 152590
rect 455420 152526 455472 152532
rect 454224 149728 454276 149734
rect 454224 149670 454276 149676
rect 454236 124778 454264 149670
rect 454316 146940 454368 146946
rect 454316 146882 454368 146888
rect 454328 135250 454356 146882
rect 454316 135244 454368 135250
rect 454316 135186 454368 135192
rect 454224 124772 454276 124778
rect 454224 124714 454276 124720
rect 455524 115870 455552 226306
rect 455604 159384 455656 159390
rect 455604 159326 455656 159332
rect 455616 140486 455644 159326
rect 455972 147824 456024 147830
rect 455972 147766 456024 147772
rect 455984 142154 456012 147766
rect 456064 147688 456116 147694
rect 456064 147630 456116 147636
rect 456076 145586 456104 147630
rect 456064 145580 456116 145586
rect 456064 145522 456116 145528
rect 455984 142126 456104 142154
rect 455604 140480 455656 140486
rect 455604 140422 455656 140428
rect 455512 115864 455564 115870
rect 455512 115806 455564 115812
rect 456076 113150 456104 142126
rect 456064 113144 456116 113150
rect 456064 113086 456116 113092
rect 454224 104916 454276 104922
rect 454224 104858 454276 104864
rect 454132 103080 454184 103086
rect 454132 103022 454184 103028
rect 454040 98932 454092 98938
rect 454040 98874 454092 98880
rect 452622 97430 452700 97458
rect 452566 97407 452622 97416
rect 453304 97300 453356 97306
rect 453304 97242 453356 97248
rect 453316 93809 453344 97242
rect 453302 93800 453358 93809
rect 453302 93735 453358 93744
rect 454236 88262 454264 104858
rect 456812 93702 456840 302262
rect 456904 238066 456932 373966
rect 458192 323610 458220 399758
rect 458180 323604 458232 323610
rect 458180 323546 458232 323552
rect 458180 312588 458232 312594
rect 458180 312530 458232 312536
rect 458192 311914 458220 312530
rect 458180 311908 458232 311914
rect 458180 311850 458232 311856
rect 457444 311840 457496 311846
rect 457444 311782 457496 311788
rect 456892 238060 456944 238066
rect 456892 238002 456944 238008
rect 456892 152516 456944 152522
rect 456892 152458 456944 152464
rect 456904 110362 456932 152458
rect 456892 110356 456944 110362
rect 456892 110298 456944 110304
rect 456800 93696 456852 93702
rect 456800 93638 456852 93644
rect 457456 93634 457484 311782
rect 458192 306374 458220 311850
rect 460952 311846 460980 399758
rect 464264 398682 464292 399758
rect 464252 398676 464304 398682
rect 464252 398618 464304 398624
rect 466196 397526 466224 399758
rect 464344 397520 464396 397526
rect 464344 397462 464396 397468
rect 466184 397520 466236 397526
rect 466184 397462 466236 397468
rect 460940 311840 460992 311846
rect 460940 311782 460992 311788
rect 458364 308440 458416 308446
rect 458364 308382 458416 308388
rect 458376 307834 458404 308382
rect 458364 307828 458416 307834
rect 458364 307770 458416 307776
rect 458192 306346 458312 306374
rect 458180 303816 458232 303822
rect 458180 303758 458232 303764
rect 458192 93770 458220 303758
rect 458284 238678 458312 306346
rect 458272 238672 458324 238678
rect 458272 238614 458324 238620
rect 458376 237386 458404 307770
rect 463700 305040 463752 305046
rect 463700 304982 463752 304988
rect 459652 302592 459704 302598
rect 459652 302534 459704 302540
rect 458364 237380 458416 237386
rect 458364 237322 458416 237328
rect 458272 229900 458324 229906
rect 458272 229842 458324 229848
rect 458284 128314 458312 229842
rect 458376 138922 458404 237322
rect 458824 203584 458876 203590
rect 458824 203526 458876 203532
rect 458836 152522 458864 203526
rect 459560 189100 459612 189106
rect 459560 189042 459612 189048
rect 458824 152516 458876 152522
rect 458824 152458 458876 152464
rect 458364 138916 458416 138922
rect 458364 138858 458416 138864
rect 458272 128308 458324 128314
rect 458272 128250 458324 128256
rect 458836 94926 458864 152458
rect 459572 149161 459600 189042
rect 459558 149152 459614 149161
rect 459558 149087 459614 149096
rect 459560 147008 459612 147014
rect 459560 146950 459612 146956
rect 459572 122670 459600 146950
rect 459560 122664 459612 122670
rect 459560 122606 459612 122612
rect 459664 95062 459692 302534
rect 463608 273964 463660 273970
rect 463608 273906 463660 273912
rect 463620 273290 463648 273906
rect 462320 273284 462372 273290
rect 462320 273226 462372 273232
rect 463608 273284 463660 273290
rect 463608 273226 463660 273232
rect 460204 266416 460256 266422
rect 460204 266358 460256 266364
rect 459744 236972 459796 236978
rect 459744 236914 459796 236920
rect 459652 95056 459704 95062
rect 459652 94998 459704 95004
rect 458824 94920 458876 94926
rect 458824 94862 458876 94868
rect 458180 93764 458232 93770
rect 458180 93706 458232 93712
rect 457444 93628 457496 93634
rect 457444 93570 457496 93576
rect 459756 93566 459784 236914
rect 460216 189786 460244 266358
rect 460940 251252 460992 251258
rect 460940 251194 460992 251200
rect 460204 189780 460256 189786
rect 460204 189722 460256 189728
rect 460216 189106 460244 189722
rect 460204 189100 460256 189106
rect 460204 189042 460256 189048
rect 460204 146396 460256 146402
rect 460204 146338 460256 146344
rect 459744 93560 459796 93566
rect 459744 93502 459796 93508
rect 454224 88256 454276 88262
rect 454224 88198 454276 88204
rect 451740 69828 451792 69834
rect 451740 69770 451792 69776
rect 451372 66904 451424 66910
rect 451372 66846 451424 66852
rect 460216 60722 460244 146338
rect 460952 95334 460980 251194
rect 461032 221468 461084 221474
rect 461032 221410 461084 221416
rect 460940 95328 460992 95334
rect 460940 95270 460992 95276
rect 461044 92342 461072 221410
rect 462332 92410 462360 273226
rect 462412 251864 462464 251870
rect 462412 251806 462464 251812
rect 462320 92404 462372 92410
rect 462320 92346 462372 92352
rect 461032 92336 461084 92342
rect 461032 92278 461084 92284
rect 462424 90982 462452 251806
rect 463712 94994 463740 304982
rect 464356 204950 464384 397462
rect 466460 318844 466512 318850
rect 466460 318786 466512 318792
rect 465080 308508 465132 308514
rect 465080 308450 465132 308456
rect 464344 204944 464396 204950
rect 464344 204886 464396 204892
rect 464344 178084 464396 178090
rect 464344 178026 464396 178032
rect 464356 125594 464384 178026
rect 465092 129742 465120 308450
rect 465080 129736 465132 129742
rect 465080 129678 465132 129684
rect 464344 125588 464396 125594
rect 464344 125530 464396 125536
rect 466472 111722 466500 318786
rect 467104 262268 467156 262274
rect 467104 262210 467156 262216
rect 467116 245614 467144 262210
rect 467104 245608 467156 245614
rect 467104 245550 467156 245556
rect 467116 228410 467144 245550
rect 467104 228404 467156 228410
rect 467104 228346 467156 228352
rect 467104 206304 467156 206310
rect 467104 206246 467156 206252
rect 466552 148368 466604 148374
rect 466552 148310 466604 148316
rect 466564 147762 466592 148310
rect 466552 147756 466604 147762
rect 466552 147698 466604 147704
rect 466460 111716 466512 111722
rect 466460 111658 466512 111664
rect 463700 94988 463752 94994
rect 463700 94930 463752 94936
rect 462412 90976 462464 90982
rect 462412 90918 462464 90924
rect 466564 84182 466592 147698
rect 467116 144906 467144 206246
rect 467104 144900 467156 144906
rect 467104 144842 467156 144848
rect 467852 97306 467880 399758
rect 469220 306400 469272 306406
rect 469220 306342 469272 306348
rect 467932 277432 467984 277438
rect 467932 277374 467984 277380
rect 467944 235958 467972 277374
rect 467932 235952 467984 235958
rect 467932 235894 467984 235900
rect 467840 97300 467892 97306
rect 467840 97242 467892 97248
rect 467944 89622 467972 235894
rect 469232 111790 469260 306342
rect 470612 188358 470640 399758
rect 472624 393984 472676 393990
rect 472624 393926 472676 393932
rect 471980 303680 472032 303686
rect 471980 303622 472032 303628
rect 470692 302388 470744 302394
rect 470692 302330 470744 302336
rect 470600 188352 470652 188358
rect 470600 188294 470652 188300
rect 469220 111784 469272 111790
rect 469220 111726 469272 111732
rect 470704 90914 470732 302330
rect 470692 90908 470744 90914
rect 470692 90850 470744 90856
rect 467932 89616 467984 89622
rect 467932 89558 467984 89564
rect 466552 84176 466604 84182
rect 466552 84118 466604 84124
rect 471992 73166 472020 303622
rect 472636 132462 472664 393926
rect 473372 373318 473400 399758
rect 473360 373312 473412 373318
rect 473360 373254 473412 373260
rect 474752 226234 474780 399774
rect 477512 399758 478506 399786
rect 480272 399758 481082 399786
rect 482986 399786 483014 400044
rect 485562 399786 485590 400044
rect 488138 399786 488166 400044
rect 490714 399786 490742 400044
rect 482986 399758 483060 399786
rect 477512 366382 477540 399758
rect 477500 366376 477552 366382
rect 477500 366318 477552 366324
rect 477960 334688 478012 334694
rect 477960 334630 478012 334636
rect 477972 334014 478000 334630
rect 477500 334008 477552 334014
rect 477500 333950 477552 333956
rect 477960 334008 478012 334014
rect 477960 333950 478012 333956
rect 476212 299532 476264 299538
rect 476212 299474 476264 299480
rect 476120 280832 476172 280838
rect 476120 280774 476172 280780
rect 476132 280226 476160 280774
rect 476120 280220 476172 280226
rect 476120 280162 476172 280168
rect 476132 240786 476160 280162
rect 476120 240780 476172 240786
rect 476120 240722 476172 240728
rect 474740 226228 474792 226234
rect 474740 226170 474792 226176
rect 472624 132456 472676 132462
rect 472624 132398 472676 132404
rect 476132 93838 476160 240722
rect 476224 206990 476252 299474
rect 476212 206984 476264 206990
rect 476212 206926 476264 206932
rect 476224 206310 476252 206926
rect 476212 206304 476264 206310
rect 476212 206246 476264 206252
rect 476212 166320 476264 166326
rect 476212 166262 476264 166268
rect 476224 165646 476252 166262
rect 476212 165640 476264 165646
rect 476212 165582 476264 165588
rect 476224 126954 476252 165582
rect 476212 126948 476264 126954
rect 476212 126890 476264 126896
rect 477512 100706 477540 333950
rect 480272 184210 480300 399758
rect 482284 388476 482336 388482
rect 482284 388418 482336 388424
rect 480352 285728 480404 285734
rect 480352 285670 480404 285676
rect 480260 184204 480312 184210
rect 480260 184146 480312 184152
rect 477500 100700 477552 100706
rect 477500 100642 477552 100648
rect 480364 95266 480392 285670
rect 482296 133890 482324 388418
rect 483032 319462 483060 399758
rect 485516 399758 485590 399786
rect 487172 399758 488166 399786
rect 489932 399758 490742 399786
rect 492646 399786 492674 400044
rect 495222 399838 495250 400044
rect 494060 399832 494112 399838
rect 492646 399758 492720 399786
rect 494060 399774 494112 399780
rect 495210 399832 495262 399838
rect 497798 399786 497826 400044
rect 499730 399786 499758 400044
rect 495210 399774 495262 399780
rect 485516 398614 485544 399758
rect 485504 398608 485556 398614
rect 485504 398550 485556 398556
rect 483020 319456 483072 319462
rect 483020 319398 483072 319404
rect 484400 300960 484452 300966
rect 484400 300902 484452 300908
rect 482284 133884 482336 133890
rect 482284 133826 482336 133832
rect 484412 118658 484440 300902
rect 485780 233912 485832 233918
rect 485780 233854 485832 233860
rect 485792 233345 485820 233854
rect 485778 233336 485834 233345
rect 485778 233271 485834 233280
rect 484400 118652 484452 118658
rect 484400 118594 484452 118600
rect 485792 114510 485820 233271
rect 487172 181490 487200 399758
rect 489184 396772 489236 396778
rect 489184 396714 489236 396720
rect 489196 229838 489224 396714
rect 489932 359514 489960 399758
rect 492692 393990 492720 399758
rect 492680 393984 492732 393990
rect 492680 393926 492732 393932
rect 489920 359508 489972 359514
rect 489920 359450 489972 359456
rect 489184 229832 489236 229838
rect 489184 229774 489236 229780
rect 487160 181484 487212 181490
rect 487160 181426 487212 181432
rect 485780 114504 485832 114510
rect 485780 114446 485832 114452
rect 480352 95260 480404 95266
rect 480352 95202 480404 95208
rect 476120 93832 476172 93838
rect 476120 93774 476172 93780
rect 494072 88194 494100 399774
rect 497752 399758 497826 399786
rect 499592 399758 499758 399786
rect 502306 399786 502334 400044
rect 504882 399838 504910 400044
rect 503720 399832 503772 399838
rect 502306 399758 502380 399786
rect 503720 399774 503772 399780
rect 504870 399832 504922 399838
rect 507458 399786 507486 400044
rect 509390 399786 509418 400044
rect 504870 399774 504922 399780
rect 497752 398546 497780 399758
rect 497740 398540 497792 398546
rect 497740 398482 497792 398488
rect 498842 396672 498898 396681
rect 498842 396607 498898 396616
rect 496084 393984 496136 393990
rect 496084 393926 496136 393932
rect 496096 280838 496124 393926
rect 496084 280832 496136 280838
rect 496084 280774 496136 280780
rect 498856 171086 498884 396607
rect 499592 377466 499620 399758
rect 502352 397526 502380 399758
rect 502984 398132 503036 398138
rect 502984 398074 503036 398080
rect 500224 397520 500276 397526
rect 500224 397462 500276 397468
rect 502340 397520 502392 397526
rect 502340 397462 502392 397468
rect 499580 377460 499632 377466
rect 499580 377402 499632 377408
rect 498844 171080 498896 171086
rect 498844 171022 498896 171028
rect 498844 142180 498896 142186
rect 498844 142122 498896 142128
rect 494060 88188 494112 88194
rect 494060 88130 494112 88136
rect 471980 73160 472032 73166
rect 471980 73102 472032 73108
rect 460204 60716 460256 60722
rect 460204 60658 460256 60664
rect 451280 38616 451332 38622
rect 451280 38558 451332 38564
rect 464620 35216 464672 35222
rect 464620 35158 464672 35164
rect 464632 33114 464660 35158
rect 464620 33108 464672 33114
rect 464620 33050 464672 33056
rect 498856 20670 498884 142122
rect 500236 89690 500264 397462
rect 502996 342242 503024 398074
rect 502984 342236 503036 342242
rect 502984 342178 503036 342184
rect 503732 117298 503760 399774
rect 506492 399758 507486 399786
rect 509252 399758 509418 399786
rect 511966 399786 511994 400044
rect 514542 399838 514570 400044
rect 513380 399832 513432 399838
rect 511966 399758 512040 399786
rect 513380 399774 513432 399780
rect 514530 399832 514582 399838
rect 516474 399786 516502 400044
rect 519050 399786 519078 400044
rect 514530 399774 514582 399780
rect 506492 185638 506520 399758
rect 508502 395448 508558 395457
rect 508502 395383 508558 395392
rect 508516 371210 508544 395383
rect 508504 371204 508556 371210
rect 508504 371146 508556 371152
rect 509252 322250 509280 399758
rect 512012 398750 512040 399758
rect 512000 398744 512052 398750
rect 512000 398686 512052 398692
rect 512012 397526 512040 398686
rect 512000 397520 512052 397526
rect 512000 397462 512052 397468
rect 512644 397520 512696 397526
rect 512644 397462 512696 397468
rect 512656 334626 512684 397462
rect 512644 334620 512696 334626
rect 512644 334562 512696 334568
rect 513392 333266 513420 399774
rect 516152 399758 516502 399786
rect 518912 399758 519078 399786
rect 521626 399786 521654 400044
rect 524202 399838 524230 400044
rect 523040 399832 523092 399838
rect 521626 399758 521700 399786
rect 523040 399774 523092 399780
rect 524190 399832 524242 399838
rect 526134 399786 526162 400044
rect 528710 399786 528738 400044
rect 524190 399774 524242 399780
rect 513380 333260 513432 333266
rect 513380 333202 513432 333208
rect 509240 322244 509292 322250
rect 509240 322186 509292 322192
rect 506480 185632 506532 185638
rect 506480 185574 506532 185580
rect 516152 173194 516180 399758
rect 518912 388482 518940 399758
rect 520924 395412 520976 395418
rect 520924 395354 520976 395360
rect 518900 388476 518952 388482
rect 518900 388418 518952 388424
rect 520936 193866 520964 395354
rect 521672 374678 521700 399758
rect 522304 395344 522356 395350
rect 522304 395286 522356 395292
rect 521660 374672 521712 374678
rect 521660 374614 521712 374620
rect 520924 193860 520976 193866
rect 520924 193802 520976 193808
rect 516140 173188 516192 173194
rect 516140 173130 516192 173136
rect 522316 148374 522344 395286
rect 523052 369170 523080 399774
rect 526088 399758 526162 399786
rect 528572 399758 528738 399786
rect 531286 399786 531314 400044
rect 531286 399758 531360 399786
rect 526088 397526 526116 399758
rect 526444 399492 526496 399498
rect 526444 399434 526496 399440
rect 525064 397520 525116 397526
rect 525064 397462 525116 397468
rect 526076 397520 526128 397526
rect 526076 397462 526128 397468
rect 523040 369164 523092 369170
rect 523040 369106 523092 369112
rect 522304 148368 522356 148374
rect 522304 148310 522356 148316
rect 503720 117292 503772 117298
rect 503720 117234 503772 117240
rect 525076 95198 525104 397462
rect 526456 217326 526484 399434
rect 528572 340202 528600 399758
rect 530584 398268 530636 398274
rect 530584 398210 530636 398216
rect 528560 340196 528612 340202
rect 528560 340138 528612 340144
rect 526444 217320 526496 217326
rect 526444 217262 526496 217268
rect 530596 215966 530624 398210
rect 530676 398200 530728 398206
rect 530676 398142 530728 398148
rect 530688 358057 530716 398142
rect 531332 393990 531360 399758
rect 531320 393984 531372 393990
rect 531320 393926 531372 393932
rect 531964 389224 532016 389230
rect 531964 389166 532016 389172
rect 531976 384334 532004 389166
rect 531964 384328 532016 384334
rect 531964 384270 532016 384276
rect 530674 358048 530730 358057
rect 530674 357983 530730 357992
rect 531976 273970 532004 384270
rect 531964 273964 532016 273970
rect 531964 273906 532016 273912
rect 533356 229770 533384 409550
rect 533434 409527 533490 409536
rect 533988 400648 534040 400654
rect 533988 400590 534040 400596
rect 533434 400072 533490 400081
rect 533434 400007 533490 400016
rect 533448 398886 533476 400007
rect 533436 398880 533488 398886
rect 533436 398822 533488 398828
rect 534000 245614 534028 400590
rect 534092 246362 534120 490447
rect 534184 345710 534212 566607
rect 534276 407561 534304 607854
rect 534368 551041 534396 618870
rect 536932 614168 536984 614174
rect 536932 614110 536984 614116
rect 536840 601860 536892 601866
rect 536840 601802 536892 601808
rect 535458 600400 535514 600409
rect 535458 600335 535514 600344
rect 535472 574161 535500 600335
rect 535552 596420 535604 596426
rect 535552 596362 535604 596368
rect 535458 574152 535514 574161
rect 535458 574087 535514 574096
rect 535460 569220 535512 569226
rect 535460 569162 535512 569168
rect 535472 568721 535500 569162
rect 535458 568712 535514 568721
rect 535458 568647 535514 568656
rect 535458 563952 535514 563961
rect 535458 563887 535460 563896
rect 535512 563887 535514 563896
rect 535460 563858 535512 563864
rect 535458 556472 535514 556481
rect 535458 556407 535514 556416
rect 535472 554826 535500 556407
rect 535380 554798 535500 554826
rect 535380 553602 535408 554798
rect 535460 554736 535512 554742
rect 535460 554678 535512 554684
rect 535472 553761 535500 554678
rect 535458 553752 535514 553761
rect 535458 553687 535514 553696
rect 535380 553574 535500 553602
rect 534354 551032 534410 551041
rect 534354 550967 534410 550976
rect 534354 429992 534410 430001
rect 534354 429927 534410 429936
rect 534262 407552 534318 407561
rect 534262 407487 534318 407496
rect 534276 380186 534304 407487
rect 534368 387122 534396 429927
rect 535472 404954 535500 553574
rect 535564 536081 535592 596362
rect 535734 596320 535790 596329
rect 535734 596255 535790 596264
rect 535748 596174 535776 596255
rect 535748 596146 535960 596174
rect 535828 594924 535880 594930
rect 535828 594866 535880 594872
rect 535644 594584 535696 594590
rect 535642 594552 535644 594561
rect 535696 594552 535698 594561
rect 535642 594487 535698 594496
rect 535642 591832 535698 591841
rect 535642 591767 535698 591776
rect 535656 590714 535684 591767
rect 535644 590708 535696 590714
rect 535644 590650 535696 590656
rect 535840 590458 535868 594866
rect 535656 590430 535868 590458
rect 535656 571441 535684 590430
rect 535932 586514 535960 596146
rect 535748 586486 535960 586514
rect 535748 584361 535776 586486
rect 535734 584352 535790 584361
rect 535734 584287 535790 584296
rect 535734 581632 535790 581641
rect 535734 581567 535790 581576
rect 535748 581058 535776 581567
rect 535736 581052 535788 581058
rect 535736 580994 535788 581000
rect 535736 579216 535788 579222
rect 535736 579158 535788 579164
rect 535748 578921 535776 579158
rect 535734 578912 535790 578921
rect 535734 578847 535790 578856
rect 535736 576904 535788 576910
rect 535734 576872 535736 576881
rect 535788 576872 535790 576881
rect 535734 576807 535790 576816
rect 535642 571432 535698 571441
rect 535642 571367 535698 571376
rect 535642 561232 535698 561241
rect 535642 561167 535698 561176
rect 535550 536072 535606 536081
rect 535550 536007 535606 536016
rect 535552 533452 535604 533458
rect 535552 533394 535604 533400
rect 535564 533361 535592 533394
rect 535550 533352 535606 533361
rect 535550 533287 535606 533296
rect 535552 528624 535604 528630
rect 535550 528592 535552 528601
rect 535604 528592 535606 528601
rect 535550 528527 535606 528536
rect 535550 521112 535606 521121
rect 535550 521047 535606 521056
rect 535564 520334 535592 521047
rect 535552 520328 535604 520334
rect 535552 520270 535604 520276
rect 535552 518900 535604 518906
rect 535552 518842 535604 518848
rect 535564 518401 535592 518842
rect 535550 518392 535606 518401
rect 535550 518327 535606 518336
rect 535550 515672 535606 515681
rect 535550 515607 535606 515616
rect 535564 515098 535592 515607
rect 535552 515092 535604 515098
rect 535552 515034 535604 515040
rect 535550 513632 535606 513641
rect 535550 513567 535606 513576
rect 535564 513398 535592 513567
rect 535552 513392 535604 513398
rect 535552 513334 535604 513340
rect 535550 508192 535606 508201
rect 535550 508127 535606 508136
rect 535564 507890 535592 508127
rect 535552 507884 535604 507890
rect 535552 507826 535604 507832
rect 535552 506456 535604 506462
rect 535552 506398 535604 506404
rect 535564 506161 535592 506398
rect 535550 506152 535606 506161
rect 535550 506087 535606 506096
rect 535550 503432 535606 503441
rect 535550 503367 535606 503376
rect 535564 502382 535592 503367
rect 535552 502376 535604 502382
rect 535552 502318 535604 502324
rect 535550 500712 535606 500721
rect 535550 500647 535606 500656
rect 535564 499594 535592 500647
rect 535552 499588 535604 499594
rect 535552 499530 535604 499536
rect 535550 495952 535606 495961
rect 535550 495887 535606 495896
rect 535564 495514 535592 495887
rect 535552 495508 535604 495514
rect 535552 495450 535604 495456
rect 535550 493232 535606 493241
rect 535550 493167 535606 493176
rect 535564 492726 535592 493167
rect 535552 492720 535604 492726
rect 535552 492662 535604 492668
rect 535550 485752 535606 485761
rect 535550 485687 535606 485696
rect 535564 484430 535592 485687
rect 535552 484424 535604 484430
rect 535552 484366 535604 484372
rect 535552 483064 535604 483070
rect 535550 483032 535552 483041
rect 535604 483032 535606 483041
rect 535550 482967 535606 482976
rect 535552 482928 535604 482934
rect 535552 482870 535604 482876
rect 535380 404926 535500 404954
rect 535380 404274 535408 404926
rect 535458 404832 535514 404841
rect 535458 404767 535514 404776
rect 535472 404394 535500 404767
rect 535460 404388 535512 404394
rect 535460 404330 535512 404336
rect 535380 404246 535500 404274
rect 534356 387116 534408 387122
rect 534356 387058 534408 387064
rect 534264 380180 534316 380186
rect 534264 380122 534316 380128
rect 534172 345704 534224 345710
rect 534172 345646 534224 345652
rect 534080 246356 534132 246362
rect 534080 246298 534132 246304
rect 533988 245608 534040 245614
rect 533988 245550 534040 245556
rect 533344 229764 533396 229770
rect 533344 229706 533396 229712
rect 530584 215960 530636 215966
rect 530584 215902 530636 215908
rect 535472 197266 535500 404246
rect 535460 197260 535512 197266
rect 535460 197202 535512 197208
rect 535564 151774 535592 482870
rect 535656 378826 535684 561167
rect 535826 523832 535882 523841
rect 535826 523767 535882 523776
rect 535840 523734 535868 523767
rect 536852 523734 536880 601802
rect 536944 549001 536972 614110
rect 537024 612740 537076 612746
rect 537024 612682 537076 612688
rect 537036 611454 537064 612682
rect 537024 611448 537076 611454
rect 537024 611390 537076 611396
rect 537036 605834 537064 611390
rect 537036 605806 537156 605834
rect 537024 599072 537076 599078
rect 537024 599014 537076 599020
rect 536930 548992 536986 549001
rect 536930 548927 536986 548936
rect 537036 546281 537064 599014
rect 537128 594590 537156 605806
rect 537116 594584 537168 594590
rect 537116 594526 537168 594532
rect 538232 579222 538260 702578
rect 543476 699718 543504 703520
rect 559668 699718 559696 703520
rect 540244 699712 540296 699718
rect 540244 699654 540296 699660
rect 543464 699712 543516 699718
rect 543464 699654 543516 699660
rect 552664 699712 552716 699718
rect 552664 699654 552716 699660
rect 559656 699712 559708 699718
rect 559656 699654 559708 699660
rect 540256 612746 540284 699654
rect 549904 683188 549956 683194
rect 549904 683130 549956 683136
rect 543004 670744 543056 670750
rect 543004 670686 543056 670692
rect 540244 612740 540296 612746
rect 540244 612682 540296 612688
rect 542452 599140 542504 599146
rect 542452 599082 542504 599088
rect 538312 597780 538364 597786
rect 538312 597722 538364 597728
rect 538220 579216 538272 579222
rect 538220 579158 538272 579164
rect 538220 563916 538272 563922
rect 538220 563858 538272 563864
rect 537022 546272 537078 546281
rect 537022 546207 537078 546216
rect 537022 538792 537078 538801
rect 537022 538727 537078 538736
rect 535828 523728 535880 523734
rect 535828 523670 535880 523676
rect 536840 523728 536892 523734
rect 536840 523670 536892 523676
rect 536746 510912 536802 510921
rect 536802 510870 536880 510898
rect 536746 510847 536802 510856
rect 535734 488472 535790 488481
rect 535734 488407 535790 488416
rect 535748 482934 535776 488407
rect 535736 482928 535788 482934
rect 535736 482870 535788 482876
rect 535734 478272 535790 478281
rect 535734 478207 535790 478216
rect 535748 477562 535776 478207
rect 535736 477556 535788 477562
rect 535736 477498 535788 477504
rect 535734 475552 535790 475561
rect 535734 475487 535790 475496
rect 535748 474774 535776 475487
rect 535736 474768 535788 474774
rect 535736 474710 535788 474716
rect 535734 472832 535790 472841
rect 535734 472767 535790 472776
rect 535748 472258 535776 472767
rect 535736 472252 535788 472258
rect 535736 472194 535788 472200
rect 535734 470792 535790 470801
rect 535734 470727 535790 470736
rect 535748 470626 535776 470727
rect 535736 470620 535788 470626
rect 535736 470562 535788 470568
rect 535734 468072 535790 468081
rect 535734 468007 535736 468016
rect 535788 468007 535790 468016
rect 535736 467978 535788 467984
rect 535734 465352 535790 465361
rect 535734 465287 535790 465296
rect 535748 465118 535776 465287
rect 535736 465112 535788 465118
rect 535736 465054 535788 465060
rect 535734 462632 535790 462641
rect 535734 462567 535790 462576
rect 535748 462398 535776 462567
rect 535736 462392 535788 462398
rect 535736 462334 535788 462340
rect 535734 460592 535790 460601
rect 535734 460527 535790 460536
rect 535748 459610 535776 460527
rect 535736 459604 535788 459610
rect 535736 459546 535788 459552
rect 535734 457872 535790 457881
rect 535734 457807 535790 457816
rect 535748 456822 535776 457807
rect 535736 456816 535788 456822
rect 535736 456758 535788 456764
rect 535734 453112 535790 453121
rect 535734 453047 535790 453056
rect 535748 452674 535776 453047
rect 535736 452668 535788 452674
rect 535736 452610 535788 452616
rect 535734 447672 535790 447681
rect 535734 447607 535790 447616
rect 535748 447166 535776 447607
rect 535736 447160 535788 447166
rect 535736 447102 535788 447108
rect 535734 444952 535790 444961
rect 535734 444887 535790 444896
rect 535748 444446 535776 444887
rect 535736 444440 535788 444446
rect 535736 444382 535788 444388
rect 535734 442912 535790 442921
rect 535734 442847 535790 442856
rect 535748 441658 535776 442847
rect 535736 441652 535788 441658
rect 535736 441594 535788 441600
rect 535734 435432 535790 435441
rect 535734 435367 535790 435376
rect 535748 434790 535776 435367
rect 535736 434784 535788 434790
rect 535736 434726 535788 434732
rect 535734 432712 535790 432721
rect 535734 432647 535790 432656
rect 535644 378820 535696 378826
rect 535644 378762 535696 378768
rect 535748 367810 535776 432647
rect 535826 427272 535882 427281
rect 535826 427207 535882 427216
rect 535840 426494 535868 427207
rect 535828 426488 535880 426494
rect 535828 426430 535880 426436
rect 535826 422512 535882 422521
rect 535826 422447 535882 422456
rect 535840 422346 535868 422447
rect 535828 422340 535880 422346
rect 535828 422282 535880 422288
rect 535826 419792 535882 419801
rect 535826 419727 535882 419736
rect 535840 419558 535868 419727
rect 535828 419552 535880 419558
rect 535828 419494 535880 419500
rect 535826 417752 535882 417761
rect 535826 417687 535882 417696
rect 535840 417382 535868 417687
rect 535828 417376 535880 417382
rect 535828 417318 535880 417324
rect 535826 415032 535882 415041
rect 535826 414967 535882 414976
rect 535840 414050 535868 414967
rect 535828 414044 535880 414050
rect 535828 413986 535880 413992
rect 535826 412312 535882 412321
rect 535826 412247 535882 412256
rect 535840 411330 535868 412247
rect 535828 411324 535880 411330
rect 535828 411266 535880 411272
rect 535826 402112 535882 402121
rect 535826 402047 535882 402056
rect 535840 401674 535868 402047
rect 535828 401668 535880 401674
rect 535828 401610 535880 401616
rect 535736 367804 535788 367810
rect 535736 367746 535788 367752
rect 536852 160750 536880 510870
rect 536930 440192 536986 440201
rect 536930 440127 536986 440136
rect 536944 189854 536972 440127
rect 537036 327729 537064 538727
rect 537116 528624 537168 528630
rect 537116 528566 537168 528572
rect 537022 327720 537078 327729
rect 537022 327655 537078 327664
rect 537128 326398 537156 528566
rect 537116 326392 537168 326398
rect 537116 326334 537168 326340
rect 538232 198014 538260 563858
rect 538324 400654 538352 597722
rect 539692 596488 539744 596494
rect 539692 596430 539744 596436
rect 538864 594992 538916 594998
rect 538864 594934 538916 594940
rect 538402 594824 538458 594833
rect 538402 594759 538458 594768
rect 538416 569226 538444 594759
rect 538404 569220 538456 569226
rect 538404 569162 538456 569168
rect 538876 563718 538904 594934
rect 539600 576904 539652 576910
rect 539600 576846 539652 576852
rect 538864 563712 538916 563718
rect 538864 563654 538916 563660
rect 538404 515092 538456 515098
rect 538404 515034 538456 515040
rect 538312 400648 538364 400654
rect 538312 400590 538364 400596
rect 538416 338774 538444 515034
rect 538496 472252 538548 472258
rect 538496 472194 538548 472200
rect 538508 395962 538536 472194
rect 538496 395956 538548 395962
rect 538496 395898 538548 395904
rect 538404 338768 538456 338774
rect 538404 338710 538456 338716
rect 538220 198008 538272 198014
rect 538220 197950 538272 197956
rect 536932 189848 536984 189854
rect 536932 189790 536984 189796
rect 539612 169046 539640 576846
rect 539704 533458 539732 596430
rect 539692 533452 539744 533458
rect 539692 533394 539744 533400
rect 539692 468036 539744 468042
rect 539692 467978 539744 467984
rect 539704 398138 539732 467978
rect 540980 462392 541032 462398
rect 540980 462334 541032 462340
rect 539784 422340 539836 422346
rect 539784 422282 539836 422288
rect 539692 398132 539744 398138
rect 539692 398074 539744 398080
rect 539796 389842 539824 422282
rect 539876 417376 539928 417382
rect 539876 417318 539928 417324
rect 539888 398274 539916 417318
rect 539876 398268 539928 398274
rect 539876 398210 539928 398216
rect 540992 396030 541020 462334
rect 541072 452668 541124 452674
rect 541072 452610 541124 452616
rect 541084 398206 541112 452610
rect 541164 411324 541216 411330
rect 541164 411266 541216 411272
rect 541072 398200 541124 398206
rect 541072 398142 541124 398148
rect 540980 396024 541032 396030
rect 540980 395966 541032 395972
rect 539784 389836 539836 389842
rect 539784 389778 539836 389784
rect 541176 385014 541204 411266
rect 542360 404388 542412 404394
rect 542360 404330 542412 404336
rect 541256 401668 541308 401674
rect 541256 401610 541308 401616
rect 541268 391950 541296 401610
rect 541256 391944 541308 391950
rect 541256 391886 541308 391892
rect 541164 385008 541216 385014
rect 541164 384950 541216 384956
rect 542372 266354 542400 404330
rect 542464 395418 542492 599082
rect 542544 447160 542596 447166
rect 542544 447102 542596 447108
rect 542452 395412 542504 395418
rect 542452 395354 542504 395360
rect 542556 394670 542584 447102
rect 543016 398818 543044 670686
rect 549916 601798 549944 683130
rect 552676 616146 552704 699654
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 570604 696992 570656 696998
rect 570604 696934 570656 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 552664 616140 552716 616146
rect 552664 616082 552716 616088
rect 562324 607300 562376 607306
rect 562324 607242 562376 607248
rect 549260 601792 549312 601798
rect 549260 601734 549312 601740
rect 549904 601792 549956 601798
rect 549904 601734 549956 601740
rect 544476 600364 544528 600370
rect 544476 600306 544528 600312
rect 543740 597712 543792 597718
rect 543740 597654 543792 597660
rect 543004 398812 543056 398818
rect 543004 398754 543056 398760
rect 542544 394664 542596 394670
rect 542544 394606 542596 394612
rect 543752 328438 543780 597654
rect 544384 595128 544436 595134
rect 544384 595070 544436 595076
rect 543832 474768 543884 474774
rect 543832 474710 543884 474716
rect 543844 381546 543872 474710
rect 543924 456816 543976 456822
rect 543924 456758 543976 456764
rect 543936 399498 543964 456758
rect 543924 399492 543976 399498
rect 543924 399434 543976 399440
rect 543832 381540 543884 381546
rect 543832 381482 543884 381488
rect 544396 365702 544424 595070
rect 544488 525774 544516 600306
rect 547880 597848 547932 597854
rect 545118 597816 545174 597825
rect 547880 597790 547932 597796
rect 545118 597751 545174 597760
rect 544476 525768 544528 525774
rect 544476 525710 544528 525716
rect 545132 395350 545160 597751
rect 546500 502376 546552 502382
rect 546500 502318 546552 502324
rect 545212 470620 545264 470626
rect 545212 470562 545264 470568
rect 545224 397390 545252 470562
rect 545304 465112 545356 465118
rect 545304 465054 545356 465060
rect 545316 397458 545344 465054
rect 545396 419552 545448 419558
rect 545396 419494 545448 419500
rect 545304 397452 545356 397458
rect 545304 397394 545356 397400
rect 545212 397384 545264 397390
rect 545212 397326 545264 397332
rect 545120 395344 545172 395350
rect 545120 395286 545172 395292
rect 545408 386374 545436 419494
rect 546512 398585 546540 502318
rect 546592 495508 546644 495514
rect 546592 495450 546644 495456
rect 546498 398576 546554 398585
rect 546498 398511 546554 398520
rect 546604 396778 546632 495450
rect 546684 434784 546736 434790
rect 546684 434726 546736 434732
rect 546592 396772 546644 396778
rect 546592 396714 546644 396720
rect 545396 386368 545448 386374
rect 545396 386310 545448 386316
rect 546696 383042 546724 434726
rect 546684 383036 546736 383042
rect 546684 382978 546736 382984
rect 544384 365696 544436 365702
rect 544384 365638 544436 365644
rect 547892 350538 547920 597790
rect 549272 518906 549300 601734
rect 552020 597916 552072 597922
rect 552020 597858 552072 597864
rect 549352 520328 549404 520334
rect 549352 520270 549404 520276
rect 549260 518900 549312 518906
rect 549260 518842 549312 518848
rect 548524 513392 548576 513398
rect 548524 513334 548576 513340
rect 547972 499588 548024 499594
rect 547972 499530 548024 499536
rect 547984 398721 548012 499530
rect 548156 441652 548208 441658
rect 548156 441594 548208 441600
rect 548064 426488 548116 426494
rect 548064 426430 548116 426436
rect 547970 398712 548026 398721
rect 547970 398647 548026 398656
rect 548076 351898 548104 426430
rect 548168 376038 548196 441594
rect 548536 431254 548564 513334
rect 549260 477556 549312 477562
rect 549260 477498 549312 477504
rect 548524 431248 548576 431254
rect 548524 431190 548576 431196
rect 548156 376032 548208 376038
rect 548156 375974 548208 375980
rect 548064 351892 548116 351898
rect 548064 351834 548116 351840
rect 547880 350532 547932 350538
rect 547880 350474 547932 350480
rect 543740 328432 543792 328438
rect 543740 328374 543792 328380
rect 542360 266348 542412 266354
rect 542360 266290 542412 266296
rect 539600 169040 539652 169046
rect 539600 168982 539652 168988
rect 536840 160744 536892 160750
rect 536840 160686 536892 160692
rect 535552 151768 535604 151774
rect 535552 151710 535604 151716
rect 525064 95192 525116 95198
rect 525064 95134 525116 95140
rect 500224 89684 500276 89690
rect 500224 89626 500276 89632
rect 549272 88330 549300 477498
rect 549364 382226 549392 520270
rect 550640 507884 550692 507890
rect 550640 507826 550692 507832
rect 549444 484424 549496 484430
rect 549444 484366 549496 484372
rect 549456 395894 549484 484366
rect 550652 399809 550680 507826
rect 550732 492720 550784 492726
rect 550732 492662 550784 492668
rect 550744 399945 550772 492662
rect 550824 444440 550876 444446
rect 550824 444382 550876 444388
rect 550730 399936 550786 399945
rect 550730 399871 550786 399880
rect 550638 399800 550694 399809
rect 550638 399735 550694 399744
rect 549444 395888 549496 395894
rect 549444 395830 549496 395836
rect 550836 394466 550864 444382
rect 550824 394460 550876 394466
rect 550824 394402 550876 394408
rect 549352 382220 549404 382226
rect 549352 382162 549404 382168
rect 552032 334694 552060 597858
rect 561680 597576 561732 597582
rect 561680 597518 561732 597524
rect 553492 595060 553544 595066
rect 553492 595002 553544 595008
rect 553400 483064 553452 483070
rect 553400 483006 553452 483012
rect 552112 459604 552164 459610
rect 552112 459546 552164 459552
rect 552124 397322 552152 459546
rect 552112 397316 552164 397322
rect 552112 397258 552164 397264
rect 552020 334688 552072 334694
rect 552020 334630 552072 334636
rect 553412 175982 553440 483006
rect 553504 299470 553532 595002
rect 554044 590708 554096 590714
rect 554044 590650 554096 590656
rect 554056 406434 554084 590650
rect 560944 576904 560996 576910
rect 560944 576846 560996 576852
rect 558184 523728 558236 523734
rect 558184 523670 558236 523676
rect 556804 456816 556856 456822
rect 556804 456758 556856 456764
rect 554044 406428 554096 406434
rect 554044 406370 554096 406376
rect 556816 315314 556844 456758
rect 558196 419490 558224 523670
rect 558184 419484 558236 419490
rect 558184 419426 558236 419432
rect 560956 398750 560984 576846
rect 560944 398744 560996 398750
rect 560944 398686 560996 398692
rect 556804 315308 556856 315314
rect 556804 315250 556856 315256
rect 553492 299464 553544 299470
rect 553492 299406 553544 299412
rect 561692 236706 561720 597518
rect 562336 591326 562364 607242
rect 570616 595678 570644 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 574744 597644 574796 597650
rect 574744 597586 574796 597592
rect 569960 595672 570012 595678
rect 569960 595614 570012 595620
rect 570604 595672 570656 595678
rect 570604 595614 570656 595620
rect 569972 594862 570000 595614
rect 569960 594856 570012 594862
rect 569960 594798 570012 594804
rect 562324 591320 562376 591326
rect 562324 591262 562376 591268
rect 562336 554742 562364 591262
rect 563704 581052 563756 581058
rect 563704 580994 563756 581000
rect 562324 554736 562376 554742
rect 562324 554678 562376 554684
rect 563716 511290 563744 580994
rect 563704 511284 563756 511290
rect 563704 511226 563756 511232
rect 569972 506462 570000 594798
rect 574756 538218 574784 597586
rect 582380 596284 582432 596290
rect 582380 596226 582432 596232
rect 579804 591320 579856 591326
rect 579804 591262 579856 591268
rect 579816 591025 579844 591262
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 575480 563712 575532 563718
rect 575480 563654 575532 563660
rect 575492 563106 575520 563654
rect 579816 563106 579844 564295
rect 575480 563100 575532 563106
rect 575480 563042 575532 563048
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 574744 538212 574796 538218
rect 574744 538154 574796 538160
rect 569960 506456 570012 506462
rect 569960 506398 570012 506404
rect 571248 431248 571300 431254
rect 571248 431190 571300 431196
rect 571260 429894 571288 431190
rect 570604 429888 570656 429894
rect 570604 429830 570656 429836
rect 571248 429888 571300 429894
rect 571248 429830 571300 429836
rect 563060 414044 563112 414050
rect 563060 413986 563112 413992
rect 563072 384334 563100 413986
rect 563060 384328 563112 384334
rect 563060 384270 563112 384276
rect 563072 379506 563100 384270
rect 563060 379500 563112 379506
rect 563060 379442 563112 379448
rect 570616 261526 570644 429830
rect 574744 405000 574796 405006
rect 574744 404942 574796 404948
rect 574756 348430 574784 404942
rect 574744 348424 574796 348430
rect 574744 348366 574796 348372
rect 575492 308446 575520 563042
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 579804 525768 579856 525774
rect 579804 525710 579856 525716
rect 579816 524521 579844 525710
rect 579802 524512 579858 524521
rect 579802 524447 579858 524456
rect 579618 511320 579674 511329
rect 579618 511255 579620 511264
rect 579672 511255 579674 511264
rect 579620 511226 579672 511232
rect 576860 406428 576912 406434
rect 576860 406370 576912 406376
rect 576872 405006 576900 406370
rect 576860 405000 576912 405006
rect 576860 404942 576912 404948
rect 579632 392630 579660 511226
rect 580262 484664 580318 484673
rect 580262 484599 580318 484608
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 429894 580212 431559
rect 580172 429888 580224 429894
rect 580172 429830 580224 429836
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 579712 405000 579764 405006
rect 579710 404968 579712 404977
rect 579764 404968 579766 404977
rect 579710 404903 579766 404912
rect 580276 394534 580304 484599
rect 582392 458153 582420 596226
rect 582470 471472 582526 471481
rect 582470 471407 582526 471416
rect 580906 458144 580962 458153
rect 580906 458079 580962 458088
rect 582378 458144 582434 458153
rect 582378 458079 582434 458088
rect 580920 456822 580948 458079
rect 580908 456816 580960 456822
rect 580908 456758 580960 456764
rect 582484 394602 582512 471407
rect 582472 394596 582524 394602
rect 582472 394538 582524 394544
rect 580264 394528 580316 394534
rect 580264 394470 580316 394476
rect 579620 392624 579672 392630
rect 579620 392566 579672 392572
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 575480 308440 575532 308446
rect 575480 308382 575532 308388
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580276 239426 580304 325207
rect 582378 272232 582434 272241
rect 582378 272167 582434 272176
rect 580264 239420 580316 239426
rect 580264 239362 580316 239368
rect 561680 236700 561732 236706
rect 561680 236642 561732 236648
rect 582392 233918 582420 272167
rect 582380 233912 582432 233918
rect 582380 233854 582432 233860
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 579620 224256 579672 224262
rect 579620 224198 579672 224204
rect 553400 175976 553452 175982
rect 553400 175918 553452 175924
rect 576124 99408 576176 99414
rect 576124 99350 576176 99356
rect 576136 92274 576164 99350
rect 576124 92268 576176 92274
rect 576124 92210 576176 92216
rect 549260 88324 549312 88330
rect 549260 88266 549312 88272
rect 498844 20664 498896 20670
rect 498844 20606 498896 20612
rect 450084 12436 450136 12442
rect 450084 12378 450136 12384
rect 429844 9648 429896 9654
rect 429844 9590 429896 9596
rect 414020 6860 414072 6866
rect 414020 6802 414072 6808
rect 418804 6860 418856 6866
rect 418804 6802 418856 6808
rect 403624 4140 403676 4146
rect 403624 4082 403676 4088
rect 355324 3460 355376 3466
rect 355324 3402 355376 3408
rect 348026 326 348464 354
rect 348026 -960 348138 326
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579632 354 579660 224198
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 579988 206984 580040 206990
rect 579988 206926 580040 206932
rect 580000 205737 580028 206926
rect 579986 205728 580042 205737
rect 579986 205663 580042 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580184 152522 580212 152623
rect 580172 152516 580224 152522
rect 580172 152458 580224 152464
rect 580356 146328 580408 146334
rect 580356 146270 580408 146276
rect 580264 145580 580316 145586
rect 580264 145522 580316 145528
rect 580276 126041 580304 145522
rect 580368 139369 580396 146270
rect 580354 139360 580410 139369
rect 580354 139295 580410 139304
rect 580262 126032 580318 126041
rect 580262 125967 580318 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579894 33144 579950 33153
rect 579894 33079 579896 33088
rect 579948 33079 579950 33088
rect 579896 33050 579948 33056
rect 579896 20664 579948 20670
rect 579896 20606 579948 20612
rect 579908 19825 579936 20606
rect 579894 19816 579950 19825
rect 579894 19751 579950 19760
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 579774 354 579886 480
rect 579632 326 579886 354
rect 579774 -960 579886 326
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3146 553832 3202 553888
rect 3422 527856 3478 527912
rect 3422 514800 3478 514856
rect 3054 501744 3110 501800
rect 3882 475632 3938 475688
rect 3422 462612 3424 462632
rect 3424 462612 3476 462632
rect 3476 462612 3478 462632
rect 3422 462576 3478 462612
rect 3422 449556 3424 449576
rect 3424 449556 3476 449576
rect 3476 449556 3478 449576
rect 3422 449520 3478 449556
rect 4066 423544 4122 423600
rect 3146 410488 3202 410544
rect 3974 397432 4030 397488
rect 2962 371320 3018 371376
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 3330 345344 3386 345400
rect 3146 319232 3202 319288
rect 3238 306176 3294 306232
rect 3238 293120 3294 293176
rect 3514 267144 3570 267200
rect 3422 254088 3478 254144
rect 3330 241032 3386 241088
rect 3514 214920 3570 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 2778 84632 2834 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 16578 72392 16634 72448
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3514 32408 3570 32464
rect 3514 19352 3570 19408
rect 8298 24112 8354 24168
rect 3514 6432 3570 6488
rect 9678 10240 9734 10296
rect 17958 29552 18014 29608
rect 16302 2624 16358 2680
rect 38566 252456 38622 252512
rect 31758 68176 31814 68232
rect 42706 587968 42762 588024
rect 44822 586608 44878 586664
rect 43994 585248 44050 585304
rect 43902 197240 43958 197296
rect 53470 217232 53526 217288
rect 54850 275848 54906 275904
rect 54758 238312 54814 238368
rect 56506 583888 56562 583944
rect 58990 584024 59046 584080
rect 56414 195200 56470 195256
rect 56506 192480 56562 192536
rect 50986 186904 51042 186960
rect 57702 251096 57758 251152
rect 58622 391992 58678 392048
rect 59082 393216 59138 393272
rect 59082 391992 59138 392048
rect 60462 511808 60518 511864
rect 61382 585112 61438 585168
rect 60646 579128 60702 579184
rect 60738 572328 60794 572384
rect 60738 568928 60794 568984
rect 60738 565528 60794 565584
rect 60738 555328 60794 555384
rect 60738 552608 60794 552664
rect 60738 549208 60794 549264
rect 60738 545828 60794 545864
rect 60738 545808 60740 545828
rect 60740 545808 60792 545828
rect 60792 545808 60794 545828
rect 60738 542428 60794 542464
rect 60738 542408 60740 542428
rect 60740 542408 60792 542428
rect 60792 542408 60794 542428
rect 60738 539008 60794 539064
rect 60738 532208 60794 532264
rect 60738 528808 60794 528864
rect 60738 525408 60794 525464
rect 60738 492088 60794 492144
rect 60738 488688 60794 488744
rect 60738 485288 60794 485344
rect 60738 481888 60794 481944
rect 60738 478488 60794 478544
rect 60738 468288 60794 468344
rect 60738 464888 60794 464944
rect 60738 458088 60794 458144
rect 60738 451968 60794 452024
rect 60738 445168 60794 445224
rect 60738 441768 60794 441824
rect 60738 431568 60794 431624
rect 60738 428168 60794 428224
rect 60738 424768 60794 424824
rect 60738 421368 60794 421424
rect 61014 417968 61070 418024
rect 60830 414568 60886 414624
rect 61566 575728 61622 575784
rect 61566 535608 61622 535664
rect 61474 508408 61530 508464
rect 62302 505008 62358 505064
rect 63130 505008 63186 505064
rect 62026 502288 62082 502344
rect 61934 498888 61990 498944
rect 61842 448568 61898 448624
rect 60738 407788 60794 407824
rect 60738 407768 60740 407788
rect 60740 407768 60792 407788
rect 60792 407768 60794 407788
rect 60646 238448 60702 238504
rect 62762 495488 62818 495544
rect 63130 461488 63186 461544
rect 63222 436736 63278 436792
rect 74354 585248 74410 585304
rect 80702 586608 80758 586664
rect 118698 593408 118754 593464
rect 119342 593408 119398 593464
rect 115570 586744 115626 586800
rect 134246 585112 134302 585168
rect 156786 587968 156842 588024
rect 178590 592184 178646 592240
rect 175462 585112 175518 585168
rect 188250 592048 188306 592104
rect 210422 586336 210478 586392
rect 210882 586336 210938 586392
rect 220542 586608 220598 586664
rect 220726 586608 220782 586664
rect 64786 584568 64842 584624
rect 63498 579128 63554 579184
rect 63406 471708 63462 471744
rect 63406 471688 63408 471708
rect 63408 471688 63460 471708
rect 63460 471688 63462 471708
rect 63406 434968 63462 435024
rect 63314 414568 63370 414624
rect 63222 411304 63278 411360
rect 63498 417968 63554 418024
rect 64878 404368 64934 404424
rect 62854 238176 62910 238232
rect 65982 297336 66038 297392
rect 65798 233824 65854 233880
rect 68282 291760 68338 291816
rect 67730 291080 67786 291136
rect 67638 290400 67694 290456
rect 67730 289720 67786 289776
rect 67638 289040 67694 289096
rect 67638 287680 67694 287736
rect 67730 287000 67786 287056
rect 68006 284824 68062 284880
rect 67638 284316 67640 284336
rect 67640 284316 67692 284336
rect 67692 284316 67694 284336
rect 67638 284280 67694 284316
rect 68006 283600 68062 283656
rect 67730 282920 67786 282976
rect 68926 290808 68982 290864
rect 68926 286320 68982 286376
rect 68742 285640 68798 285696
rect 68650 284960 68706 285016
rect 68926 283600 68982 283656
rect 68558 281560 68614 281616
rect 67638 280880 67694 280936
rect 67638 280220 67694 280256
rect 67638 280200 67640 280220
rect 67640 280200 67692 280220
rect 67692 280200 67694 280220
rect 67638 279520 67694 279576
rect 67362 278840 67418 278896
rect 67638 278160 67694 278216
rect 67638 277480 67694 277536
rect 67730 276800 67786 276856
rect 67638 276120 67694 276176
rect 67638 275440 67694 275496
rect 68282 274760 68338 274816
rect 67638 274080 67694 274136
rect 67822 273400 67878 273456
rect 67638 272720 67694 272776
rect 67454 272040 67510 272096
rect 67362 250280 67418 250336
rect 67270 241576 67326 241632
rect 67730 271360 67786 271416
rect 67638 270680 67694 270736
rect 67638 270000 67694 270056
rect 67730 269320 67786 269376
rect 67730 268640 67786 268696
rect 67638 267960 67694 268016
rect 67638 267280 67694 267336
rect 67730 266600 67786 266656
rect 67638 265240 67694 265296
rect 67730 264560 67786 264616
rect 67638 263880 67694 263936
rect 67730 263200 67786 263256
rect 67638 262520 67694 262576
rect 67730 261840 67786 261896
rect 67638 261160 67694 261216
rect 67638 260480 67694 260536
rect 67730 259800 67786 259856
rect 67730 259120 67786 259176
rect 67638 257760 67694 257816
rect 67730 256400 67786 256456
rect 67638 255720 67694 255776
rect 67638 255040 67694 255096
rect 67730 254360 67786 254416
rect 67638 253680 67694 253736
rect 67546 252320 67602 252376
rect 67638 251640 67694 251696
rect 67638 250960 67694 251016
rect 67638 249600 67694 249656
rect 68006 248920 68062 248976
rect 67638 248240 67694 248296
rect 67730 247560 67786 247616
rect 67638 246880 67694 246936
rect 68098 246200 68154 246256
rect 67638 245556 67640 245576
rect 67640 245556 67692 245576
rect 67692 245556 67694 245576
rect 67638 245520 67694 245556
rect 67546 244840 67602 244896
rect 67638 244196 67640 244216
rect 67640 244196 67692 244216
rect 67692 244196 67694 244216
rect 67638 244160 67694 244196
rect 67730 243480 67786 243536
rect 67730 242800 67786 242856
rect 67638 242120 67694 242176
rect 67638 241460 67694 241496
rect 67638 241440 67640 241460
rect 67640 241440 67692 241460
rect 67692 241440 67694 241460
rect 67638 240780 67694 240816
rect 67638 240760 67640 240780
rect 67640 240760 67692 240780
rect 67692 240760 67694 240780
rect 71962 295296 72018 295352
rect 73066 295296 73122 295352
rect 80702 402192 80758 402248
rect 77942 309032 77998 309088
rect 78586 309032 78642 309088
rect 77942 307808 77998 307864
rect 75274 294208 75330 294264
rect 75826 294208 75882 294264
rect 77758 292712 77814 292768
rect 84842 400832 84898 400888
rect 80702 295976 80758 296032
rect 88982 399472 89038 399528
rect 98826 400832 98882 400888
rect 92570 292576 92626 292632
rect 97722 295976 97778 296032
rect 97722 295432 97778 295488
rect 98734 364928 98790 364984
rect 104990 403552 105046 403608
rect 108486 402192 108542 402248
rect 116582 391176 116638 391232
rect 104162 298152 104218 298208
rect 106738 295568 106794 295624
rect 109130 302232 109186 302288
rect 110326 302232 110382 302288
rect 113822 370504 113878 370560
rect 110878 299512 110934 299568
rect 111706 299512 111762 299568
rect 112442 297608 112498 297664
rect 116674 296792 116730 296848
rect 117226 297608 117282 297664
rect 117686 294072 117742 294128
rect 117226 293936 117282 293992
rect 117226 292032 117282 292088
rect 119710 295568 119766 295624
rect 118974 293936 119030 293992
rect 118606 291896 118662 291952
rect 69110 288360 69166 288416
rect 120170 291896 120226 291952
rect 120078 278160 120134 278216
rect 69018 265376 69074 265432
rect 69018 258440 69074 258496
rect 68926 210296 68982 210352
rect 66166 181328 66222 181384
rect 120262 286320 120318 286376
rect 120170 261840 120226 261896
rect 120170 250960 120226 251016
rect 120630 250960 120686 251016
rect 119986 248648 120042 248704
rect 120078 241440 120134 241496
rect 119894 241168 119950 241224
rect 70674 239808 70730 239864
rect 73894 238584 73950 238640
rect 72606 238448 72662 238504
rect 81622 238448 81678 238504
rect 82266 238176 82322 238232
rect 93214 235864 93270 235920
rect 93766 235864 93822 235920
rect 100666 177520 100722 177576
rect 106186 177520 106242 177576
rect 107566 177520 107622 177576
rect 97814 176704 97870 176760
rect 99194 176704 99250 176760
rect 100758 176724 100814 176760
rect 100758 176704 100760 176724
rect 100760 176704 100812 176724
rect 100812 176704 100814 176724
rect 108118 176740 108120 176760
rect 108120 176740 108172 176760
rect 108172 176740 108174 176760
rect 108118 176704 108174 176740
rect 110050 176704 110106 176760
rect 69018 175888 69074 175944
rect 121550 291080 121606 291136
rect 121642 290400 121698 290456
rect 121550 289756 121552 289776
rect 121552 289756 121604 289776
rect 121604 289756 121606 289776
rect 121550 289720 121606 289756
rect 121642 289040 121698 289096
rect 121550 287680 121606 287736
rect 121458 284280 121514 284336
rect 121458 283620 121514 283656
rect 121458 283600 121460 283620
rect 121460 283600 121512 283620
rect 121512 283600 121514 283620
rect 121550 282240 121606 282296
rect 121458 281580 121514 281616
rect 121458 281560 121460 281580
rect 121460 281560 121512 281580
rect 121512 281560 121514 281580
rect 121366 280880 121422 280936
rect 121458 280220 121514 280256
rect 121458 280200 121460 280220
rect 121460 280200 121512 280220
rect 121512 280200 121514 280220
rect 121458 278840 121514 278896
rect 121550 277480 121606 277536
rect 121458 276800 121514 276856
rect 121458 276120 121514 276176
rect 121458 275440 121514 275496
rect 121550 274760 121606 274816
rect 121458 274080 121514 274136
rect 121458 273420 121514 273456
rect 121458 273400 121460 273420
rect 121460 273400 121512 273420
rect 121512 273400 121514 273420
rect 121458 272720 121514 272776
rect 121734 287000 121790 287056
rect 121458 271360 121514 271416
rect 121458 270000 121514 270056
rect 121550 269320 121606 269376
rect 121458 268640 121514 268696
rect 121458 267960 121514 268016
rect 122470 284980 122526 285016
rect 122470 284960 122472 284980
rect 122472 284960 122524 284980
rect 122524 284960 122526 284980
rect 125598 386960 125654 387016
rect 122746 285640 122802 285696
rect 122746 282920 122802 282976
rect 122654 279520 122710 279576
rect 122470 278160 122526 278216
rect 122194 272040 122250 272096
rect 122102 266600 122158 266656
rect 121642 265920 121698 265976
rect 121458 265240 121514 265296
rect 121458 263880 121514 263936
rect 121458 263200 121514 263256
rect 121550 262520 121606 262576
rect 120906 261840 120962 261896
rect 121458 261160 121514 261216
rect 121458 260480 121514 260536
rect 121458 259800 121514 259856
rect 122102 259120 122158 259176
rect 121458 258440 121514 258496
rect 121550 257760 121606 257816
rect 121458 257080 121514 257136
rect 121458 256400 121514 256456
rect 121458 255720 121514 255776
rect 121458 254360 121514 254416
rect 121458 253680 121514 253736
rect 121550 253000 121606 253056
rect 121550 252320 121606 252376
rect 121458 251640 121514 251696
rect 121458 250280 121514 250336
rect 121458 249636 121460 249656
rect 121460 249636 121512 249656
rect 121512 249636 121514 249656
rect 121458 249600 121514 249636
rect 120906 249056 120962 249112
rect 121550 248920 121606 248976
rect 121550 248240 121606 248296
rect 121458 247560 121514 247616
rect 121550 246880 121606 246936
rect 121458 246200 121514 246256
rect 121550 245520 121606 245576
rect 121458 244840 121514 244896
rect 121458 244180 121514 244216
rect 121458 244160 121460 244180
rect 121460 244160 121512 244180
rect 121512 244160 121514 244180
rect 121642 243480 121698 243536
rect 121458 242836 121460 242856
rect 121460 242836 121512 242856
rect 121512 242836 121514 242856
rect 121458 242800 121514 242836
rect 121550 242120 121606 242176
rect 121458 240760 121514 240816
rect 121642 240080 121698 240136
rect 115846 192616 115902 192672
rect 113086 191120 113142 191176
rect 114374 182144 114430 182200
rect 112626 177520 112682 177576
rect 114374 177520 114430 177576
rect 121642 235864 121698 235920
rect 122286 267280 122342 267336
rect 122194 255040 122250 255096
rect 122194 230424 122250 230480
rect 122470 264560 122526 264616
rect 124310 296792 124366 296848
rect 125782 205572 125784 205592
rect 125784 205572 125836 205592
rect 125836 205572 125838 205592
rect 125782 205536 125838 205572
rect 130382 389816 130438 389872
rect 133786 262792 133842 262848
rect 130382 184184 130438 184240
rect 114466 177248 114522 177304
rect 115846 177112 115902 177168
rect 116950 177112 117006 177168
rect 121182 177520 121238 177576
rect 124126 177520 124182 177576
rect 124954 177112 125010 177168
rect 135166 289040 135222 289096
rect 135994 368600 136050 368656
rect 140594 405048 140650 405104
rect 140042 401648 140098 401704
rect 138754 189624 138810 189680
rect 134522 180104 134578 180160
rect 127806 177520 127862 177576
rect 142986 300872 143042 300928
rect 146298 322924 146354 322960
rect 146298 322904 146300 322924
rect 146300 322904 146352 322924
rect 146352 322904 146354 322924
rect 147494 244316 147550 244352
rect 147494 244296 147496 244316
rect 147496 244296 147548 244316
rect 147548 244296 147550 244316
rect 152462 217912 152518 217968
rect 154394 283464 154450 283520
rect 156602 298152 156658 298208
rect 155222 184320 155278 184376
rect 149794 181600 149850 181656
rect 157246 239400 157302 239456
rect 158626 283464 158682 283520
rect 158258 240080 158314 240136
rect 158166 199960 158222 200016
rect 164882 297336 164938 297392
rect 163594 240760 163650 240816
rect 159362 185680 159418 185736
rect 156602 177248 156658 177304
rect 148230 177112 148286 177168
rect 118422 176704 118478 176760
rect 125782 176704 125838 176760
rect 128174 176704 128230 176760
rect 130750 176704 130806 176760
rect 132038 176704 132094 176760
rect 134430 176704 134486 176760
rect 135718 176704 135774 176760
rect 159270 176704 159326 176760
rect 104622 175344 104678 175400
rect 165066 295432 165122 295488
rect 166262 292576 166318 292632
rect 165526 269184 165582 269240
rect 165526 228248 165582 228304
rect 164974 214512 165030 214568
rect 162122 176024 162178 176080
rect 121918 175344 121974 175400
rect 129462 175344 129518 175400
rect 133142 175344 133198 175400
rect 119434 174936 119490 174992
rect 66166 129240 66222 129296
rect 65522 128016 65578 128072
rect 66074 122576 66130 122632
rect 66074 102312 66130 102368
rect 67638 126248 67694 126304
rect 67546 125160 67602 125216
rect 67454 123528 67510 123584
rect 67362 120808 67418 120864
rect 67270 100680 67326 100736
rect 67362 89664 67418 89720
rect 168194 356088 168250 356144
rect 168286 293936 168342 293992
rect 168010 171536 168066 171592
rect 170678 239536 170734 239592
rect 176382 373224 176438 373280
rect 176290 371864 176346 371920
rect 175186 362208 175242 362264
rect 171506 182824 171562 182880
rect 170494 179968 170550 180024
rect 151726 94832 151782 94888
rect 94962 94696 95018 94752
rect 113178 94696 113234 94752
rect 115846 94696 115902 94752
rect 126518 94696 126574 94752
rect 130750 93608 130806 93664
rect 97262 93472 97318 93528
rect 113822 93472 113878 93528
rect 110142 93200 110198 93256
rect 87142 92384 87198 92440
rect 98182 92420 98184 92440
rect 98184 92420 98236 92440
rect 98236 92420 98238 92440
rect 98182 92384 98238 92420
rect 98642 92384 98698 92440
rect 107382 92384 107438 92440
rect 75366 91160 75422 91216
rect 85486 91160 85542 91216
rect 86406 91160 86462 91216
rect 86866 91160 86922 91216
rect 89626 91160 89682 91216
rect 90638 91160 90694 91216
rect 92386 91160 92442 91216
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97906 91160 97962 91216
rect 99746 91704 99802 91760
rect 99286 91160 99342 91216
rect 101954 91296 102010 91352
rect 104806 91296 104862 91352
rect 100666 91160 100722 91216
rect 101678 91160 101734 91216
rect 101678 85448 101734 85504
rect 102046 91160 102102 91216
rect 102966 91160 103022 91216
rect 103334 91160 103390 91216
rect 104714 91160 104770 91216
rect 102046 80008 102102 80064
rect 108946 91296 109002 91352
rect 105726 91160 105782 91216
rect 107474 91160 107530 91216
rect 108854 91160 108910 91216
rect 109774 91160 109830 91216
rect 116766 92384 116822 92440
rect 120354 92404 120410 92440
rect 120354 92384 120356 92404
rect 120356 92384 120408 92404
rect 120408 92384 120410 92404
rect 124034 92384 124090 92440
rect 125782 92420 125784 92440
rect 125784 92420 125836 92440
rect 125836 92420 125838 92440
rect 125782 92384 125838 92420
rect 129462 92384 129518 92440
rect 133142 92384 133198 92440
rect 135718 92384 135774 92440
rect 151542 92384 151598 92440
rect 152094 92384 152150 92440
rect 117134 91704 117190 91760
rect 110326 91568 110382 91624
rect 112442 91296 112498 91352
rect 111062 91160 111118 91216
rect 111706 91160 111762 91216
rect 109774 88168 109830 88224
rect 113086 91160 113142 91216
rect 115294 91160 115350 91216
rect 115846 91160 115902 91216
rect 122838 91432 122894 91488
rect 118054 91160 118110 91216
rect 118606 91160 118662 91216
rect 119894 91160 119950 91216
rect 121366 91160 121422 91216
rect 121918 91160 121974 91216
rect 122746 91160 122802 91216
rect 125414 91296 125470 91352
rect 124126 91160 124182 91216
rect 125506 91160 125562 91216
rect 126886 91160 126942 91216
rect 132222 91568 132278 91624
rect 151358 91568 151414 91624
rect 134798 91160 134854 91216
rect 168286 111732 168288 111752
rect 168288 111732 168340 111752
rect 168340 111732 168342 111752
rect 168286 111696 168342 111732
rect 167826 110064 167882 110120
rect 168102 108704 168158 108760
rect 170402 88168 170458 88224
rect 175002 237088 175058 237144
rect 125874 3304 125930 3360
rect 135258 12960 135314 13016
rect 176658 348064 176714 348120
rect 176658 345480 176714 345536
rect 177670 342216 177726 342272
rect 176658 341264 176714 341320
rect 176658 339224 176714 339280
rect 176566 336640 176622 336696
rect 176658 334620 176714 334656
rect 176658 334600 176660 334620
rect 176660 334600 176712 334620
rect 176712 334600 176714 334620
rect 176658 332560 176714 332616
rect 176566 327664 176622 327720
rect 176474 301144 176530 301200
rect 176382 263880 176438 263936
rect 176382 250824 176438 250880
rect 176382 240216 176438 240272
rect 175922 95104 175978 95160
rect 176658 325760 176714 325816
rect 177578 321580 177580 321600
rect 177580 321580 177632 321600
rect 177632 321580 177634 321600
rect 177578 321544 177634 321580
rect 176658 312704 176714 312760
rect 176658 310120 176714 310176
rect 176658 306076 176660 306096
rect 176660 306076 176712 306096
rect 176712 306076 176714 306096
rect 176658 306040 176714 306076
rect 176658 299240 176714 299296
rect 176658 297064 176714 297120
rect 176658 295024 176714 295080
rect 176658 290436 176660 290456
rect 176660 290436 176712 290456
rect 176712 290436 176714 290456
rect 176658 290400 176714 290436
rect 176658 288260 176660 288280
rect 176660 288260 176712 288280
rect 176712 288260 176714 288280
rect 176658 288224 176714 288260
rect 177302 286184 177358 286240
rect 176658 283600 176714 283656
rect 176658 281560 176714 281616
rect 176658 279520 176714 279576
rect 176658 277480 176714 277536
rect 176658 274780 176714 274816
rect 176658 274760 176660 274780
rect 176660 274760 176712 274780
rect 176712 274760 176714 274780
rect 176658 272584 176714 272640
rect 176658 268504 176714 268560
rect 176658 265920 176714 265976
rect 176658 261704 176714 261760
rect 176658 256944 176714 257000
rect 176658 255040 176714 255096
rect 176658 246064 176714 246120
rect 176658 241984 176714 242040
rect 177854 343440 177910 343496
rect 177854 342216 177910 342272
rect 177854 330384 177910 330440
rect 177762 259664 177818 259720
rect 179142 355272 179198 355328
rect 178682 354864 178738 354920
rect 179234 354320 179290 354376
rect 179142 318960 179198 319016
rect 179142 316784 179198 316840
rect 177946 303864 178002 303920
rect 180798 368464 180854 368520
rect 184938 357448 184994 357504
rect 186962 355272 187018 355328
rect 191746 360168 191802 360224
rect 225694 402192 225750 402248
rect 200118 354728 200174 354784
rect 228362 366288 228418 366344
rect 238022 389136 238078 389192
rect 238666 389136 238722 389192
rect 233790 358808 233846 358864
rect 244186 579808 244242 579864
rect 245014 586608 245070 586664
rect 244278 543088 244334 543144
rect 244186 532888 244242 532944
rect 244186 398656 244242 398712
rect 244370 418648 244426 418704
rect 245750 583208 245806 583264
rect 245658 576408 245714 576464
rect 245658 573008 245714 573064
rect 245658 569608 245714 569664
rect 245566 562808 245622 562864
rect 245014 558184 245070 558240
rect 245658 556688 245714 556744
rect 245290 543088 245346 543144
rect 245934 566208 245990 566264
rect 245934 560088 245990 560144
rect 245934 553288 245990 553344
rect 245934 549888 245990 549944
rect 245934 546508 245990 546544
rect 245934 546488 245936 546508
rect 245936 546488 245988 546508
rect 245988 546488 245990 546508
rect 246946 540232 247002 540288
rect 245842 536288 245898 536344
rect 246854 529488 246910 529544
rect 245842 526088 245898 526144
rect 245842 525000 245898 525056
rect 245842 522688 245898 522744
rect 245842 519288 245898 519344
rect 245842 515888 245898 515944
rect 245658 512488 245714 512544
rect 245014 492768 245070 492824
rect 245842 509768 245898 509824
rect 245842 506368 245898 506424
rect 245842 499568 245898 499624
rect 245842 496168 245898 496224
rect 245842 485968 245898 486024
rect 245750 482568 245806 482624
rect 245750 475768 245806 475824
rect 245842 472368 245898 472424
rect 245842 468968 245898 469024
rect 245842 465568 245898 465624
rect 245842 462168 245898 462224
rect 245842 459448 245898 459504
rect 245842 456048 245898 456104
rect 245842 452648 245898 452704
rect 245842 445848 245898 445904
rect 245842 439048 245898 439104
rect 245750 435648 245806 435704
rect 245842 432248 245898 432304
rect 245750 428848 245806 428904
rect 245842 425448 245898 425504
rect 245750 422048 245806 422104
rect 245842 415248 245898 415304
rect 245842 411848 245898 411904
rect 245842 409148 245898 409184
rect 245842 409128 245844 409148
rect 245844 409128 245896 409148
rect 245896 409128 245898 409148
rect 245842 405728 245898 405784
rect 246946 502968 247002 503024
rect 246394 442448 246450 442504
rect 248418 557368 248474 557424
rect 246578 399880 246634 399936
rect 249706 557368 249762 557424
rect 267646 702480 267702 702536
rect 252466 357448 252522 357504
rect 260746 360848 260802 360904
rect 271142 586336 271198 586392
rect 280802 398248 280858 398304
rect 281446 398248 281502 398304
rect 282090 358672 282146 358728
rect 282826 358672 282882 358728
rect 282090 357584 282146 357640
rect 293866 594904 293922 594960
rect 291106 355952 291162 356008
rect 291842 355000 291898 355056
rect 291842 354728 291898 354784
rect 291198 354592 291254 354648
rect 293866 464344 293922 464400
rect 292578 354592 292634 354648
rect 179878 349968 179934 350024
rect 179510 314812 179566 314868
rect 179510 308012 179566 308068
rect 179234 292304 179290 292360
rect 179418 270544 179474 270600
rect 179326 252864 179382 252920
rect 293314 354492 293316 354512
rect 293316 354492 293368 354512
rect 293368 354492 293370 354512
rect 293314 354456 293370 354492
rect 293130 331880 293186 331936
rect 293866 331880 293922 331936
rect 293130 325760 293186 325816
rect 293038 276936 293094 276992
rect 179694 270612 179750 270668
rect 293038 258848 293094 258904
rect 179510 243480 179566 243536
rect 271142 240624 271198 240680
rect 182822 240216 182878 240272
rect 180798 214376 180854 214432
rect 182086 214376 182142 214432
rect 182086 213968 182142 214024
rect 185582 239536 185638 239592
rect 187698 222128 187754 222184
rect 188986 222128 189042 222184
rect 185582 221448 185638 221504
rect 188986 220904 189042 220960
rect 208398 220768 208454 220824
rect 209686 220768 209742 220824
rect 207754 92248 207810 92304
rect 211802 227024 211858 227080
rect 210422 199280 210478 199336
rect 211802 184184 211858 184240
rect 214562 239400 214618 239456
rect 213918 175616 213974 175672
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 213918 173576 213974 173632
rect 214102 172896 214158 172952
rect 213918 172216 213974 172272
rect 214010 171536 214066 171592
rect 213918 171028 213920 171048
rect 213920 171028 213972 171048
rect 213972 171028 213974 171048
rect 213918 170992 213974 171028
rect 213918 169668 213920 169688
rect 213920 169668 213972 169688
rect 213972 169668 213974 169688
rect 213918 169632 213974 169668
rect 214010 168952 214066 169008
rect 213918 168308 213920 168328
rect 213920 168308 213972 168328
rect 213972 168308 213974 168328
rect 213918 168272 213974 168308
rect 214010 167592 214066 167648
rect 213918 166932 213974 166968
rect 213918 166912 213920 166932
rect 213920 166912 213972 166932
rect 213972 166912 213974 166932
rect 214102 166368 214158 166424
rect 214010 165688 214066 165744
rect 213918 165008 213974 165064
rect 213918 163648 213974 163704
rect 214010 162968 214066 163024
rect 213918 161744 213974 161800
rect 213918 161064 213974 161120
rect 214010 160384 214066 160440
rect 213918 159704 213974 159760
rect 214010 159024 214066 159080
rect 213458 157800 213514 157856
rect 213458 157392 213514 157448
rect 214102 157120 214158 157176
rect 213918 156440 213974 156496
rect 213918 155760 213974 155816
rect 214562 155080 214618 155136
rect 214010 154400 214066 154456
rect 213918 153720 213974 153776
rect 213918 153040 213974 153096
rect 214010 152496 214066 152552
rect 213918 151836 213974 151872
rect 213918 151816 213920 151836
rect 213920 151816 213972 151836
rect 213972 151816 213974 151836
rect 214010 151136 214066 151192
rect 213918 150492 213920 150512
rect 213920 150492 213972 150512
rect 213972 150492 213974 150512
rect 213918 150456 213974 150492
rect 214930 170312 214986 170368
rect 214654 149776 214710 149832
rect 213918 149096 213974 149152
rect 213918 148416 213974 148472
rect 214562 147872 214618 147928
rect 213918 147192 213974 147248
rect 214010 145832 214066 145888
rect 213918 145152 213974 145208
rect 213918 144472 213974 144528
rect 213918 143248 213974 143304
rect 213918 142568 213974 142624
rect 214010 141888 214066 141944
rect 213918 141208 213974 141264
rect 213182 140528 213238 140584
rect 213918 139848 213974 139904
rect 213918 138624 213974 138680
rect 214102 137944 214158 138000
rect 213918 137264 213974 137320
rect 214010 136584 214066 136640
rect 214102 135904 214158 135960
rect 213918 135224 213974 135280
rect 214010 134544 214066 134600
rect 213918 133900 213920 133920
rect 213920 133900 213972 133920
rect 213972 133900 213974 133920
rect 213918 133864 213974 133900
rect 214010 133320 214066 133376
rect 213918 132640 213974 132696
rect 213274 131280 213330 131336
rect 213918 130600 213974 130656
rect 213918 128696 213974 128752
rect 213918 127336 213974 127392
rect 214010 126656 214066 126712
rect 213918 125976 213974 126032
rect 214010 125296 214066 125352
rect 213918 124616 213974 124672
rect 214010 124072 214066 124128
rect 213918 123392 213974 123448
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 214010 121352 214066 121408
rect 213918 120672 213974 120728
rect 214010 119992 214066 120048
rect 213918 119448 213974 119504
rect 214102 118804 214104 118824
rect 214104 118804 214156 118824
rect 214156 118804 214158 118824
rect 214102 118768 214158 118804
rect 214010 118088 214066 118144
rect 213918 117408 213974 117464
rect 214010 116728 214066 116784
rect 213918 116068 213974 116104
rect 213918 116048 213920 116068
rect 213920 116048 213972 116068
rect 213972 116048 213974 116068
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 214010 114144 214066 114200
rect 213918 113464 213974 113520
rect 214010 112784 214066 112840
rect 213918 112104 213974 112160
rect 213918 111424 213974 111480
rect 214010 110200 214066 110256
rect 213918 109520 213974 109576
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 214010 107480 214066 107536
rect 213918 106800 213974 106856
rect 213918 106120 213974 106176
rect 214010 105576 214066 105632
rect 213918 104916 213974 104952
rect 213918 104896 213920 104916
rect 213920 104896 213972 104916
rect 213972 104896 213974 104916
rect 214010 104216 214066 104272
rect 213918 103556 213974 103592
rect 213918 103536 213920 103556
rect 213920 103536 213972 103556
rect 213972 103536 213974 103556
rect 214010 102856 214066 102912
rect 213918 102196 213974 102232
rect 213918 102176 213920 102196
rect 213920 102176 213972 102196
rect 213972 102176 213974 102196
rect 214654 146512 214710 146568
rect 214838 128016 214894 128072
rect 214746 110744 214802 110800
rect 213918 100952 213974 101008
rect 214010 100272 214066 100328
rect 213918 99592 213974 99648
rect 214010 98912 214066 98968
rect 213918 98232 213974 98288
rect 213918 97552 213974 97608
rect 214562 96872 214618 96928
rect 213918 96328 213974 96384
rect 214562 88984 214618 89040
rect 215022 101496 215078 101552
rect 215022 89664 215078 89720
rect 232502 178880 232558 178936
rect 242254 237904 242310 237960
rect 239402 235184 239458 235240
rect 259366 233144 259422 233200
rect 264978 238448 265034 238504
rect 265530 236952 265586 237008
rect 264058 236000 264114 236056
rect 265530 236000 265586 236056
rect 262126 232464 262182 232520
rect 253938 224848 253994 224904
rect 246302 178744 246358 178800
rect 245658 177520 245714 177576
rect 247866 177792 247922 177848
rect 246946 175752 247002 175808
rect 249062 172488 249118 172544
rect 249246 175208 249302 175264
rect 249154 171808 249210 171864
rect 249338 171400 249394 171456
rect 249798 154400 249854 154456
rect 249982 176024 250038 176080
rect 249982 173712 250038 173768
rect 250074 170856 250130 170912
rect 251178 159568 251234 159624
rect 251178 153448 251234 153504
rect 250626 149640 250682 149696
rect 249890 149232 249946 149288
rect 240138 15136 240194 15192
rect 240782 15136 240838 15192
rect 245658 86128 245714 86184
rect 249798 96600 249854 96656
rect 251454 164328 251510 164384
rect 251362 160520 251418 160576
rect 252466 170448 252522 170504
rect 252466 169088 252522 169144
rect 252374 168544 252430 168600
rect 252466 168136 252522 168192
rect 252374 167592 252430 167648
rect 252006 167184 252062 167240
rect 251914 166268 251916 166288
rect 251916 166268 251968 166288
rect 251968 166268 251970 166288
rect 251914 166232 251970 166268
rect 252466 166640 252522 166696
rect 252374 165688 252430 165744
rect 252466 165280 252522 165336
rect 251914 164736 251970 164792
rect 251914 163376 251970 163432
rect 252190 162968 252246 163024
rect 252098 162424 252154 162480
rect 252466 162016 252522 162072
rect 252466 161508 252468 161528
rect 252468 161508 252520 161528
rect 252520 161508 252522 161528
rect 252466 161472 252522 161508
rect 252466 161064 252522 161120
rect 251914 160112 251970 160168
rect 251638 159160 251694 159216
rect 252466 158208 252522 158264
rect 252374 157800 252430 157856
rect 252466 156848 252522 156904
rect 251546 156304 251602 156360
rect 252466 155916 252522 155952
rect 252466 155896 252468 155916
rect 252468 155896 252520 155916
rect 252520 155896 252522 155916
rect 252466 155352 252522 155408
rect 252374 154944 252430 155000
rect 251730 153992 251786 154048
rect 252466 153076 252468 153096
rect 252468 153076 252520 153096
rect 252520 153076 252522 153096
rect 252466 153040 252522 153076
rect 252006 152088 252062 152144
rect 252466 151700 252522 151736
rect 252466 151680 252468 151700
rect 252468 151680 252520 151700
rect 252520 151680 252522 151700
rect 252374 150728 252430 150784
rect 251914 150184 251970 150240
rect 251546 149776 251602 149832
rect 252742 169496 252798 169552
rect 252650 151136 252706 151192
rect 252374 148824 252430 148880
rect 251270 147872 251326 147928
rect 251178 146956 251180 146976
rect 251180 146956 251232 146976
rect 251232 146956 251234 146976
rect 251178 146920 251234 146956
rect 251546 144608 251602 144664
rect 251914 145968 251970 146024
rect 252466 148280 252522 148336
rect 252466 147484 252522 147520
rect 252466 147464 252468 147484
rect 252468 147464 252520 147484
rect 252520 147464 252522 147484
rect 252374 146512 252430 146568
rect 251730 143112 251786 143168
rect 251086 142568 251142 142624
rect 250626 136992 250682 137048
rect 251730 141344 251786 141400
rect 251730 139476 251732 139496
rect 251732 139476 251784 139496
rect 251784 139476 251786 139496
rect 251730 139440 251786 139476
rect 251730 138488 251786 138544
rect 251362 137944 251418 138000
rect 251730 135632 251786 135688
rect 251454 134680 251510 134736
rect 251362 133728 251418 133784
rect 251546 131824 251602 131880
rect 251454 129104 251510 129160
rect 251638 127608 251694 127664
rect 251362 124344 251418 124400
rect 251178 122984 251234 123040
rect 252466 145560 252522 145616
rect 252098 145016 252154 145072
rect 252466 144084 252522 144120
rect 252466 144064 252468 144084
rect 252468 144064 252520 144084
rect 252520 144064 252522 144084
rect 252650 144064 252706 144120
rect 252190 143656 252246 143712
rect 252466 142704 252522 142760
rect 251914 127200 251970 127256
rect 251914 125332 251916 125352
rect 251916 125332 251968 125352
rect 251968 125332 251970 125352
rect 251914 125296 251970 125332
rect 252466 138896 252522 138952
rect 252466 137536 252522 137592
rect 252466 136176 252522 136232
rect 252374 135224 252430 135280
rect 252466 134272 252522 134328
rect 252374 133320 252430 133376
rect 252466 132776 252522 132832
rect 252466 132404 252468 132424
rect 252468 132404 252520 132424
rect 252520 132404 252522 132424
rect 252466 132368 252522 132404
rect 252098 131416 252154 131472
rect 252466 130872 252522 130928
rect 252466 130500 252468 130520
rect 252468 130500 252520 130520
rect 252520 130500 252522 130520
rect 252466 130464 252522 130500
rect 252374 130056 252430 130112
rect 252466 129512 252522 129568
rect 252374 128560 252430 128616
rect 252466 128188 252468 128208
rect 252468 128188 252520 128208
rect 252520 128188 252522 128208
rect 252466 128152 252522 128188
rect 252098 125704 252154 125760
rect 252466 126656 252522 126712
rect 251362 122032 251418 122088
rect 251362 119584 251418 119640
rect 251822 120536 251878 120592
rect 251822 117816 251878 117872
rect 251730 117272 251786 117328
rect 251362 116864 251418 116920
rect 252006 121488 252062 121544
rect 251730 114416 251786 114472
rect 251638 114008 251694 114064
rect 251362 113464 251418 113520
rect 251914 114960 251970 115016
rect 251638 112104 251694 112160
rect 251086 109112 251142 109168
rect 251362 105032 251418 105088
rect 252466 124752 252522 124808
rect 252466 123936 252522 123992
rect 252374 123392 252430 123448
rect 252466 122440 252522 122496
rect 252466 121080 252522 121136
rect 252282 120128 252338 120184
rect 252282 118768 252338 118824
rect 252466 119176 252522 119232
rect 252466 118224 252522 118280
rect 252374 116320 252430 116376
rect 252466 115912 252522 115968
rect 252282 115368 252338 115424
rect 252466 113056 252522 113112
rect 252466 112648 252522 112704
rect 252098 111696 252154 111752
rect 252006 111152 252062 111208
rect 251914 110200 251970 110256
rect 252098 109248 252154 109304
rect 251822 106936 251878 106992
rect 251914 105984 251970 106040
rect 251914 104624 251970 104680
rect 251730 103672 251786 103728
rect 252466 109792 252522 109848
rect 252466 108876 252468 108896
rect 252468 108876 252520 108896
rect 252520 108876 252522 108896
rect 252466 108840 252522 108876
rect 252374 108296 252430 108352
rect 252282 107888 252338 107944
rect 252190 107480 252246 107536
rect 252098 106528 252154 106584
rect 252466 105576 252522 105632
rect 251730 99864 251786 99920
rect 251178 98912 251234 98968
rect 251822 98504 251878 98560
rect 251546 97960 251602 98016
rect 252006 103128 252062 103184
rect 252466 104080 252522 104136
rect 252374 102720 252430 102776
rect 252466 102176 252522 102232
rect 252282 101768 252338 101824
rect 252006 100852 252008 100872
rect 252008 100852 252060 100872
rect 252060 100852 252062 100872
rect 252006 100816 252062 100852
rect 251178 97008 251234 97064
rect 251914 97008 251970 97064
rect 251270 96192 251326 96248
rect 252466 101360 252522 101416
rect 252466 100408 252522 100464
rect 252374 99456 252430 99512
rect 252190 97588 252192 97608
rect 252192 97588 252244 97608
rect 252244 97588 252246 97608
rect 252190 97552 252246 97588
rect 252098 96600 252154 96656
rect 252374 3440 252430 3496
rect 257618 152904 257674 152960
rect 258262 3440 258318 3496
rect 261206 176604 261208 176624
rect 261208 176604 261260 176624
rect 261260 176604 261262 176624
rect 261206 176568 261262 176604
rect 262126 21936 262182 21992
rect 266266 175888 266322 175944
rect 264978 149640 265034 149696
rect 273994 238720 274050 238776
rect 271786 238448 271842 238504
rect 279422 238312 279478 238368
rect 277950 238176 278006 238232
rect 278686 232464 278742 232520
rect 271234 232056 271290 232112
rect 270406 231104 270462 231160
rect 269118 60052 269120 60072
rect 269120 60052 269172 60072
rect 269172 60052 269174 60072
rect 269118 60016 269174 60052
rect 270038 134408 270094 134464
rect 270406 11736 270462 11792
rect 271786 113872 271842 113928
rect 271694 46860 271696 46880
rect 271696 46860 271748 46880
rect 271748 46860 271750 46880
rect 271694 46824 271750 46860
rect 273902 181328 273958 181384
rect 278134 113736 278190 113792
rect 292946 240488 293002 240544
rect 285586 174528 285642 174584
rect 288530 233144 288586 233200
rect 286966 218592 287022 218648
rect 287978 32408 288034 32464
rect 289726 19252 289728 19272
rect 289728 19252 289780 19272
rect 289780 19252 289782 19272
rect 289726 19216 289782 19252
rect 292670 198076 292726 198112
rect 292670 198056 292672 198076
rect 292672 198056 292724 198076
rect 292724 198056 292726 198076
rect 293866 259120 293922 259176
rect 294326 323040 294382 323096
rect 294050 305380 294106 305416
rect 294050 305360 294052 305380
rect 294052 305360 294104 305380
rect 294104 305360 294106 305380
rect 294050 299240 294106 299296
rect 293958 246200 294014 246256
rect 293314 241848 293370 241904
rect 293314 241168 293370 241224
rect 293222 238448 293278 238504
rect 295430 354320 295486 354376
rect 295430 352280 295486 352336
rect 295430 349560 295486 349616
rect 295430 347520 295486 347576
rect 295430 343440 295486 343496
rect 295430 340720 295486 340776
rect 295430 338680 295486 338736
rect 295430 334328 295486 334384
rect 295430 329840 295486 329896
rect 296718 354592 296774 354648
rect 295614 345480 295670 345536
rect 295522 327800 295578 327856
rect 295338 321000 295394 321056
rect 295338 318960 295394 319016
rect 295338 316920 295394 316976
rect 295338 314200 295394 314256
rect 295338 312160 295394 312216
rect 295338 310120 295394 310176
rect 295338 307828 295394 307864
rect 295338 307808 295340 307828
rect 295340 307808 295392 307828
rect 295392 307808 295394 307828
rect 295338 303320 295394 303376
rect 295338 301280 295394 301336
rect 295338 296520 295394 296576
rect 295338 292476 295340 292496
rect 295340 292476 295392 292496
rect 295392 292476 295394 292496
rect 295338 292440 295394 292476
rect 295338 290400 295394 290456
rect 294786 283600 294842 283656
rect 295246 283600 295302 283656
rect 295338 281580 295394 281616
rect 295338 281560 295340 281580
rect 295340 281560 295392 281580
rect 295392 281560 295394 281580
rect 295338 274760 295394 274816
rect 295338 272720 295394 272776
rect 294234 267960 294290 268016
rect 295338 261180 295394 261216
rect 295338 261160 295340 261180
rect 295340 261160 295392 261180
rect 295392 261160 295394 261180
rect 295338 257080 295394 257136
rect 295338 255040 295394 255096
rect 295338 252320 295394 252376
rect 295338 250280 295394 250336
rect 295338 248240 295394 248296
rect 294326 246200 294382 246256
rect 295706 336640 295762 336696
rect 295982 336640 296038 336696
rect 296166 287136 296222 287192
rect 296626 294480 296682 294536
rect 296534 278840 296590 278896
rect 296074 270408 296130 270464
rect 296350 263508 296352 263528
rect 296352 263508 296404 263528
rect 296404 263508 296406 263528
rect 296350 263472 296406 263508
rect 296258 243480 296314 243536
rect 296442 241460 296498 241496
rect 296442 241440 296444 241460
rect 296444 241440 296496 241460
rect 296496 241440 296498 241460
rect 296718 231240 296774 231296
rect 298006 357856 298062 357912
rect 298190 240760 298246 240816
rect 298006 225528 298062 225584
rect 299478 353232 299534 353288
rect 295338 84224 295394 84280
rect 297362 22616 297418 22672
rect 297362 8200 297418 8256
rect 303526 522280 303582 522336
rect 302238 241848 302294 241904
rect 302238 25472 302294 25528
rect 299570 11736 299626 11792
rect 305090 354864 305146 354920
rect 305550 291760 305606 291816
rect 305090 240216 305146 240272
rect 305642 240216 305698 240272
rect 305090 238720 305146 238776
rect 309230 369824 309286 369880
rect 307666 175616 307722 175672
rect 307022 175208 307078 175264
rect 306930 173168 306986 173224
rect 306562 170584 306618 170640
rect 306562 169224 306618 169280
rect 306562 166776 306618 166832
rect 306378 166368 306434 166424
rect 306470 165824 306526 165880
rect 306470 165416 306526 165472
rect 306378 164600 306434 164656
rect 306378 164228 306380 164248
rect 306380 164228 306432 164248
rect 306432 164228 306434 164248
rect 306378 164192 306434 164228
rect 306562 163784 306618 163840
rect 306378 163376 306434 163432
rect 306470 162968 306526 163024
rect 306470 162424 306526 162480
rect 306378 161608 306434 161664
rect 306562 162016 306618 162072
rect 306470 161200 306526 161256
rect 306378 160792 306434 160848
rect 306562 160384 306618 160440
rect 306562 159976 306618 160032
rect 306378 159568 306434 159624
rect 306470 159024 306526 159080
rect 306562 158616 306618 158672
rect 306378 158208 306434 158264
rect 306470 157800 306526 157856
rect 306930 157392 306986 157448
rect 306746 155624 306802 155680
rect 306654 153176 306710 153232
rect 306562 152632 306618 152688
rect 305734 152224 305790 152280
rect 305642 149232 305698 149288
rect 307482 174800 307538 174856
rect 307574 174392 307630 174448
rect 307666 173984 307722 174040
rect 307666 173576 307722 173632
rect 307298 172660 307300 172680
rect 307300 172660 307352 172680
rect 307352 172660 307354 172680
rect 307298 172624 307354 172660
rect 307574 172216 307630 172272
rect 307482 171400 307538 171456
rect 307666 171808 307722 171864
rect 307298 170992 307354 171048
rect 307666 170176 307722 170232
rect 307666 169788 307722 169824
rect 307666 169768 307668 169788
rect 307668 169768 307720 169788
rect 307720 169768 307722 169788
rect 307666 168816 307722 168872
rect 307298 168408 307354 168464
rect 307114 165008 307170 165064
rect 306562 145016 306618 145072
rect 306562 139984 306618 140040
rect 306746 137808 306802 137864
rect 307482 168000 307538 168056
rect 307574 167592 307630 167648
rect 307666 167204 307722 167240
rect 307666 167184 307668 167204
rect 307668 167184 307720 167204
rect 307720 167184 307722 167204
rect 307482 156984 307538 157040
rect 307574 156576 307630 156632
rect 307666 156168 307722 156224
rect 307482 155216 307538 155272
rect 307390 154808 307446 154864
rect 307574 154400 307630 154456
rect 307482 153584 307538 153640
rect 307666 153992 307722 154048
rect 307666 151852 307668 151872
rect 307668 151852 307720 151872
rect 307720 151852 307722 151872
rect 307666 151816 307722 151852
rect 307482 151408 307538 151464
rect 307298 151000 307354 151056
rect 307666 150592 307722 150648
rect 307482 150184 307538 150240
rect 307666 149776 307722 149832
rect 307574 148824 307630 148880
rect 307482 148008 307538 148064
rect 307666 148416 307722 148472
rect 307574 147600 307630 147656
rect 307482 147192 307538 147248
rect 307482 145832 307538 145888
rect 307206 144608 307262 144664
rect 306746 136584 306802 136640
rect 306562 136176 306618 136232
rect 306930 135632 306986 135688
rect 307114 131008 307170 131064
rect 306562 129240 306618 129296
rect 307114 128832 307170 128888
rect 307114 127608 307170 127664
rect 306746 127200 306802 127256
rect 306746 125840 306802 125896
rect 306746 125432 306802 125488
rect 307022 124616 307078 124672
rect 306562 123800 306618 123856
rect 306746 121216 306802 121272
rect 306562 118224 306618 118280
rect 306746 117000 306802 117056
rect 306930 114416 306986 114472
rect 306562 114008 306618 114064
rect 305642 107616 305698 107672
rect 305734 106256 305790 106312
rect 305918 105440 305974 105496
rect 305826 101088 305882 101144
rect 306746 101632 306802 101688
rect 307114 124228 307170 124264
rect 307114 124208 307116 124228
rect 307116 124208 307168 124228
rect 307168 124208 307170 124228
rect 307114 123392 307170 123448
rect 307114 115640 307170 115696
rect 307666 146784 307722 146840
rect 307666 145424 307722 145480
rect 307390 144200 307446 144256
rect 307298 143384 307354 143440
rect 307298 116184 307354 116240
rect 307206 98640 307262 98696
rect 307482 143792 307538 143848
rect 307666 142976 307722 143032
rect 307482 142432 307538 142488
rect 307666 142024 307722 142080
rect 307574 141208 307630 141264
rect 307666 140820 307722 140856
rect 307666 140800 307668 140820
rect 307668 140800 307720 140820
rect 307720 140800 307722 140820
rect 307574 140392 307630 140448
rect 307666 139576 307722 139632
rect 307482 139032 307538 139088
rect 307666 138624 307722 138680
rect 307574 138216 307630 138272
rect 307666 137400 307722 137456
rect 307666 135224 307722 135280
rect 307482 134816 307538 134872
rect 307574 134408 307630 134464
rect 307666 134036 307668 134056
rect 307668 134036 307720 134056
rect 307720 134036 307722 134056
rect 307666 134000 307722 134036
rect 307482 133592 307538 133648
rect 307574 133184 307630 133240
rect 307666 132660 307722 132696
rect 307666 132640 307668 132660
rect 307668 132640 307720 132660
rect 307720 132640 307722 132660
rect 307482 132232 307538 132288
rect 307574 131824 307630 131880
rect 307666 131416 307722 131472
rect 307574 130600 307630 130656
rect 307482 130192 307538 130248
rect 307666 129784 307722 129840
rect 307666 128016 307722 128072
rect 307666 126792 307722 126848
rect 307666 125024 307722 125080
rect 307666 122984 307722 123040
rect 307482 122440 307538 122496
rect 307574 122032 307630 122088
rect 307666 121644 307722 121680
rect 307666 121624 307668 121644
rect 307668 121624 307720 121644
rect 307720 121624 307722 121644
rect 307574 120808 307630 120864
rect 307666 120400 307722 120456
rect 307574 119992 307630 120048
rect 307482 119584 307538 119640
rect 307666 119040 307722 119096
rect 307574 118632 307630 118688
rect 307666 117816 307722 117872
rect 307666 117428 307722 117464
rect 307666 117408 307668 117428
rect 307668 117408 307720 117428
rect 307720 117408 307722 117428
rect 307482 116592 307538 116648
rect 307574 115232 307630 115288
rect 307666 114824 307722 114880
rect 307666 113212 307722 113248
rect 307666 113192 307668 113212
rect 307668 113192 307720 113212
rect 307720 113192 307722 113212
rect 307482 112240 307538 112296
rect 307666 111868 307668 111888
rect 307668 111868 307720 111888
rect 307720 111868 307722 111888
rect 307666 111832 307722 111868
rect 307482 111424 307538 111480
rect 307574 111016 307630 111072
rect 307666 110608 307722 110664
rect 307482 110200 307538 110256
rect 307574 109792 307630 109848
rect 307666 109248 307722 109304
rect 307482 108840 307538 108896
rect 307666 108432 307722 108488
rect 307574 108024 307630 108080
rect 307482 107616 307538 107672
rect 307666 107616 307722 107672
rect 307482 107208 307538 107264
rect 308494 146376 308550 146432
rect 307574 106800 307630 106856
rect 307666 106428 307668 106448
rect 307668 106428 307720 106448
rect 307720 106428 307722 106448
rect 307666 106392 307722 106428
rect 307482 106256 307538 106312
rect 307574 105848 307630 105904
rect 307666 105052 307722 105088
rect 307666 105032 307668 105052
rect 307668 105032 307720 105052
rect 307720 105032 307722 105052
rect 307482 104624 307538 104680
rect 307666 104216 307722 104272
rect 307574 103808 307630 103864
rect 307574 103400 307630 103456
rect 307482 102992 307538 103048
rect 307666 102448 307722 102504
rect 307482 102040 307538 102096
rect 307574 101224 307630 101280
rect 307482 101088 307538 101144
rect 307666 100816 307722 100872
rect 307574 100408 307630 100464
rect 307666 99592 307722 99648
rect 307574 99048 307630 99104
rect 307666 98232 307722 98288
rect 307666 97416 307722 97472
rect 307574 97008 307630 97064
rect 307666 96636 307668 96656
rect 307668 96636 307720 96656
rect 307720 96636 307722 96656
rect 307666 96600 307722 96636
rect 307666 96192 307722 96248
rect 309230 100136 309286 100192
rect 307758 42064 307814 42120
rect 305642 5480 305698 5536
rect 313922 599120 313978 599176
rect 313186 217368 313242 217424
rect 313186 216688 313242 216744
rect 313922 243480 313978 243536
rect 313922 187176 313978 187232
rect 317418 597896 317474 597952
rect 314658 216688 314714 216744
rect 314474 178880 314530 178936
rect 318154 235864 318210 235920
rect 318706 226888 318762 226944
rect 315946 177384 316002 177440
rect 320086 582936 320142 582992
rect 322202 583888 322258 583944
rect 320822 356088 320878 356144
rect 318154 176160 318210 176216
rect 321466 176024 321522 176080
rect 321282 165008 321338 165064
rect 322754 230424 322810 230480
rect 322846 209772 322902 209808
rect 322846 209752 322848 209772
rect 322848 209752 322900 209772
rect 322900 209752 322902 209772
rect 323122 226888 323178 226944
rect 322938 207032 322994 207088
rect 321558 142840 321614 142896
rect 324410 190984 324466 191040
rect 324318 172388 324320 172408
rect 324320 172388 324372 172408
rect 324372 172388 324374 172408
rect 324318 172352 324374 172388
rect 324318 170040 324374 170096
rect 324318 169360 324374 169416
rect 324410 168544 324466 168600
rect 324318 167728 324374 167784
rect 324318 165416 324374 165472
rect 324318 163920 324374 163976
rect 324410 163104 324466 163160
rect 324318 160792 324374 160848
rect 324594 174664 324650 174720
rect 324502 160112 324558 160168
rect 324318 159296 324374 159352
rect 324318 158480 324374 158536
rect 324410 157800 324466 157856
rect 324318 157020 324320 157040
rect 324320 157020 324372 157040
rect 324372 157020 324374 157040
rect 324318 156984 324374 157020
rect 324410 156304 324466 156360
rect 324686 155488 324742 155544
rect 324318 154672 324374 154728
rect 324318 153992 324374 154048
rect 323214 153176 323270 153232
rect 324318 152360 324374 152416
rect 323030 149368 323086 149424
rect 323306 136992 323362 137048
rect 324318 151716 324320 151736
rect 324320 151716 324372 151736
rect 324372 151716 324374 151736
rect 324318 151680 324374 151716
rect 324318 150864 324374 150920
rect 325606 150048 325662 150104
rect 327354 405592 327410 405648
rect 327354 404912 327410 404968
rect 325790 171672 325846 171728
rect 324318 148552 324374 148608
rect 324410 147736 324466 147792
rect 324318 147056 324374 147112
rect 324318 146260 324374 146296
rect 324318 146240 324320 146260
rect 324320 146240 324372 146260
rect 324372 146240 324374 146260
rect 324410 145424 324466 145480
rect 324318 144780 324320 144800
rect 324320 144780 324372 144800
rect 324372 144780 324374 144800
rect 324318 144744 324374 144780
rect 324410 143928 324466 143984
rect 324318 143112 324374 143168
rect 324318 141616 324374 141672
rect 324410 140800 324466 140856
rect 324318 140120 324374 140176
rect 324318 138488 324374 138544
rect 324318 137808 324374 137864
rect 323398 136312 323454 136368
rect 324318 135496 324374 135552
rect 324318 134680 324374 134736
rect 324410 134000 324466 134056
rect 324318 133184 324374 133240
rect 323490 131824 323546 131880
rect 323490 131144 323546 131200
rect 324318 130872 324374 130928
rect 324410 130056 324466 130112
rect 324318 129412 324320 129432
rect 324320 129412 324372 129432
rect 324372 129412 324374 129432
rect 324318 129376 324374 129412
rect 324410 128560 324466 128616
rect 324318 127744 324374 127800
rect 324410 127064 324466 127120
rect 324318 124752 324374 124808
rect 323490 123392 323546 123448
rect 323490 122848 323546 122904
rect 324318 122440 324374 122496
rect 321650 122168 321706 122224
rect 324318 120808 324374 120864
rect 324410 120128 324466 120184
rect 324318 119312 324374 119368
rect 325606 126248 325662 126304
rect 325974 177248 326030 177304
rect 325882 161608 325938 161664
rect 331126 601704 331182 601760
rect 328366 600480 328422 600536
rect 327814 405592 327870 405648
rect 329102 594768 329158 594824
rect 328366 396616 328422 396672
rect 324962 118496 325018 118552
rect 324318 117816 324374 117872
rect 324318 116320 324374 116376
rect 324318 115504 324374 115560
rect 321558 109112 321614 109168
rect 321466 97280 321522 97336
rect 313738 84768 313794 84824
rect 316038 91704 316094 91760
rect 322938 106256 322994 106312
rect 323306 106256 323362 106312
rect 321650 102720 321706 102776
rect 321742 101088 321798 101144
rect 324318 114008 324374 114064
rect 324410 113192 324466 113248
rect 324962 110880 325018 110936
rect 324318 110064 324374 110120
rect 324410 108568 324466 108624
rect 324318 108296 324374 108352
rect 326342 112376 326398 112432
rect 325054 107072 325110 107128
rect 324318 105440 324374 105496
rect 324502 104760 324558 104816
rect 324318 103944 324374 104000
rect 324318 102448 324374 102504
rect 324410 100816 324466 100872
rect 324318 100136 324374 100192
rect 324410 99320 324466 99376
rect 324318 97008 324374 97064
rect 324502 93744 324558 93800
rect 324410 93608 324466 93664
rect 324318 92384 324374 92440
rect 331126 396752 331182 396808
rect 332598 236000 332654 236056
rect 331402 198736 331458 198792
rect 336094 601840 336150 601896
rect 334622 595040 334678 595096
rect 333334 237224 333390 237280
rect 333334 236000 333390 236056
rect 333242 197240 333298 197296
rect 333242 196016 333298 196072
rect 332782 181464 332838 181520
rect 336002 597624 336058 597680
rect 336554 594496 336610 594552
rect 334622 206896 334678 206952
rect 334622 205672 334678 205728
rect 332046 84768 332102 84824
rect 337106 591776 337162 591832
rect 337658 589056 337714 589112
rect 337658 586336 337714 586392
rect 337658 584296 337714 584352
rect 337658 581576 337714 581632
rect 337658 578856 337714 578912
rect 337658 576852 337660 576872
rect 337660 576852 337712 576872
rect 337712 576852 337714 576872
rect 337658 576816 337714 576852
rect 337842 574096 337898 574152
rect 337658 571376 337714 571432
rect 337658 568676 337714 568712
rect 337658 568656 337660 568676
rect 337660 568656 337712 568676
rect 337712 568656 337714 568676
rect 336922 559136 336978 559192
rect 337658 561176 337714 561232
rect 337382 553696 337438 553752
rect 337382 550976 337438 551032
rect 337658 548936 337714 548992
rect 337382 546488 337438 546544
rect 337382 546216 337438 546272
rect 337290 536016 337346 536072
rect 336830 531256 336886 531312
rect 337658 543496 337714 543552
rect 337474 541456 337530 541512
rect 337658 538736 337714 538792
rect 337658 533296 337714 533352
rect 337934 556416 337990 556472
rect 337842 525816 337898 525872
rect 337474 523776 337530 523832
rect 337474 521056 337530 521112
rect 337658 515616 337714 515672
rect 337658 513576 337714 513632
rect 337658 510856 337714 510912
rect 337106 506096 337162 506152
rect 337658 503376 337714 503432
rect 337750 500656 337806 500712
rect 337658 497936 337714 497992
rect 337474 495896 337530 495952
rect 337474 493176 337530 493232
rect 337658 490456 337714 490512
rect 337750 485696 337806 485752
rect 336738 480256 336794 480312
rect 337934 482976 337990 483032
rect 337750 478216 337806 478272
rect 337658 475496 337714 475552
rect 336830 472776 336886 472832
rect 336738 470736 336794 470792
rect 337658 465296 337714 465352
rect 337658 460536 337714 460592
rect 337658 457816 337714 457872
rect 337658 455096 337714 455152
rect 337566 453056 337622 453112
rect 337290 450336 337346 450392
rect 337106 447616 337162 447672
rect 337290 440136 337346 440192
rect 337290 437416 337346 437472
rect 337382 435376 337438 435432
rect 337658 432656 337714 432712
rect 336922 429936 336978 429992
rect 336922 427216 336978 427272
rect 337658 425176 337714 425232
rect 337658 422456 337714 422512
rect 337842 417696 337898 417752
rect 336830 414976 336886 415032
rect 337382 412256 337438 412312
rect 336922 409536 336978 409592
rect 337658 407496 337714 407552
rect 337750 404776 337806 404832
rect 337474 401648 337530 401704
rect 338946 598984 339002 599040
rect 338762 563896 338818 563952
rect 338026 468016 338082 468072
rect 338026 444896 338082 444952
rect 338026 401648 338082 401704
rect 335450 196016 335506 196072
rect 335634 185544 335690 185600
rect 333242 65456 333298 65512
rect 333242 45464 333298 45520
rect 332690 44240 332746 44296
rect 333242 44240 333298 44296
rect 336830 178744 336886 178800
rect 340326 597760 340382 597816
rect 355138 596400 355194 596456
rect 364798 597896 364854 597952
rect 419538 603200 419594 603256
rect 420182 603200 420238 603256
rect 429198 599120 429254 599176
rect 433614 601840 433670 601896
rect 445850 601704 445906 601760
rect 462594 600480 462650 600536
rect 467194 597760 467250 597816
rect 479338 598984 479394 599040
rect 507858 603064 507914 603120
rect 505742 598984 505798 599040
rect 515402 604424 515458 604480
rect 522946 597760 523002 597816
rect 359646 595040 359702 595096
rect 362222 594904 362278 594960
rect 534170 566616 534226 566672
rect 534078 531256 534134 531312
rect 534078 490456 534134 490512
rect 339314 488416 339370 488472
rect 339406 398792 339462 398848
rect 337474 158752 337530 158808
rect 343638 396752 343694 396808
rect 340142 362752 340198 362808
rect 340142 362208 340198 362264
rect 336830 26188 336832 26208
rect 336832 26188 336884 26208
rect 336884 26188 336886 26208
rect 336830 26152 336886 26188
rect 336830 25472 336886 25528
rect 340142 28872 340198 28928
rect 340142 28192 340198 28248
rect 342442 187040 342498 187096
rect 342994 224440 343050 224496
rect 345754 382880 345810 382936
rect 343730 178608 343786 178664
rect 343822 151000 343878 151056
rect 347778 196560 347834 196616
rect 347226 117292 347282 117328
rect 347226 117272 347228 117292
rect 347228 117272 347280 117292
rect 347280 117272 347282 117292
rect 347870 179968 347926 180024
rect 349250 202136 349306 202192
rect 349250 201456 349306 201512
rect 342902 28872 342958 28928
rect 349894 242120 349950 242176
rect 351182 240760 351238 240816
rect 353298 357448 353354 357504
rect 354678 396616 354734 396672
rect 363602 335960 363658 336016
rect 362958 231784 363014 231840
rect 364154 231784 364210 231840
rect 364706 246200 364762 246256
rect 376758 398384 376814 398440
rect 377954 398384 378010 398440
rect 373722 241848 373778 241904
rect 374642 102720 374698 102776
rect 376942 297064 376998 297120
rect 377402 292984 377458 293040
rect 376942 290944 376998 291000
rect 376942 288904 376998 288960
rect 376942 286864 376998 286920
rect 377310 284144 377366 284200
rect 376942 282104 376998 282160
rect 376942 280220 376998 280256
rect 376942 280200 376944 280220
rect 376944 280200 376996 280220
rect 376996 280200 376998 280220
rect 376758 278024 376814 278080
rect 376942 265104 376998 265160
rect 376114 250144 376170 250200
rect 377310 263200 377366 263256
rect 376942 258984 376998 259040
rect 377310 254360 377366 254416
rect 376942 252184 376998 252240
rect 376942 248104 376998 248160
rect 376942 246064 376998 246120
rect 376666 241984 376722 242040
rect 377954 299240 378010 299296
rect 379150 295160 379206 295216
rect 377770 276020 377772 276040
rect 377772 276020 377824 276040
rect 377824 276020 377826 276040
rect 377770 275984 377826 276020
rect 377770 273944 377826 274000
rect 378046 254360 378102 254416
rect 377954 244024 378010 244080
rect 377954 237088 378010 237144
rect 377954 236136 378010 236192
rect 378046 228248 378102 228304
rect 378046 227704 378102 227760
rect 378874 272040 378930 272096
rect 379242 272040 379298 272096
rect 379242 267144 379298 267200
rect 410522 353368 410578 353424
rect 421010 395392 421066 395448
rect 434810 387640 434866 387696
rect 379610 299240 379666 299296
rect 440330 291080 440386 291136
rect 440422 288768 440478 288824
rect 379518 275984 379574 276040
rect 440330 275984 440386 276040
rect 379426 273944 379482 274000
rect 379334 261160 379390 261216
rect 440238 259120 440294 259176
rect 379702 242256 379758 242312
rect 381634 240624 381690 240680
rect 382278 240216 382334 240272
rect 383014 236000 383070 236056
rect 389822 237904 389878 237960
rect 390190 136584 390246 136640
rect 396722 119040 396778 119096
rect 398746 179968 398802 180024
rect 398102 174528 398158 174584
rect 397458 145560 397514 145616
rect 397458 144236 397460 144256
rect 397460 144236 397512 144256
rect 397512 144236 397514 144256
rect 397458 144200 397514 144236
rect 397550 143656 397606 143712
rect 397550 142180 397606 142216
rect 397550 142160 397552 142180
rect 397552 142160 397604 142180
rect 397604 142160 397606 142180
rect 397458 141616 397514 141672
rect 397366 140256 397422 140312
rect 397458 138896 397514 138952
rect 397458 137536 397514 137592
rect 397550 136856 397606 136912
rect 397458 135360 397514 135416
rect 397458 134700 397514 134736
rect 397458 134680 397460 134700
rect 397460 134680 397512 134700
rect 397512 134680 397514 134700
rect 397458 133320 397514 133376
rect 397550 132640 397606 132696
rect 397550 130600 397606 130656
rect 397458 129920 397514 129976
rect 398194 129920 398250 129976
rect 397458 128696 397514 128752
rect 397458 127880 397514 127936
rect 397458 126656 397514 126712
rect 397550 125976 397606 126032
rect 397458 125296 397514 125352
rect 397458 123800 397514 123856
rect 398194 123120 398250 123176
rect 397458 121896 397514 121952
rect 397458 121216 397514 121272
rect 397458 119856 397514 119912
rect 397458 117136 397514 117192
rect 397458 115096 397514 115152
rect 397458 114452 397460 114472
rect 397460 114452 397512 114472
rect 397512 114452 397514 114472
rect 397458 114416 397514 114452
rect 397458 113092 397460 113112
rect 397460 113092 397512 113112
rect 397512 113092 397514 113112
rect 397458 113056 397514 113092
rect 397458 111016 397514 111072
rect 397458 110372 397460 110392
rect 397460 110372 397512 110392
rect 397512 110372 397514 110392
rect 397458 110336 397514 110372
rect 397458 108160 397514 108216
rect 397458 105596 397514 105632
rect 397734 109520 397790 109576
rect 397642 106256 397698 106312
rect 397458 105576 397460 105596
rect 397460 105576 397512 105596
rect 397512 105576 397514 105596
rect 396906 96600 396962 96656
rect 398010 104080 398066 104136
rect 397550 103536 397606 103592
rect 397550 102856 397606 102912
rect 397550 101496 397606 101552
rect 397642 100816 397698 100872
rect 397550 99456 397606 99512
rect 397550 97280 397606 97336
rect 398746 132096 398802 132152
rect 398654 127880 398710 127936
rect 398286 117816 398342 117872
rect 398930 116456 398986 116512
rect 399114 98776 399170 98832
rect 414294 226888 414350 226944
rect 417422 238312 417478 238368
rect 422206 146920 422262 146976
rect 427910 238720 427966 238776
rect 438858 239400 438914 239456
rect 439502 147736 439558 147792
rect 439962 147736 440018 147792
rect 440974 287000 441030 287056
rect 441526 287036 441528 287056
rect 441528 287036 441580 287056
rect 441580 287036 441582 287056
rect 441526 287000 441582 287036
rect 440882 275984 440938 276040
rect 440514 257080 440570 257136
rect 442814 297064 442870 297120
rect 441710 295024 441766 295080
rect 442814 295024 442870 295080
rect 442170 284960 442226 285016
rect 442722 282104 442778 282160
rect 442814 280220 442870 280256
rect 442814 280200 442816 280220
rect 442816 280200 442868 280220
rect 442868 280200 442870 280220
rect 442630 278024 442686 278080
rect 442722 273944 442778 274000
rect 442814 272076 442816 272096
rect 442816 272076 442868 272096
rect 442868 272076 442870 272096
rect 442814 272040 442870 272076
rect 442262 269864 442318 269920
rect 442814 267144 442870 267200
rect 442354 265124 442410 265160
rect 442354 265104 442356 265124
rect 442356 265104 442408 265124
rect 442408 265104 442410 265124
rect 442722 263064 442778 263120
rect 441710 261160 441766 261216
rect 442814 261160 442870 261216
rect 441618 248104 441674 248160
rect 441618 247016 441674 247072
rect 441618 246200 441674 246256
rect 442906 252320 442962 252376
rect 442722 250280 442778 250336
rect 441802 247016 441858 247072
rect 442906 246200 442962 246256
rect 442170 244024 442226 244080
rect 442906 242156 442908 242176
rect 442908 242156 442960 242176
rect 442960 242156 442962 242176
rect 442906 242120 442962 242156
rect 443182 292984 443238 293040
rect 443090 255040 443146 255096
rect 443182 236972 443238 237008
rect 443182 236952 443184 236972
rect 443184 236952 443236 236972
rect 443236 236952 443238 236972
rect 446586 201456 446642 201512
rect 449254 145560 449310 145616
rect 449346 143384 449402 143440
rect 400126 139984 400182 140040
rect 399574 111832 399630 111888
rect 427726 91024 427782 91080
rect 430394 93744 430450 93800
rect 442998 95240 443054 95296
rect 443826 95240 443882 95296
rect 449530 143248 449586 143304
rect 449438 141480 449494 141536
rect 449438 130076 449494 130112
rect 449438 130056 449440 130076
rect 449440 130056 449492 130076
rect 449492 130056 449494 130076
rect 449990 137944 450046 138000
rect 451554 147736 451610 147792
rect 451462 142296 451518 142352
rect 451278 138896 451334 138952
rect 450542 136584 450598 136640
rect 450082 135496 450138 135552
rect 449990 131144 450046 131200
rect 449898 129104 449954 129160
rect 449346 117000 449402 117056
rect 449898 101904 449954 101960
rect 451554 125296 451610 125352
rect 451278 124616 451334 124672
rect 452566 144336 452622 144392
rect 452474 142840 452530 142896
rect 451922 140256 451978 140312
rect 452106 138216 452162 138272
rect 451922 134136 451978 134192
rect 452198 133456 452254 133512
rect 452566 130736 452622 130792
rect 452566 129376 452622 129432
rect 452106 127336 452162 127392
rect 452566 126656 452622 126712
rect 452566 125296 452622 125352
rect 451646 123936 451702 123992
rect 452566 122612 452568 122632
rect 452568 122612 452620 122632
rect 452620 122612 452622 122632
rect 452566 122576 452622 122612
rect 450082 120400 450138 120456
rect 452474 117816 452530 117872
rect 451554 115812 451556 115832
rect 451556 115812 451608 115832
rect 451608 115812 451610 115832
rect 451554 115776 451610 115812
rect 451370 114960 451426 115016
rect 451278 106256 451334 106312
rect 450174 104080 450230 104136
rect 452474 113736 452530 113792
rect 452566 111716 452622 111752
rect 452566 111696 452568 111716
rect 452568 111696 452620 111716
rect 452620 111696 452622 111716
rect 452474 111016 452530 111072
rect 452106 109656 452162 109712
rect 451554 108976 451610 109032
rect 451738 108160 451794 108216
rect 452566 106936 452622 106992
rect 452842 108976 452898 109032
rect 452566 104916 452622 104952
rect 452566 104896 452568 104916
rect 452568 104896 452620 104916
rect 452620 104896 452622 104916
rect 452566 102856 452622 102912
rect 452566 100136 452622 100192
rect 452290 98096 452346 98152
rect 452566 97416 452622 97472
rect 454130 224848 454186 224904
rect 453302 93744 453358 93800
rect 459558 149096 459614 149152
rect 485778 233280 485834 233336
rect 498842 396616 498898 396672
rect 508502 395392 508558 395448
rect 530674 357992 530730 358048
rect 533434 409536 533490 409592
rect 533434 400016 533490 400072
rect 535458 600344 535514 600400
rect 535458 574096 535514 574152
rect 535458 568656 535514 568712
rect 535458 563916 535514 563952
rect 535458 563896 535460 563916
rect 535460 563896 535512 563916
rect 535512 563896 535514 563916
rect 535458 556416 535514 556472
rect 535458 553696 535514 553752
rect 534354 550976 534410 551032
rect 534354 429936 534410 429992
rect 534262 407496 534318 407552
rect 535734 596264 535790 596320
rect 535642 594532 535644 594552
rect 535644 594532 535696 594552
rect 535696 594532 535698 594552
rect 535642 594496 535698 594532
rect 535642 591776 535698 591832
rect 535734 584296 535790 584352
rect 535734 581576 535790 581632
rect 535734 578856 535790 578912
rect 535734 576852 535736 576872
rect 535736 576852 535788 576872
rect 535788 576852 535790 576872
rect 535734 576816 535790 576852
rect 535642 571376 535698 571432
rect 535642 561176 535698 561232
rect 535550 536016 535606 536072
rect 535550 533296 535606 533352
rect 535550 528572 535552 528592
rect 535552 528572 535604 528592
rect 535604 528572 535606 528592
rect 535550 528536 535606 528572
rect 535550 521056 535606 521112
rect 535550 518336 535606 518392
rect 535550 515616 535606 515672
rect 535550 513576 535606 513632
rect 535550 508136 535606 508192
rect 535550 506096 535606 506152
rect 535550 503376 535606 503432
rect 535550 500656 535606 500712
rect 535550 495896 535606 495952
rect 535550 493176 535606 493232
rect 535550 485696 535606 485752
rect 535550 483012 535552 483032
rect 535552 483012 535604 483032
rect 535604 483012 535606 483032
rect 535550 482976 535606 483012
rect 535458 404776 535514 404832
rect 535826 523776 535882 523832
rect 536930 548936 536986 548992
rect 537022 546216 537078 546272
rect 537022 538736 537078 538792
rect 536746 510856 536802 510912
rect 535734 488416 535790 488472
rect 535734 478216 535790 478272
rect 535734 475496 535790 475552
rect 535734 472776 535790 472832
rect 535734 470736 535790 470792
rect 535734 468036 535790 468072
rect 535734 468016 535736 468036
rect 535736 468016 535788 468036
rect 535788 468016 535790 468036
rect 535734 465296 535790 465352
rect 535734 462576 535790 462632
rect 535734 460536 535790 460592
rect 535734 457816 535790 457872
rect 535734 453056 535790 453112
rect 535734 447616 535790 447672
rect 535734 444896 535790 444952
rect 535734 442856 535790 442912
rect 535734 435376 535790 435432
rect 535734 432656 535790 432712
rect 535826 427216 535882 427272
rect 535826 422456 535882 422512
rect 535826 419736 535882 419792
rect 535826 417696 535882 417752
rect 535826 414976 535882 415032
rect 535826 412256 535882 412312
rect 535826 402056 535882 402112
rect 536930 440136 536986 440192
rect 537022 327664 537078 327720
rect 538402 594768 538458 594824
rect 580170 697176 580226 697232
rect 545118 597760 545174 597816
rect 546498 398520 546554 398576
rect 547970 398656 548026 398712
rect 550730 399880 550786 399936
rect 550638 399744 550694 399800
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 579802 524456 579858 524512
rect 579618 511284 579674 511320
rect 579618 511264 579620 511284
rect 579620 511264 579672 511284
rect 579672 511264 579674 511284
rect 580262 484608 580318 484664
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 579710 404948 579712 404968
rect 579712 404948 579764 404968
rect 579764 404948 579766 404968
rect 579710 404912 579766 404948
rect 582470 471416 582526 471472
rect 580906 458088 580962 458144
rect 582378 458088 582434 458144
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580262 325216 580318 325272
rect 579986 312024 580042 312080
rect 579618 298696 579674 298752
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 582378 272176 582434 272232
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579986 205672 580042 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580354 139304 580410 139360
rect 580262 125976 580318 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 579894 33108 579950 33144
rect 579894 33088 579896 33108
rect 579896 33088 579948 33108
rect 579948 33088 579950 33108
rect 579894 19760 579950 19816
rect 580170 6568 580226 6624
<< obsm2 >>
rect 68800 95100 164756 174600
<< metal3 >>
rect 63350 702476 63356 702540
rect 63420 702538 63426 702540
rect 267641 702538 267707 702541
rect 63420 702536 267707 702538
rect 63420 702480 267646 702536
rect 267702 702480 267707 702536
rect 63420 702478 267707 702480
rect 63420 702476 63426 702478
rect 267641 702475 267707 702478
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect -960 671198 674 671258
rect -960 671122 480 671198
rect 614 671122 674 671198
rect -960 671108 674 671122
rect 246 671062 674 671108
rect 246 670714 306 671062
rect 243486 670714 243492 670716
rect 246 670654 243492 670714
rect 243486 670652 243492 670654
rect 243556 670652 243562 670716
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 336038 604420 336044 604484
rect 336108 604482 336114 604484
rect 515397 604482 515463 604485
rect 336108 604480 515463 604482
rect 336108 604424 515402 604480
rect 515458 604424 515463 604480
rect 336108 604422 515463 604424
rect 336108 604420 336114 604422
rect 515397 604419 515463 604422
rect 583520 604060 584960 604300
rect 340086 603196 340092 603260
rect 340156 603258 340162 603260
rect 419533 603258 419599 603261
rect 420177 603258 420243 603261
rect 340156 603256 420243 603258
rect 340156 603200 419538 603256
rect 419594 603200 420182 603256
rect 420238 603200 420243 603256
rect 340156 603198 420243 603200
rect 340156 603196 340162 603198
rect 419533 603195 419599 603198
rect 420177 603195 420243 603198
rect 337326 603060 337332 603124
rect 337396 603122 337402 603124
rect 507853 603122 507919 603125
rect 337396 603120 507919 603122
rect 337396 603064 507858 603120
rect 507914 603064 507919 603120
rect 337396 603062 507919 603064
rect 337396 603060 337402 603062
rect 507853 603059 507919 603062
rect 336089 601898 336155 601901
rect 433609 601898 433675 601901
rect 336089 601896 433675 601898
rect 336089 601840 336094 601896
rect 336150 601840 433614 601896
rect 433670 601840 433675 601896
rect 336089 601838 433675 601840
rect 336089 601835 336155 601838
rect 433609 601835 433675 601838
rect 331121 601762 331187 601765
rect 445845 601762 445911 601765
rect 331121 601760 445911 601762
rect 331121 601704 331126 601760
rect 331182 601704 445850 601760
rect 445906 601704 445911 601760
rect 331121 601702 445911 601704
rect 331121 601699 331187 601702
rect 445845 601699 445911 601702
rect 328361 600538 328427 600541
rect 462589 600538 462655 600541
rect 328361 600536 462655 600538
rect 328361 600480 328366 600536
rect 328422 600480 462594 600536
rect 462650 600480 462655 600536
rect 328361 600478 462655 600480
rect 328361 600475 328427 600478
rect 462589 600475 462655 600478
rect 335854 600340 335860 600404
rect 335924 600402 335930 600404
rect 535453 600402 535519 600405
rect 335924 600400 535519 600402
rect 335924 600344 535458 600400
rect 535514 600344 535519 600400
rect 335924 600342 535519 600344
rect 335924 600340 335930 600342
rect 535453 600339 535519 600342
rect 313917 599178 313983 599181
rect 429193 599178 429259 599181
rect 313917 599176 429259 599178
rect 313917 599120 313922 599176
rect 313978 599120 429198 599176
rect 429254 599120 429259 599176
rect 313917 599118 429259 599120
rect 313917 599115 313983 599118
rect 429193 599115 429259 599118
rect 338941 599042 339007 599045
rect 479333 599042 479399 599045
rect 338941 599040 479399 599042
rect 338941 598984 338946 599040
rect 339002 598984 479338 599040
rect 479394 598984 479399 599040
rect 338941 598982 479399 598984
rect 338941 598979 339007 598982
rect 479333 598979 479399 598982
rect 505737 599042 505803 599045
rect 539542 599042 539548 599044
rect 505737 599040 539548 599042
rect 505737 598984 505742 599040
rect 505798 598984 539548 599040
rect 505737 598982 539548 598984
rect 505737 598979 505803 598982
rect 539542 598980 539548 598982
rect 539612 598980 539618 599044
rect 317413 597954 317479 597957
rect 364793 597954 364859 597957
rect 317413 597952 364859 597954
rect 317413 597896 317418 597952
rect 317474 597896 364798 597952
rect 364854 597896 364859 597952
rect 317413 597894 364859 597896
rect 317413 597891 317479 597894
rect 364793 597891 364859 597894
rect 313774 597756 313780 597820
rect 313844 597818 313850 597820
rect 340321 597818 340387 597821
rect 313844 597816 340387 597818
rect 313844 597760 340326 597816
rect 340382 597760 340387 597816
rect 313844 597758 340387 597760
rect 313844 597756 313850 597758
rect 340321 597755 340387 597758
rect 340638 597756 340644 597820
rect 340708 597818 340714 597820
rect 467189 597818 467255 597821
rect 340708 597816 467255 597818
rect 340708 597760 467194 597816
rect 467250 597760 467255 597816
rect 340708 597758 467255 597760
rect 340708 597756 340714 597758
rect 467189 597755 467255 597758
rect 522941 597818 523007 597821
rect 545113 597818 545179 597821
rect 522941 597816 545179 597818
rect 522941 597760 522946 597816
rect 523002 597760 545118 597816
rect 545174 597760 545179 597816
rect 522941 597758 545179 597760
rect 522941 597755 523007 597758
rect 545113 597755 545179 597758
rect 335997 597682 336063 597685
rect 534022 597682 534028 597684
rect 335997 597680 534028 597682
rect 335997 597624 336002 597680
rect 336058 597624 534028 597680
rect 335997 597622 534028 597624
rect 335997 597619 336063 597622
rect 534022 597620 534028 597622
rect 534092 597620 534098 597684
rect 311014 596396 311020 596460
rect 311084 596458 311090 596460
rect 355133 596458 355199 596461
rect 311084 596456 355199 596458
rect 311084 596400 355138 596456
rect 355194 596400 355199 596456
rect 311084 596398 355199 596400
rect 311084 596396 311090 596398
rect 355133 596395 355199 596398
rect 338614 596260 338620 596324
rect 338684 596322 338690 596324
rect 535729 596322 535795 596325
rect 338684 596320 535795 596322
rect 338684 596264 535734 596320
rect 535790 596264 535795 596320
rect 338684 596262 535795 596264
rect 338684 596260 338690 596262
rect 535729 596259 535795 596262
rect 334617 595098 334683 595101
rect 359641 595098 359707 595101
rect 334617 595096 359707 595098
rect 334617 595040 334622 595096
rect 334678 595040 359646 595096
rect 359702 595040 359707 595096
rect 334617 595038 359707 595040
rect 334617 595035 334683 595038
rect 359641 595035 359707 595038
rect 293861 594962 293927 594965
rect 362217 594962 362283 594965
rect 293861 594960 362283 594962
rect 293861 594904 293866 594960
rect 293922 594904 362222 594960
rect 362278 594904 362283 594960
rect 293861 594902 362283 594904
rect 293861 594899 293927 594902
rect 362217 594899 362283 594902
rect 329097 594826 329163 594829
rect 538397 594826 538463 594829
rect 329097 594824 538463 594826
rect 329097 594768 329102 594824
rect 329158 594768 538402 594824
rect 538458 594768 538463 594824
rect 329097 594766 538463 594768
rect 329097 594763 329163 594766
rect 538397 594763 538463 594766
rect 336549 594554 336615 594557
rect 535637 594554 535703 594557
rect 336549 594552 340124 594554
rect 336549 594496 336554 594552
rect 336610 594496 340124 594552
rect 336549 594494 340124 594496
rect 533140 594552 535703 594554
rect 533140 594496 535642 594552
rect 535698 594496 535703 594552
rect 533140 594494 535703 594496
rect 336549 594491 336615 594494
rect 535637 594491 535703 594494
rect 55070 593404 55076 593468
rect 55140 593466 55146 593468
rect 118693 593466 118759 593469
rect 119337 593466 119403 593469
rect 55140 593464 119403 593466
rect 55140 593408 118698 593464
rect 118754 593408 119342 593464
rect 119398 593408 119403 593464
rect 55140 593406 119403 593408
rect 55140 593404 55146 593406
rect 118693 593403 118759 593406
rect 119337 593403 119403 593406
rect -960 592908 480 593148
rect 340638 592650 340644 592652
rect 190410 592590 340644 592650
rect 50838 592180 50844 592244
rect 50908 592242 50914 592244
rect 178585 592242 178651 592245
rect 50908 592240 178651 592242
rect 50908 592184 178590 592240
rect 178646 592184 178651 592240
rect 50908 592182 178651 592184
rect 50908 592180 50914 592182
rect 178585 592179 178651 592182
rect 59118 592044 59124 592108
rect 59188 592106 59194 592108
rect 188245 592106 188311 592109
rect 190410 592106 190470 592590
rect 340638 592588 340644 592590
rect 340708 592588 340714 592652
rect 59188 592104 190470 592106
rect 59188 592048 188250 592104
rect 188306 592048 190470 592104
rect 59188 592046 190470 592048
rect 59188 592044 59194 592046
rect 188245 592043 188311 592046
rect 337101 591834 337167 591837
rect 535637 591834 535703 591837
rect 337101 591832 340124 591834
rect 337101 591776 337106 591832
rect 337162 591776 340124 591832
rect 337101 591774 340124 591776
rect 533140 591832 535703 591834
rect 533140 591776 535642 591832
rect 535698 591776 535703 591832
rect 533140 591774 535703 591776
rect 337101 591771 337167 591774
rect 535637 591771 535703 591774
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 337653 589114 337719 589117
rect 535494 589114 535500 589116
rect 337653 589112 340124 589114
rect 337653 589056 337658 589112
rect 337714 589056 340124 589112
rect 337653 589054 340124 589056
rect 533140 589054 535500 589114
rect 337653 589051 337719 589054
rect 535494 589052 535500 589054
rect 535564 589052 535570 589116
rect 42701 588026 42767 588029
rect 156781 588026 156847 588029
rect 42701 588024 156847 588026
rect 42701 587968 42706 588024
rect 42762 587968 156786 588024
rect 156842 587968 156847 588024
rect 42701 587966 156847 587968
rect 42701 587963 42767 587966
rect 156781 587963 156847 587966
rect 60038 586740 60044 586804
rect 60108 586802 60114 586804
rect 115565 586802 115631 586805
rect 60108 586800 115631 586802
rect 60108 586744 115570 586800
rect 115626 586744 115631 586800
rect 60108 586742 115631 586744
rect 60108 586740 60114 586742
rect 115565 586739 115631 586742
rect 44817 586666 44883 586669
rect 80697 586666 80763 586669
rect 44817 586664 80763 586666
rect 44817 586608 44822 586664
rect 44878 586608 80702 586664
rect 80758 586608 80763 586664
rect 44817 586606 80763 586608
rect 44817 586603 44883 586606
rect 80697 586603 80763 586606
rect 220537 586666 220603 586669
rect 220721 586666 220787 586669
rect 245009 586666 245075 586669
rect 220537 586664 245075 586666
rect 220537 586608 220542 586664
rect 220598 586608 220726 586664
rect 220782 586608 245014 586664
rect 245070 586608 245075 586664
rect 220537 586606 245075 586608
rect 220537 586603 220603 586606
rect 220721 586603 220787 586606
rect 245009 586603 245075 586606
rect 210417 586394 210483 586397
rect 210877 586394 210943 586397
rect 271137 586394 271203 586397
rect 210417 586392 271203 586394
rect 210417 586336 210422 586392
rect 210478 586336 210882 586392
rect 210938 586336 271142 586392
rect 271198 586336 271203 586392
rect 210417 586334 271203 586336
rect 210417 586331 210483 586334
rect 210877 586331 210943 586334
rect 271137 586331 271203 586334
rect 337653 586394 337719 586397
rect 533654 586394 533660 586396
rect 337653 586392 340124 586394
rect 337653 586336 337658 586392
rect 337714 586336 340124 586392
rect 337653 586334 340124 586336
rect 533140 586334 533660 586394
rect 337653 586331 337719 586334
rect 533654 586332 533660 586334
rect 533724 586332 533730 586396
rect 43989 585306 44055 585309
rect 74349 585306 74415 585309
rect 43989 585304 74415 585306
rect 43989 585248 43994 585304
rect 44050 585248 74354 585304
rect 74410 585248 74415 585304
rect 43989 585246 74415 585248
rect 43989 585243 44055 585246
rect 74349 585243 74415 585246
rect 61377 585170 61443 585173
rect 134241 585170 134307 585173
rect 61377 585168 134307 585170
rect 61377 585112 61382 585168
rect 61438 585112 134246 585168
rect 134302 585112 134307 585168
rect 61377 585110 134307 585112
rect 61377 585107 61443 585110
rect 134241 585107 134307 585110
rect 175457 585170 175523 585173
rect 243670 585170 243676 585172
rect 175457 585168 243676 585170
rect 175457 585112 175462 585168
rect 175518 585112 243676 585168
rect 175457 585110 243676 585112
rect 175457 585107 175523 585110
rect 243670 585108 243676 585110
rect 243740 585108 243746 585172
rect 64638 584564 64644 584628
rect 64708 584626 64714 584628
rect 64781 584626 64847 584629
rect 64708 584624 64847 584626
rect 64708 584568 64786 584624
rect 64842 584568 64847 584624
rect 64708 584566 64847 584568
rect 64708 584564 64714 584566
rect 64781 584563 64847 584566
rect 337653 584354 337719 584357
rect 535729 584354 535795 584357
rect 337653 584352 340124 584354
rect 337653 584296 337658 584352
rect 337714 584296 340124 584352
rect 337653 584294 340124 584296
rect 533140 584352 535795 584354
rect 533140 584296 535734 584352
rect 535790 584296 535795 584352
rect 533140 584294 535795 584296
rect 337653 584291 337719 584294
rect 535729 584291 535795 584294
rect 58985 584082 59051 584085
rect 337510 584082 337516 584084
rect 58985 584080 337516 584082
rect 58985 584024 58990 584080
rect 59046 584024 337516 584080
rect 58985 584022 337516 584024
rect 58985 584019 59051 584022
rect 337510 584020 337516 584022
rect 337580 584020 337586 584084
rect 56501 583946 56567 583949
rect 322197 583946 322263 583949
rect 56501 583944 322263 583946
rect 56501 583888 56506 583944
rect 56562 583888 322202 583944
rect 322258 583888 322263 583944
rect 56501 583886 322263 583888
rect 56501 583883 56567 583886
rect 322197 583883 322263 583886
rect 245745 583266 245811 583269
rect 243892 583264 245811 583266
rect 243892 583208 245750 583264
rect 245806 583208 245811 583264
rect 243892 583206 245811 583208
rect 245745 583203 245811 583206
rect 320081 582994 320147 582997
rect 337326 582994 337332 582996
rect 320081 582992 337332 582994
rect 320081 582936 320086 582992
rect 320142 582936 337332 582992
rect 320081 582934 337332 582936
rect 320081 582931 320147 582934
rect 337326 582932 337332 582934
rect 337396 582932 337402 582996
rect 61878 582524 61884 582588
rect 61948 582586 61954 582588
rect 61948 582526 64124 582586
rect 61948 582524 61954 582526
rect 243486 582388 243492 582452
rect 243556 582450 243562 582452
rect 245694 582450 245700 582452
rect 243556 582390 245700 582450
rect 243556 582388 243562 582390
rect 245694 582388 245700 582390
rect 245764 582388 245770 582452
rect 337653 581634 337719 581637
rect 535729 581634 535795 581637
rect 337653 581632 340124 581634
rect 337653 581576 337658 581632
rect 337714 581576 340124 581632
rect 337653 581574 340124 581576
rect 533140 581632 535795 581634
rect 533140 581576 535734 581632
rect 535790 581576 535795 581632
rect 533140 581574 535795 581576
rect 337653 581571 337719 581574
rect 535729 581571 535795 581574
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 244181 579866 244247 579869
rect 243892 579864 244247 579866
rect 243892 579808 244186 579864
rect 244242 579808 244247 579864
rect 243892 579806 244247 579808
rect 244181 579803 244247 579806
rect 60641 579186 60707 579189
rect 63493 579186 63559 579189
rect 60641 579184 64124 579186
rect 60641 579128 60646 579184
rect 60702 579128 63498 579184
rect 63554 579128 64124 579184
rect 60641 579126 64124 579128
rect 60641 579123 60707 579126
rect 63493 579123 63559 579126
rect 337653 578914 337719 578917
rect 535729 578914 535795 578917
rect 337653 578912 340124 578914
rect 337653 578856 337658 578912
rect 337714 578856 340124 578912
rect 337653 578854 340124 578856
rect 533140 578912 535795 578914
rect 533140 578856 535734 578912
rect 535790 578856 535795 578912
rect 533140 578854 535795 578856
rect 337653 578851 337719 578854
rect 535729 578851 535795 578854
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 337653 576874 337719 576877
rect 535729 576874 535795 576877
rect 337653 576872 340124 576874
rect 337653 576816 337658 576872
rect 337714 576816 340124 576872
rect 337653 576814 340124 576816
rect 533140 576872 535795 576874
rect 533140 576816 535734 576872
rect 535790 576816 535795 576872
rect 533140 576814 535795 576816
rect 337653 576811 337719 576814
rect 535729 576811 535795 576814
rect 245653 576466 245719 576469
rect 243892 576464 245719 576466
rect 243892 576408 245658 576464
rect 245714 576408 245719 576464
rect 243892 576406 245719 576408
rect 245653 576403 245719 576406
rect 61561 575786 61627 575789
rect 61561 575784 64124 575786
rect 61561 575728 61566 575784
rect 61622 575728 64124 575784
rect 61561 575726 64124 575728
rect 61561 575723 61627 575726
rect 337837 574154 337903 574157
rect 535453 574154 535519 574157
rect 337837 574152 340124 574154
rect 337837 574096 337842 574152
rect 337898 574096 340124 574152
rect 337837 574094 340124 574096
rect 533140 574152 535519 574154
rect 533140 574096 535458 574152
rect 535514 574096 535519 574152
rect 533140 574094 535519 574096
rect 337837 574091 337903 574094
rect 535453 574091 535519 574094
rect 245653 573066 245719 573069
rect 243892 573064 245719 573066
rect 243892 573008 245658 573064
rect 245714 573008 245719 573064
rect 243892 573006 245719 573008
rect 245653 573003 245719 573006
rect 60733 572386 60799 572389
rect 60733 572384 64124 572386
rect 60733 572328 60738 572384
rect 60794 572328 64124 572384
rect 60733 572326 64124 572328
rect 60733 572323 60799 572326
rect 337653 571434 337719 571437
rect 535637 571434 535703 571437
rect 337653 571432 340124 571434
rect 337653 571376 337658 571432
rect 337714 571376 340124 571432
rect 337653 571374 340124 571376
rect 533140 571432 535703 571434
rect 533140 571376 535642 571432
rect 535698 571376 535703 571432
rect 533140 571374 535703 571376
rect 337653 571371 337719 571374
rect 535637 571371 535703 571374
rect 245653 569666 245719 569669
rect 243892 569664 245719 569666
rect 243892 569608 245658 569664
rect 245714 569608 245719 569664
rect 243892 569606 245719 569608
rect 245653 569603 245719 569606
rect 60733 568986 60799 568989
rect 60733 568984 64124 568986
rect 60733 568928 60738 568984
rect 60794 568928 64124 568984
rect 60733 568926 64124 568928
rect 60733 568923 60799 568926
rect 337653 568714 337719 568717
rect 535453 568714 535519 568717
rect 337653 568712 340124 568714
rect 337653 568656 337658 568712
rect 337714 568656 340124 568712
rect 337653 568654 340124 568656
rect 533140 568712 535519 568714
rect 533140 568656 535458 568712
rect 535514 568656 535519 568712
rect 533140 568654 535519 568656
rect 337653 568651 337719 568654
rect 535453 568651 535519 568654
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 534165 566674 534231 566677
rect 533140 566672 534231 566674
rect 245929 566266 245995 566269
rect 243892 566264 245995 566266
rect 243892 566208 245934 566264
rect 245990 566208 245995 566264
rect 243892 566206 245995 566208
rect 245929 566203 245995 566206
rect 333094 565796 333100 565860
rect 333164 565858 333170 565860
rect 340094 565858 340154 566644
rect 533140 566616 534170 566672
rect 534226 566616 534231 566672
rect 533140 566614 534231 566616
rect 534165 566611 534231 566614
rect 333164 565798 340154 565858
rect 333164 565796 333170 565798
rect 60733 565586 60799 565589
rect 60733 565584 64124 565586
rect 60733 565528 60738 565584
rect 60794 565528 64124 565584
rect 60733 565526 64124 565528
rect 60733 565523 60799 565526
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect 338757 563954 338823 563957
rect 535453 563954 535519 563957
rect 338757 563952 340124 563954
rect 338757 563896 338762 563952
rect 338818 563896 340124 563952
rect 338757 563894 340124 563896
rect 533140 563952 535519 563954
rect 533140 563896 535458 563952
rect 535514 563896 535519 563952
rect 533140 563894 535519 563896
rect 338757 563891 338823 563894
rect 535453 563891 535519 563894
rect 245561 562866 245627 562869
rect 243892 562864 245627 562866
rect 243892 562808 245566 562864
rect 245622 562808 245627 562864
rect 243892 562806 245627 562808
rect 245561 562803 245627 562806
rect 57830 562124 57836 562188
rect 57900 562186 57906 562188
rect 57900 562126 64124 562186
rect 57900 562124 57906 562126
rect 337653 561234 337719 561237
rect 535637 561234 535703 561237
rect 337653 561232 340124 561234
rect 337653 561176 337658 561232
rect 337714 561176 340124 561232
rect 337653 561174 340124 561176
rect 533140 561232 535703 561234
rect 533140 561176 535642 561232
rect 535698 561176 535703 561232
rect 533140 561174 535703 561176
rect 337653 561171 337719 561174
rect 535637 561171 535703 561174
rect 245929 560146 245995 560149
rect 243892 560144 245995 560146
rect 243892 560088 245934 560144
rect 245990 560088 245995 560144
rect 243892 560086 245995 560088
rect 245929 560083 245995 560086
rect 336917 559194 336983 559197
rect 538438 559194 538444 559196
rect 336917 559192 340124 559194
rect 336917 559136 336922 559192
rect 336978 559136 340124 559192
rect 336917 559134 340124 559136
rect 533140 559134 538444 559194
rect 336917 559131 336983 559134
rect 538438 559132 538444 559134
rect 538508 559132 538514 559196
rect 55622 558724 55628 558788
rect 55692 558786 55698 558788
rect 55692 558726 64124 558786
rect 55692 558724 55698 558726
rect 245009 558242 245075 558245
rect 295374 558242 295380 558244
rect 245009 558240 295380 558242
rect 245009 558184 245014 558240
rect 245070 558184 295380 558240
rect 245009 558182 295380 558184
rect 245009 558179 245075 558182
rect 295374 558180 295380 558182
rect 295444 558180 295450 558244
rect 243670 557364 243676 557428
rect 243740 557426 243746 557428
rect 248413 557426 248479 557429
rect 249701 557426 249767 557429
rect 243740 557424 249767 557426
rect 243740 557368 248418 557424
rect 248474 557368 249706 557424
rect 249762 557368 249767 557424
rect 243740 557366 249767 557368
rect 243740 557364 243746 557366
rect 248413 557363 248479 557366
rect 249701 557363 249767 557366
rect 245653 556746 245719 556749
rect 243892 556744 245719 556746
rect 243892 556688 245658 556744
rect 245714 556688 245719 556744
rect 243892 556686 245719 556688
rect 245653 556683 245719 556686
rect 337929 556474 337995 556477
rect 535453 556474 535519 556477
rect 337929 556472 340124 556474
rect 337929 556416 337934 556472
rect 337990 556416 340124 556472
rect 337929 556414 340124 556416
rect 533140 556472 535519 556474
rect 533140 556416 535458 556472
rect 535514 556416 535519 556472
rect 533140 556414 535519 556416
rect 337929 556411 337995 556414
rect 535453 556411 535519 556414
rect 60733 555386 60799 555389
rect 60733 555384 64124 555386
rect 60733 555328 60738 555384
rect 60794 555328 64124 555384
rect 60733 555326 64124 555328
rect 60733 555323 60799 555326
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 337377 553754 337443 553757
rect 535453 553754 535519 553757
rect 337377 553752 340124 553754
rect 337377 553696 337382 553752
rect 337438 553696 340124 553752
rect 337377 553694 340124 553696
rect 533140 553752 535519 553754
rect 533140 553696 535458 553752
rect 535514 553696 535519 553752
rect 533140 553694 535519 553696
rect 337377 553691 337443 553694
rect 535453 553691 535519 553694
rect 245929 553346 245995 553349
rect 243892 553344 245995 553346
rect 243892 553288 245934 553344
rect 245990 553288 245995 553344
rect 243892 553286 245995 553288
rect 245929 553283 245995 553286
rect 60733 552666 60799 552669
rect 60733 552664 64124 552666
rect 60733 552608 60738 552664
rect 60794 552608 64124 552664
rect 60733 552606 64124 552608
rect 60733 552603 60799 552606
rect 337377 551034 337443 551037
rect 534349 551034 534415 551037
rect 337377 551032 340124 551034
rect 337377 550976 337382 551032
rect 337438 550976 340124 551032
rect 337377 550974 340124 550976
rect 533140 551032 534415 551034
rect 533140 550976 534354 551032
rect 534410 550976 534415 551032
rect 583520 551020 584960 551260
rect 533140 550974 534415 550976
rect 337377 550971 337443 550974
rect 534349 550971 534415 550974
rect 245929 549946 245995 549949
rect 243892 549944 245995 549946
rect 243892 549888 245934 549944
rect 245990 549888 245995 549944
rect 243892 549886 245995 549888
rect 245929 549883 245995 549886
rect 60733 549266 60799 549269
rect 60733 549264 64124 549266
rect 60733 549208 60738 549264
rect 60794 549208 64124 549264
rect 60733 549206 64124 549208
rect 60733 549203 60799 549206
rect 337653 548994 337719 548997
rect 536925 548994 536991 548997
rect 337653 548992 340124 548994
rect 337653 548936 337658 548992
rect 337714 548936 340124 548992
rect 337653 548934 340124 548936
rect 533140 548992 536991 548994
rect 533140 548936 536930 548992
rect 536986 548936 536991 548992
rect 533140 548934 536991 548936
rect 337653 548931 337719 548934
rect 536925 548931 536991 548934
rect 245929 546546 245995 546549
rect 243892 546544 245995 546546
rect 243892 546488 245934 546544
rect 245990 546488 245995 546544
rect 243892 546486 245995 546488
rect 245929 546483 245995 546486
rect 331806 546484 331812 546548
rect 331876 546546 331882 546548
rect 337377 546546 337443 546549
rect 331876 546544 337443 546546
rect 331876 546488 337382 546544
rect 337438 546488 337443 546544
rect 331876 546486 337443 546488
rect 331876 546484 331882 546486
rect 337377 546483 337443 546486
rect 337377 546274 337443 546277
rect 537017 546274 537083 546277
rect 337377 546272 340124 546274
rect 337377 546216 337382 546272
rect 337438 546216 340124 546272
rect 337377 546214 340124 546216
rect 533140 546272 537083 546274
rect 533140 546216 537022 546272
rect 537078 546216 537083 546272
rect 533140 546214 537083 546216
rect 337377 546211 337443 546214
rect 537017 546211 537083 546214
rect 60733 545866 60799 545869
rect 60733 545864 64124 545866
rect 60733 545808 60738 545864
rect 60794 545808 64124 545864
rect 60733 545806 64124 545808
rect 60733 545803 60799 545806
rect 337653 543554 337719 543557
rect 534390 543554 534396 543556
rect 337653 543552 340124 543554
rect 337653 543496 337658 543552
rect 337714 543496 340124 543552
rect 337653 543494 340124 543496
rect 533140 543494 534396 543554
rect 337653 543491 337719 543494
rect 534390 543492 534396 543494
rect 534460 543492 534466 543556
rect 244273 543146 244339 543149
rect 245285 543146 245351 543149
rect 243892 543144 245351 543146
rect 243892 543088 244278 543144
rect 244334 543088 245290 543144
rect 245346 543088 245351 543144
rect 243892 543086 245351 543088
rect 244273 543083 244339 543086
rect 245285 543083 245351 543086
rect 60733 542466 60799 542469
rect 60733 542464 64124 542466
rect 60733 542408 60738 542464
rect 60794 542408 64124 542464
rect 60733 542406 64124 542408
rect 60733 542403 60799 542406
rect 337469 541514 337535 541517
rect 534022 541514 534028 541516
rect 337469 541512 340124 541514
rect 337469 541456 337474 541512
rect 337530 541456 340124 541512
rect 337469 541454 340124 541456
rect 533140 541454 534028 541514
rect 337469 541451 337535 541454
rect 534022 541452 534028 541454
rect 534092 541452 534098 541516
rect -960 540684 480 540924
rect 246941 540290 247007 540293
rect 338614 540290 338620 540292
rect 243862 540288 338620 540290
rect 243862 540232 246946 540288
rect 247002 540232 338620 540288
rect 243862 540230 338620 540232
rect 243862 539716 243922 540230
rect 246941 540227 247007 540230
rect 338614 540228 338620 540230
rect 338684 540228 338690 540292
rect 60733 539066 60799 539069
rect 60733 539064 64124 539066
rect 60733 539008 60738 539064
rect 60794 539008 64124 539064
rect 60733 539006 64124 539008
rect 60733 539003 60799 539006
rect 337653 538794 337719 538797
rect 537017 538794 537083 538797
rect 337653 538792 340124 538794
rect 337653 538736 337658 538792
rect 337714 538736 340124 538792
rect 337653 538734 340124 538736
rect 533140 538792 537083 538794
rect 533140 538736 537022 538792
rect 537078 538736 537083 538792
rect 533140 538734 537083 538736
rect 337653 538731 337719 538734
rect 537017 538731 537083 538734
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 245837 536346 245903 536349
rect 243892 536344 245903 536346
rect 243892 536288 245842 536344
rect 245898 536288 245903 536344
rect 243892 536286 245903 536288
rect 245837 536283 245903 536286
rect 337285 536074 337351 536077
rect 535545 536074 535611 536077
rect 337285 536072 340124 536074
rect 337285 536016 337290 536072
rect 337346 536016 340124 536072
rect 337285 536014 340124 536016
rect 533140 536072 535611 536074
rect 533140 536016 535550 536072
rect 535606 536016 535611 536072
rect 533140 536014 535611 536016
rect 337285 536011 337351 536014
rect 535545 536011 535611 536014
rect 61561 535666 61627 535669
rect 61561 535664 64124 535666
rect 61561 535608 61566 535664
rect 61622 535608 64124 535664
rect 61561 535606 64124 535608
rect 61561 535603 61627 535606
rect 337653 533354 337719 533357
rect 535545 533354 535611 533357
rect 337653 533352 340124 533354
rect 337653 533296 337658 533352
rect 337714 533296 340124 533352
rect 337653 533294 340124 533296
rect 533140 533352 535611 533354
rect 533140 533296 535550 533352
rect 535606 533296 535611 533352
rect 533140 533294 535611 533296
rect 337653 533291 337719 533294
rect 535545 533291 535611 533294
rect 244181 532946 244247 532949
rect 243892 532944 244247 532946
rect 243892 532888 244186 532944
rect 244242 532888 244247 532944
rect 243892 532886 244247 532888
rect 244181 532883 244247 532886
rect 60733 532266 60799 532269
rect 60733 532264 64124 532266
rect 60733 532208 60738 532264
rect 60794 532208 64124 532264
rect 60733 532206 64124 532208
rect 60733 532203 60799 532206
rect 336825 531314 336891 531317
rect 534073 531314 534139 531317
rect 336825 531312 340124 531314
rect 336825 531256 336830 531312
rect 336886 531256 340124 531312
rect 336825 531254 340124 531256
rect 533140 531312 534139 531314
rect 533140 531256 534078 531312
rect 534134 531256 534139 531312
rect 533140 531254 534139 531256
rect 336825 531251 336891 531254
rect 534073 531251 534139 531254
rect 246849 529546 246915 529549
rect 243892 529544 246915 529546
rect 243892 529488 246854 529544
rect 246910 529488 246915 529544
rect 243892 529486 246915 529488
rect 246849 529483 246915 529486
rect 60733 528866 60799 528869
rect 60733 528864 64124 528866
rect 60733 528808 60738 528864
rect 60794 528808 64124 528864
rect 60733 528806 64124 528808
rect 60733 528803 60799 528806
rect 337326 528532 337332 528596
rect 337396 528594 337402 528596
rect 535545 528594 535611 528597
rect 337396 528534 340124 528594
rect 533140 528592 535611 528594
rect 533140 528536 535550 528592
rect 535606 528536 535611 528592
rect 533140 528534 535611 528536
rect 337396 528532 337402 528534
rect 535545 528531 535611 528534
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 245837 526146 245903 526149
rect 243892 526144 245903 526146
rect 243892 526088 245842 526144
rect 245898 526088 245903 526144
rect 243892 526086 245903 526088
rect 245837 526083 245903 526086
rect 337837 525874 337903 525877
rect 536782 525874 536788 525876
rect 337837 525872 340124 525874
rect 337837 525816 337842 525872
rect 337898 525816 340124 525872
rect 337837 525814 340124 525816
rect 533140 525814 536788 525874
rect 337837 525811 337903 525814
rect 536782 525812 536788 525814
rect 536852 525812 536858 525876
rect 60733 525466 60799 525469
rect 60733 525464 64124 525466
rect 60733 525408 60738 525464
rect 60794 525408 64124 525464
rect 60733 525406 64124 525408
rect 60733 525403 60799 525406
rect 245837 525058 245903 525061
rect 292614 525058 292620 525060
rect 245837 525056 292620 525058
rect 245837 525000 245842 525056
rect 245898 525000 292620 525056
rect 245837 524998 292620 525000
rect 245837 524995 245903 524998
rect 292614 524996 292620 524998
rect 292684 524996 292690 525060
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect 337469 523834 337535 523837
rect 535821 523834 535887 523837
rect 337469 523832 340124 523834
rect 337469 523776 337474 523832
rect 337530 523776 340124 523832
rect 337469 523774 340124 523776
rect 533140 523832 535887 523834
rect 533140 523776 535826 523832
rect 535882 523776 535887 523832
rect 533140 523774 535887 523776
rect 337469 523771 337535 523774
rect 535821 523771 535887 523774
rect 245837 522746 245903 522749
rect 243892 522744 245903 522746
rect 243892 522688 245842 522744
rect 245898 522688 245903 522744
rect 243892 522686 245903 522688
rect 245837 522683 245903 522686
rect 303521 522338 303587 522341
rect 336038 522338 336044 522340
rect 303521 522336 336044 522338
rect 303521 522280 303526 522336
rect 303582 522280 336044 522336
rect 303521 522278 336044 522280
rect 303521 522275 303587 522278
rect 336038 522276 336044 522278
rect 336108 522276 336114 522340
rect 57646 522004 57652 522068
rect 57716 522066 57722 522068
rect 57716 522006 64124 522066
rect 57716 522004 57722 522006
rect 337469 521114 337535 521117
rect 535545 521114 535611 521117
rect 337469 521112 340124 521114
rect 337469 521056 337474 521112
rect 337530 521056 340124 521112
rect 337469 521054 340124 521056
rect 533140 521112 535611 521114
rect 533140 521056 535550 521112
rect 535606 521056 535611 521112
rect 533140 521054 535611 521056
rect 337469 521051 337535 521054
rect 535545 521051 535611 521054
rect 245837 519346 245903 519349
rect 243892 519344 245903 519346
rect 243892 519288 245842 519344
rect 245898 519288 245903 519344
rect 243892 519286 245903 519288
rect 245837 519283 245903 519286
rect 58934 518604 58940 518668
rect 59004 518666 59010 518668
rect 59004 518606 64124 518666
rect 59004 518604 59010 518606
rect 535545 518394 535611 518397
rect 533140 518392 535611 518394
rect 301446 517516 301452 517580
rect 301516 517578 301522 517580
rect 340094 517578 340154 518364
rect 533140 518336 535550 518392
rect 535606 518336 535611 518392
rect 533140 518334 535611 518336
rect 535545 518331 535611 518334
rect 301516 517518 340154 517578
rect 301516 517516 301522 517518
rect 245694 515946 245700 515948
rect 243892 515886 245700 515946
rect 245694 515884 245700 515886
rect 245764 515946 245770 515948
rect 245837 515946 245903 515949
rect 245764 515944 245903 515946
rect 245764 515888 245842 515944
rect 245898 515888 245903 515944
rect 245764 515886 245903 515888
rect 245764 515884 245770 515886
rect 245837 515883 245903 515886
rect 337653 515674 337719 515677
rect 535545 515674 535611 515677
rect 337653 515672 340124 515674
rect 337653 515616 337658 515672
rect 337714 515616 340124 515672
rect 337653 515614 340124 515616
rect 533140 515672 535611 515674
rect 533140 515616 535550 515672
rect 535606 515616 535611 515672
rect 533140 515614 535611 515616
rect 337653 515611 337719 515614
rect 535545 515611 535611 515614
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 46606 514796 46612 514860
rect 46676 514858 46682 514860
rect 64094 514858 64154 515236
rect 46676 514798 64154 514858
rect 46676 514796 46682 514798
rect 337653 513634 337719 513637
rect 535545 513634 535611 513637
rect 337653 513632 340124 513634
rect 337653 513576 337658 513632
rect 337714 513576 340124 513632
rect 337653 513574 340124 513576
rect 533140 513632 535611 513634
rect 533140 513576 535550 513632
rect 535606 513576 535611 513632
rect 533140 513574 535611 513576
rect 337653 513571 337719 513574
rect 535545 513571 535611 513574
rect 245653 512546 245719 512549
rect 243892 512544 245719 512546
rect 243892 512488 245658 512544
rect 245714 512488 245719 512544
rect 243892 512486 245719 512488
rect 245653 512483 245719 512486
rect 60457 511866 60523 511869
rect 60457 511864 64124 511866
rect 60457 511808 60462 511864
rect 60518 511808 64124 511864
rect 60457 511806 64124 511808
rect 60457 511803 60523 511806
rect 579613 511322 579679 511325
rect 583520 511322 584960 511412
rect 579613 511320 584960 511322
rect 579613 511264 579618 511320
rect 579674 511264 584960 511320
rect 579613 511262 584960 511264
rect 579613 511259 579679 511262
rect 583520 511172 584960 511262
rect 337653 510914 337719 510917
rect 536741 510914 536807 510917
rect 337653 510912 340124 510914
rect 337653 510856 337658 510912
rect 337714 510856 340124 510912
rect 337653 510854 340124 510856
rect 533140 510912 536807 510914
rect 533140 510856 536746 510912
rect 536802 510856 536807 510912
rect 533140 510854 536807 510856
rect 337653 510851 337719 510854
rect 536741 510851 536807 510854
rect 245837 509826 245903 509829
rect 243892 509824 245903 509826
rect 243892 509768 245842 509824
rect 245898 509768 245903 509824
rect 243892 509766 245903 509768
rect 245837 509763 245903 509766
rect 61469 508466 61535 508469
rect 61469 508464 64124 508466
rect 61469 508408 61474 508464
rect 61530 508408 64124 508464
rect 61469 508406 64124 508408
rect 61469 508403 61535 508406
rect 337510 508132 337516 508196
rect 337580 508194 337586 508196
rect 535545 508194 535611 508197
rect 337580 508134 340124 508194
rect 533140 508192 535611 508194
rect 533140 508136 535550 508192
rect 535606 508136 535611 508192
rect 533140 508134 535611 508136
rect 337580 508132 337586 508134
rect 535545 508131 535611 508134
rect 245837 506426 245903 506429
rect 243892 506424 245903 506426
rect 243892 506368 245842 506424
rect 245898 506368 245903 506424
rect 243892 506366 245903 506368
rect 245837 506363 245903 506366
rect 337101 506154 337167 506157
rect 535545 506154 535611 506157
rect 337101 506152 340124 506154
rect 337101 506096 337106 506152
rect 337162 506096 340124 506152
rect 337101 506094 340124 506096
rect 533140 506152 535611 506154
rect 533140 506096 535550 506152
rect 535606 506096 535611 506152
rect 533140 506094 535611 506096
rect 337101 506091 337167 506094
rect 535545 506091 535611 506094
rect 62297 505066 62363 505069
rect 63125 505066 63191 505069
rect 62297 505064 64124 505066
rect 62297 505008 62302 505064
rect 62358 505008 63130 505064
rect 63186 505008 64124 505064
rect 62297 505006 64124 505008
rect 62297 505003 62363 505006
rect 63125 505003 63191 505006
rect 337653 503434 337719 503437
rect 535545 503434 535611 503437
rect 337653 503432 340124 503434
rect 337653 503376 337658 503432
rect 337714 503376 340124 503432
rect 337653 503374 340124 503376
rect 533140 503432 535611 503434
rect 533140 503376 535550 503432
rect 535606 503376 535611 503432
rect 533140 503374 535611 503376
rect 337653 503371 337719 503374
rect 535545 503371 535611 503374
rect 246941 503026 247007 503029
rect 335854 503026 335860 503028
rect 243892 503024 335860 503026
rect 243892 502968 246946 503024
rect 247002 502968 335860 503024
rect 243892 502966 335860 502968
rect 246941 502963 247007 502966
rect 335854 502964 335860 502966
rect 335924 502964 335930 503028
rect 62021 502346 62087 502349
rect 62021 502344 64124 502346
rect 62021 502288 62026 502344
rect 62082 502288 64124 502344
rect 62021 502286 64124 502288
rect 62021 502283 62087 502286
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 337745 500714 337811 500717
rect 535545 500714 535611 500717
rect 337745 500712 340124 500714
rect 337745 500656 337750 500712
rect 337806 500656 340124 500712
rect 337745 500654 340124 500656
rect 533140 500712 535611 500714
rect 533140 500656 535550 500712
rect 535606 500656 535611 500712
rect 533140 500654 535611 500656
rect 337745 500651 337811 500654
rect 535545 500651 535611 500654
rect 245837 499626 245903 499629
rect 243892 499624 245903 499626
rect 243892 499568 245842 499624
rect 245898 499568 245903 499624
rect 243892 499566 245903 499568
rect 245837 499563 245903 499566
rect 61929 498946 61995 498949
rect 61929 498944 64124 498946
rect 61929 498888 61934 498944
rect 61990 498888 64124 498944
rect 61929 498886 64124 498888
rect 61929 498883 61995 498886
rect 337653 497994 337719 497997
rect 535678 497994 535684 497996
rect 337653 497992 340124 497994
rect 337653 497936 337658 497992
rect 337714 497936 340124 497992
rect 337653 497934 340124 497936
rect 533140 497934 535684 497994
rect 337653 497931 337719 497934
rect 535678 497932 535684 497934
rect 535748 497932 535754 497996
rect 583520 497844 584960 498084
rect 245837 496226 245903 496229
rect 243892 496224 245903 496226
rect 243892 496168 245842 496224
rect 245898 496168 245903 496224
rect 243892 496166 245903 496168
rect 245837 496163 245903 496166
rect 337469 495954 337535 495957
rect 535545 495954 535611 495957
rect 337469 495952 340124 495954
rect 337469 495896 337474 495952
rect 337530 495896 340124 495952
rect 337469 495894 340124 495896
rect 533140 495952 535611 495954
rect 533140 495896 535550 495952
rect 535606 495896 535611 495952
rect 533140 495894 535611 495896
rect 337469 495891 337535 495894
rect 535545 495891 535611 495894
rect 62757 495546 62823 495549
rect 62757 495544 64124 495546
rect 62757 495488 62762 495544
rect 62818 495488 64124 495544
rect 62757 495486 64124 495488
rect 62757 495483 62823 495486
rect 337469 493234 337535 493237
rect 535545 493234 535611 493237
rect 337469 493232 340124 493234
rect 337469 493176 337474 493232
rect 337530 493176 340124 493232
rect 337469 493174 340124 493176
rect 533140 493232 535611 493234
rect 533140 493176 535550 493232
rect 535606 493176 535611 493232
rect 533140 493174 535611 493176
rect 337469 493171 337535 493174
rect 535545 493171 535611 493174
rect 245009 492826 245075 492829
rect 243892 492824 245075 492826
rect 243892 492768 245014 492824
rect 245070 492768 245075 492824
rect 243892 492766 245075 492768
rect 245009 492763 245075 492766
rect 60733 492146 60799 492149
rect 60733 492144 64124 492146
rect 60733 492088 60738 492144
rect 60794 492088 64124 492144
rect 60733 492086 64124 492088
rect 60733 492083 60799 492086
rect 337653 490514 337719 490517
rect 534073 490514 534139 490517
rect 337653 490512 340124 490514
rect 337653 490456 337658 490512
rect 337714 490456 340124 490512
rect 337653 490454 340124 490456
rect 533140 490512 534139 490514
rect 533140 490456 534078 490512
rect 534134 490456 534139 490512
rect 533140 490454 534139 490456
rect 337653 490451 337719 490454
rect 534073 490451 534139 490454
rect 246246 489426 246252 489428
rect 243892 489366 246252 489426
rect 246246 489364 246252 489366
rect 246316 489364 246322 489428
rect -960 488596 480 488836
rect 60733 488746 60799 488749
rect 60733 488744 64124 488746
rect 60733 488688 60738 488744
rect 60794 488688 64124 488744
rect 60733 488686 64124 488688
rect 60733 488683 60799 488686
rect 339309 488474 339375 488477
rect 535729 488474 535795 488477
rect 339309 488472 340124 488474
rect 339309 488416 339314 488472
rect 339370 488416 340124 488472
rect 339309 488414 340124 488416
rect 533140 488472 535795 488474
rect 533140 488416 535734 488472
rect 535790 488416 535795 488472
rect 533140 488414 535795 488416
rect 339309 488411 339375 488414
rect 535729 488411 535795 488414
rect 245837 486026 245903 486029
rect 243892 486024 245903 486026
rect 243892 485968 245842 486024
rect 245898 485968 245903 486024
rect 243892 485966 245903 485968
rect 245837 485963 245903 485966
rect 337745 485754 337811 485757
rect 535545 485754 535611 485757
rect 337745 485752 340124 485754
rect 337745 485696 337750 485752
rect 337806 485696 340124 485752
rect 337745 485694 340124 485696
rect 533140 485752 535611 485754
rect 533140 485696 535550 485752
rect 535606 485696 535611 485752
rect 533140 485694 535611 485696
rect 337745 485691 337811 485694
rect 535545 485691 535611 485694
rect 60733 485346 60799 485349
rect 60733 485344 64124 485346
rect 60733 485288 60738 485344
rect 60794 485288 64124 485344
rect 60733 485286 64124 485288
rect 60733 485283 60799 485286
rect 580257 484666 580323 484669
rect 583520 484666 584960 484756
rect 580257 484664 584960 484666
rect 580257 484608 580262 484664
rect 580318 484608 584960 484664
rect 580257 484606 584960 484608
rect 580257 484603 580323 484606
rect 583520 484516 584960 484606
rect 337929 483034 337995 483037
rect 338982 483034 338988 483036
rect 337929 483032 338988 483034
rect 337929 482976 337934 483032
rect 337990 482976 338988 483032
rect 337929 482974 338988 482976
rect 337929 482971 337995 482974
rect 338982 482972 338988 482974
rect 339052 483034 339058 483036
rect 535545 483034 535611 483037
rect 339052 482974 340124 483034
rect 533140 483032 535611 483034
rect 533140 482976 535550 483032
rect 535606 482976 535611 483032
rect 533140 482974 535611 482976
rect 339052 482972 339058 482974
rect 535545 482971 535611 482974
rect 245745 482626 245811 482629
rect 243892 482624 245811 482626
rect 243892 482568 245750 482624
rect 245806 482568 245811 482624
rect 243892 482566 245811 482568
rect 245745 482563 245811 482566
rect 60733 481946 60799 481949
rect 60733 481944 64124 481946
rect 60733 481888 60738 481944
rect 60794 481888 64124 481944
rect 60733 481886 64124 481888
rect 60733 481883 60799 481886
rect 336733 480314 336799 480317
rect 538254 480314 538260 480316
rect 336733 480312 340124 480314
rect 336733 480256 336738 480312
rect 336794 480256 340124 480312
rect 336733 480254 340124 480256
rect 533140 480254 538260 480314
rect 336733 480251 336799 480254
rect 538254 480252 538260 480254
rect 538324 480252 538330 480316
rect 243310 478956 243370 479196
rect 243302 478892 243308 478956
rect 243372 478892 243378 478956
rect 60733 478546 60799 478549
rect 60733 478544 64124 478546
rect 60733 478488 60738 478544
rect 60794 478488 64124 478544
rect 60733 478486 64124 478488
rect 60733 478483 60799 478486
rect 337745 478274 337811 478277
rect 535729 478274 535795 478277
rect 337745 478272 340124 478274
rect 337745 478216 337750 478272
rect 337806 478216 340124 478272
rect 337745 478214 340124 478216
rect 533140 478272 535795 478274
rect 533140 478216 535734 478272
rect 535790 478216 535795 478272
rect 533140 478214 535795 478216
rect 337745 478211 337811 478214
rect 535729 478211 535795 478214
rect 245745 475826 245811 475829
rect 243892 475824 245811 475826
rect -960 475690 480 475780
rect 243892 475768 245750 475824
rect 245806 475768 245811 475824
rect 243892 475766 245811 475768
rect 245745 475763 245811 475766
rect 3877 475690 3943 475693
rect -960 475688 3943 475690
rect -960 475632 3882 475688
rect 3938 475632 3943 475688
rect -960 475630 3943 475632
rect -960 475540 480 475630
rect 3877 475627 3943 475630
rect 337653 475554 337719 475557
rect 535729 475554 535795 475557
rect 337653 475552 340124 475554
rect 337653 475496 337658 475552
rect 337714 475496 340124 475552
rect 337653 475494 340124 475496
rect 533140 475552 535795 475554
rect 533140 475496 535734 475552
rect 535790 475496 535795 475552
rect 533140 475494 535795 475496
rect 337653 475491 337719 475494
rect 535729 475491 535795 475494
rect 63166 475084 63172 475148
rect 63236 475146 63242 475148
rect 63236 475086 64124 475146
rect 63236 475084 63242 475086
rect 336825 472834 336891 472837
rect 535729 472834 535795 472837
rect 336825 472832 340124 472834
rect 336825 472776 336830 472832
rect 336886 472776 340124 472832
rect 336825 472774 340124 472776
rect 533140 472832 535795 472834
rect 533140 472776 535734 472832
rect 535790 472776 535795 472832
rect 533140 472774 535795 472776
rect 336825 472771 336891 472774
rect 535729 472771 535795 472774
rect 245837 472426 245903 472429
rect 243892 472424 245903 472426
rect 243892 472368 245842 472424
rect 245898 472368 245903 472424
rect 243892 472366 245903 472368
rect 245837 472363 245903 472366
rect 63401 471746 63467 471749
rect 63401 471744 64124 471746
rect 63401 471688 63406 471744
rect 63462 471688 64124 471744
rect 63401 471686 64124 471688
rect 63401 471683 63467 471686
rect 582465 471474 582531 471477
rect 583520 471474 584960 471564
rect 582465 471472 584960 471474
rect 582465 471416 582470 471472
rect 582526 471416 584960 471472
rect 582465 471414 584960 471416
rect 582465 471411 582531 471414
rect 583520 471324 584960 471414
rect 336733 470794 336799 470797
rect 535729 470794 535795 470797
rect 336733 470792 340124 470794
rect 336733 470736 336738 470792
rect 336794 470736 340124 470792
rect 336733 470734 340124 470736
rect 533140 470792 535795 470794
rect 533140 470736 535734 470792
rect 535790 470736 535795 470792
rect 533140 470734 535795 470736
rect 336733 470731 336799 470734
rect 535729 470731 535795 470734
rect 245837 469026 245903 469029
rect 243892 469024 245903 469026
rect 243892 468968 245842 469024
rect 245898 468968 245903 469024
rect 243892 468966 245903 468968
rect 245837 468963 245903 468966
rect 60733 468346 60799 468349
rect 60733 468344 64124 468346
rect 60733 468288 60738 468344
rect 60794 468288 64124 468344
rect 60733 468286 64124 468288
rect 60733 468283 60799 468286
rect 338021 468074 338087 468077
rect 535729 468074 535795 468077
rect 338021 468072 340124 468074
rect 338021 468016 338026 468072
rect 338082 468016 340124 468072
rect 338021 468014 340124 468016
rect 533140 468072 535795 468074
rect 533140 468016 535734 468072
rect 535790 468016 535795 468072
rect 533140 468014 535795 468016
rect 338021 468011 338087 468014
rect 535729 468011 535795 468014
rect 245837 465626 245903 465629
rect 243892 465624 245903 465626
rect 243892 465568 245842 465624
rect 245898 465568 245903 465624
rect 243892 465566 245903 465568
rect 245837 465563 245903 465566
rect 337653 465354 337719 465357
rect 535729 465354 535795 465357
rect 337653 465352 340124 465354
rect 337653 465296 337658 465352
rect 337714 465296 340124 465352
rect 337653 465294 340124 465296
rect 533140 465352 535795 465354
rect 533140 465296 535734 465352
rect 535790 465296 535795 465352
rect 533140 465294 535795 465296
rect 337653 465291 337719 465294
rect 535729 465291 535795 465294
rect 60733 464946 60799 464949
rect 60733 464944 64124 464946
rect 60733 464888 60738 464944
rect 60794 464888 64124 464944
rect 60733 464886 64124 464888
rect 60733 464883 60799 464886
rect 293861 464402 293927 464405
rect 324262 464402 324268 464404
rect 293861 464400 324268 464402
rect 293861 464344 293866 464400
rect 293922 464344 324268 464400
rect 293861 464342 324268 464344
rect 293861 464339 293927 464342
rect 324262 464340 324268 464342
rect 324332 464340 324338 464404
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect 535729 462634 535795 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect 533140 462632 535795 462634
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 318006 462300 318012 462364
rect 318076 462362 318082 462364
rect 340094 462362 340154 462604
rect 533140 462576 535734 462632
rect 535790 462576 535795 462632
rect 533140 462574 535795 462576
rect 535729 462571 535795 462574
rect 318076 462302 340154 462362
rect 318076 462300 318082 462302
rect 245837 462226 245903 462229
rect 243892 462224 245903 462226
rect 243892 462168 245842 462224
rect 245898 462168 245903 462224
rect 243892 462166 245903 462168
rect 245837 462163 245903 462166
rect 63125 461546 63191 461549
rect 63125 461544 64124 461546
rect 63125 461488 63130 461544
rect 63186 461488 64124 461544
rect 63125 461486 64124 461488
rect 63125 461483 63191 461486
rect 337653 460594 337719 460597
rect 535729 460594 535795 460597
rect 337653 460592 340124 460594
rect 337653 460536 337658 460592
rect 337714 460536 340124 460592
rect 337653 460534 340124 460536
rect 533140 460592 535795 460594
rect 533140 460536 535734 460592
rect 535790 460536 535795 460592
rect 533140 460534 535795 460536
rect 337653 460531 337719 460534
rect 535729 460531 535795 460534
rect 245837 459506 245903 459509
rect 243892 459504 245903 459506
rect 243892 459448 245842 459504
rect 245898 459448 245903 459504
rect 243892 459446 245903 459448
rect 245837 459443 245903 459446
rect 60733 458146 60799 458149
rect 580901 458146 580967 458149
rect 582373 458146 582439 458149
rect 583520 458146 584960 458236
rect 60733 458144 64124 458146
rect 60733 458088 60738 458144
rect 60794 458088 64124 458144
rect 60733 458086 64124 458088
rect 580901 458144 584960 458146
rect 580901 458088 580906 458144
rect 580962 458088 582378 458144
rect 582434 458088 584960 458144
rect 580901 458086 584960 458088
rect 60733 458083 60799 458086
rect 580901 458083 580967 458086
rect 582373 458083 582439 458086
rect 583520 457996 584960 458086
rect 337653 457874 337719 457877
rect 535729 457874 535795 457877
rect 337653 457872 340124 457874
rect 337653 457816 337658 457872
rect 337714 457816 340124 457872
rect 337653 457814 340124 457816
rect 533140 457872 535795 457874
rect 533140 457816 535734 457872
rect 535790 457816 535795 457872
rect 533140 457814 535795 457816
rect 337653 457811 337719 457814
rect 535729 457811 535795 457814
rect 245837 456106 245903 456109
rect 243892 456104 245903 456106
rect 243892 456048 245842 456104
rect 245898 456048 245903 456104
rect 243892 456046 245903 456048
rect 245837 456043 245903 456046
rect 337653 455154 337719 455157
rect 542670 455154 542676 455156
rect 337653 455152 340124 455154
rect 337653 455096 337658 455152
rect 337714 455096 340124 455152
rect 337653 455094 340124 455096
rect 533140 455094 542676 455154
rect 337653 455091 337719 455094
rect 542670 455092 542676 455094
rect 542740 455092 542746 455156
rect 53598 454004 53604 454068
rect 53668 454066 53674 454068
rect 64094 454066 64154 454716
rect 53668 454006 64154 454066
rect 53668 454004 53674 454006
rect 337561 453114 337627 453117
rect 535729 453114 535795 453117
rect 337561 453112 340124 453114
rect 337561 453056 337566 453112
rect 337622 453056 340124 453112
rect 337561 453054 340124 453056
rect 533140 453112 535795 453114
rect 533140 453056 535734 453112
rect 535790 453056 535795 453112
rect 533140 453054 535795 453056
rect 337561 453051 337627 453054
rect 535729 453051 535795 453054
rect 245837 452706 245903 452709
rect 243892 452704 245903 452706
rect 243892 452648 245842 452704
rect 245898 452648 245903 452704
rect 243892 452646 245903 452648
rect 245837 452643 245903 452646
rect 60733 452026 60799 452029
rect 60733 452024 64124 452026
rect 60733 451968 60738 452024
rect 60794 451968 64124 452024
rect 60733 451966 64124 451968
rect 60733 451963 60799 451966
rect 337285 450394 337351 450397
rect 534206 450394 534212 450396
rect 337285 450392 340124 450394
rect 337285 450336 337290 450392
rect 337346 450336 340124 450392
rect 337285 450334 340124 450336
rect 533140 450334 534212 450394
rect 337285 450331 337351 450334
rect 534206 450332 534212 450334
rect 534276 450332 534282 450396
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 246430 449306 246436 449308
rect 243892 449246 246436 449306
rect 246430 449244 246436 449246
rect 246500 449244 246506 449308
rect 61837 448626 61903 448629
rect 61837 448624 64124 448626
rect 61837 448568 61842 448624
rect 61898 448568 64124 448624
rect 61837 448566 64124 448568
rect 61837 448563 61903 448566
rect 337101 447674 337167 447677
rect 535729 447674 535795 447677
rect 337101 447672 340124 447674
rect 337101 447616 337106 447672
rect 337162 447616 340124 447672
rect 337101 447614 340124 447616
rect 533140 447672 535795 447674
rect 533140 447616 535734 447672
rect 535790 447616 535795 447672
rect 533140 447614 535795 447616
rect 337101 447611 337167 447614
rect 535729 447611 535795 447614
rect 245837 445906 245903 445909
rect 243892 445904 245903 445906
rect 243892 445848 245842 445904
rect 245898 445848 245903 445904
rect 243892 445846 245903 445848
rect 245837 445843 245903 445846
rect 60733 445226 60799 445229
rect 60733 445224 64124 445226
rect 60733 445168 60738 445224
rect 60794 445168 64124 445224
rect 60733 445166 64124 445168
rect 60733 445163 60799 445166
rect 338021 444954 338087 444957
rect 535729 444954 535795 444957
rect 338021 444952 340124 444954
rect 338021 444896 338026 444952
rect 338082 444896 340124 444952
rect 338021 444894 340124 444896
rect 533140 444952 535795 444954
rect 533140 444896 535734 444952
rect 535790 444896 535795 444952
rect 533140 444894 535795 444896
rect 338021 444891 338087 444894
rect 535729 444891 535795 444894
rect 583520 444668 584960 444908
rect 339166 442852 339172 442916
rect 339236 442914 339242 442916
rect 535729 442914 535795 442917
rect 339236 442854 340124 442914
rect 533140 442912 535795 442914
rect 533140 442856 535734 442912
rect 535790 442856 535795 442912
rect 533140 442854 535795 442856
rect 339236 442852 339242 442854
rect 535729 442851 535795 442854
rect 246389 442506 246455 442509
rect 243892 442504 246455 442506
rect 243892 442448 246394 442504
rect 246450 442448 246455 442504
rect 243892 442446 246455 442448
rect 246389 442443 246455 442446
rect 60733 441826 60799 441829
rect 60733 441824 64124 441826
rect 60733 441768 60738 441824
rect 60794 441768 64124 441824
rect 60733 441766 64124 441768
rect 60733 441763 60799 441766
rect 337285 440194 337351 440197
rect 536925 440194 536991 440197
rect 337285 440192 340124 440194
rect 337285 440136 337290 440192
rect 337346 440136 340124 440192
rect 337285 440134 340124 440136
rect 533140 440192 536991 440194
rect 533140 440136 536930 440192
rect 536986 440136 536991 440192
rect 533140 440134 536991 440136
rect 337285 440131 337351 440134
rect 536925 440131 536991 440134
rect 245837 439106 245903 439109
rect 243892 439104 245903 439106
rect 243892 439048 245842 439104
rect 245898 439048 245903 439104
rect 243892 439046 245903 439048
rect 245837 439043 245903 439046
rect 63350 438364 63356 438428
rect 63420 438426 63426 438428
rect 63420 438366 64124 438426
rect 63420 438364 63426 438366
rect 337285 437474 337351 437477
rect 543774 437474 543780 437476
rect 337285 437472 340124 437474
rect 337285 437416 337290 437472
rect 337346 437416 340124 437472
rect 337285 437414 340124 437416
rect 533140 437414 543780 437474
rect 337285 437411 337351 437414
rect 543774 437412 543780 437414
rect 543844 437412 543850 437476
rect 63217 436794 63283 436797
rect 63534 436794 63540 436796
rect 63217 436792 63540 436794
rect -960 436508 480 436748
rect 63217 436736 63222 436792
rect 63278 436736 63540 436792
rect 63217 436734 63540 436736
rect 63217 436731 63283 436734
rect 63534 436732 63540 436734
rect 63604 436732 63610 436796
rect 245745 435706 245811 435709
rect 243892 435704 245811 435706
rect 243892 435648 245750 435704
rect 245806 435648 245811 435704
rect 243892 435646 245811 435648
rect 245745 435643 245811 435646
rect 337377 435434 337443 435437
rect 535729 435434 535795 435437
rect 337377 435432 340124 435434
rect 337377 435376 337382 435432
rect 337438 435376 340124 435432
rect 337377 435374 340124 435376
rect 533140 435432 535795 435434
rect 533140 435376 535734 435432
rect 535790 435376 535795 435432
rect 533140 435374 535795 435376
rect 337377 435371 337443 435374
rect 535729 435371 535795 435374
rect 63401 435026 63467 435029
rect 63401 435024 64124 435026
rect 63401 434968 63406 435024
rect 63462 434968 64124 435024
rect 63401 434966 64124 434968
rect 63401 434963 63467 434966
rect 337653 432714 337719 432717
rect 535729 432714 535795 432717
rect 337653 432712 340124 432714
rect 337653 432656 337658 432712
rect 337714 432656 340124 432712
rect 337653 432654 340124 432656
rect 533140 432712 535795 432714
rect 533140 432656 535734 432712
rect 535790 432656 535795 432712
rect 533140 432654 535795 432656
rect 337653 432651 337719 432654
rect 535729 432651 535795 432654
rect 245837 432306 245903 432309
rect 243892 432304 245903 432306
rect 243892 432248 245842 432304
rect 245898 432248 245903 432304
rect 243892 432246 245903 432248
rect 245837 432243 245903 432246
rect 60733 431626 60799 431629
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 60733 431624 64124 431626
rect 60733 431568 60738 431624
rect 60794 431568 64124 431624
rect 60733 431566 64124 431568
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 60733 431563 60799 431566
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 336917 429994 336983 429997
rect 534349 429994 534415 429997
rect 336917 429992 340124 429994
rect 336917 429936 336922 429992
rect 336978 429936 340124 429992
rect 336917 429934 340124 429936
rect 533140 429992 534415 429994
rect 533140 429936 534354 429992
rect 534410 429936 534415 429992
rect 533140 429934 534415 429936
rect 336917 429931 336983 429934
rect 534349 429931 534415 429934
rect 245745 428906 245811 428909
rect 243892 428904 245811 428906
rect 243892 428848 245750 428904
rect 245806 428848 245811 428904
rect 243892 428846 245811 428848
rect 245745 428843 245811 428846
rect 60733 428226 60799 428229
rect 60733 428224 64124 428226
rect 60733 428168 60738 428224
rect 60794 428168 64124 428224
rect 60733 428166 64124 428168
rect 60733 428163 60799 428166
rect 336917 427274 336983 427277
rect 535821 427274 535887 427277
rect 336917 427272 340124 427274
rect 336917 427216 336922 427272
rect 336978 427216 340124 427272
rect 336917 427214 340124 427216
rect 533140 427272 535887 427274
rect 533140 427216 535826 427272
rect 535882 427216 535887 427272
rect 533140 427214 535887 427216
rect 336917 427211 336983 427214
rect 535821 427211 535887 427214
rect 245837 425506 245903 425509
rect 243892 425504 245903 425506
rect 243892 425448 245842 425504
rect 245898 425448 245903 425504
rect 243892 425446 245903 425448
rect 245837 425443 245903 425446
rect 337653 425234 337719 425237
rect 541014 425234 541020 425236
rect 337653 425232 340124 425234
rect 337653 425176 337658 425232
rect 337714 425176 340124 425232
rect 337653 425174 340124 425176
rect 533140 425174 541020 425234
rect 337653 425171 337719 425174
rect 541014 425172 541020 425174
rect 541084 425172 541090 425236
rect 60733 424826 60799 424829
rect 60733 424824 64124 424826
rect 60733 424768 60738 424824
rect 60794 424768 64124 424824
rect 60733 424766 64124 424768
rect 60733 424763 60799 424766
rect -960 423602 480 423692
rect 4061 423602 4127 423605
rect -960 423600 4127 423602
rect -960 423544 4066 423600
rect 4122 423544 4127 423600
rect -960 423542 4127 423544
rect -960 423452 480 423542
rect 4061 423539 4127 423542
rect 337653 422514 337719 422517
rect 535821 422514 535887 422517
rect 337653 422512 340124 422514
rect 337653 422456 337658 422512
rect 337714 422456 340124 422512
rect 337653 422454 340124 422456
rect 533140 422512 535887 422514
rect 533140 422456 535826 422512
rect 535882 422456 535887 422512
rect 533140 422454 535887 422456
rect 337653 422451 337719 422454
rect 535821 422451 535887 422454
rect 245745 422106 245811 422109
rect 243892 422104 245811 422106
rect 243892 422048 245750 422104
rect 245806 422048 245811 422104
rect 243892 422046 245811 422048
rect 245745 422043 245811 422046
rect 60733 421426 60799 421429
rect 60733 421424 64124 421426
rect 60733 421368 60738 421424
rect 60794 421368 64124 421424
rect 60733 421366 64124 421368
rect 60733 421363 60799 421366
rect 337510 419732 337516 419796
rect 337580 419794 337586 419796
rect 535821 419794 535887 419797
rect 337580 419734 340124 419794
rect 533140 419792 535887 419794
rect 533140 419736 535826 419792
rect 535882 419736 535887 419792
rect 533140 419734 535887 419736
rect 337580 419732 337586 419734
rect 535821 419731 535887 419734
rect 244365 418706 244431 418709
rect 243892 418704 244431 418706
rect 243892 418648 244370 418704
rect 244426 418648 244431 418704
rect 243892 418646 244431 418648
rect 244365 418643 244431 418646
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 61009 418026 61075 418029
rect 63493 418026 63559 418029
rect 61009 418024 64124 418026
rect 61009 417968 61014 418024
rect 61070 417968 63498 418024
rect 63554 417968 64124 418024
rect 61009 417966 64124 417968
rect 61009 417963 61075 417966
rect 63493 417963 63559 417966
rect 337837 417754 337903 417757
rect 535821 417754 535887 417757
rect 337837 417752 340124 417754
rect 337837 417696 337842 417752
rect 337898 417696 340124 417752
rect 337837 417694 340124 417696
rect 533140 417752 535887 417754
rect 533140 417696 535826 417752
rect 535882 417696 535887 417752
rect 533140 417694 535887 417696
rect 337837 417691 337903 417694
rect 535821 417691 535887 417694
rect 245837 415306 245903 415309
rect 243892 415304 245903 415306
rect 243892 415248 245842 415304
rect 245898 415248 245903 415304
rect 243892 415246 245903 415248
rect 245837 415243 245903 415246
rect 335854 414972 335860 415036
rect 335924 415034 335930 415036
rect 336825 415034 336891 415037
rect 535821 415034 535887 415037
rect 335924 415032 340124 415034
rect 335924 414976 336830 415032
rect 336886 414976 340124 415032
rect 335924 414974 340124 414976
rect 533140 415032 535887 415034
rect 533140 414976 535826 415032
rect 535882 414976 535887 415032
rect 533140 414974 535887 414976
rect 335924 414972 335930 414974
rect 336825 414971 336891 414974
rect 535821 414971 535887 414974
rect 60825 414626 60891 414629
rect 63309 414626 63375 414629
rect 60825 414624 64124 414626
rect 60825 414568 60830 414624
rect 60886 414568 63314 414624
rect 63370 414568 64124 414624
rect 60825 414566 64124 414568
rect 60825 414563 60891 414566
rect 63309 414563 63375 414566
rect 337377 412314 337443 412317
rect 535821 412314 535887 412317
rect 337377 412312 340124 412314
rect 337377 412256 337382 412312
rect 337438 412256 340124 412312
rect 337377 412254 340124 412256
rect 533140 412312 535887 412314
rect 533140 412256 535826 412312
rect 535882 412256 535887 412312
rect 533140 412254 535887 412256
rect 337377 412251 337443 412254
rect 535821 412251 535887 412254
rect 245837 411906 245903 411909
rect 243892 411904 245903 411906
rect 243892 411848 245842 411904
rect 245898 411848 245903 411904
rect 243892 411846 245903 411848
rect 245837 411843 245903 411846
rect 63217 411362 63283 411365
rect 63534 411362 63540 411364
rect 63217 411360 63540 411362
rect 63217 411304 63222 411360
rect 63278 411304 63540 411360
rect 63217 411302 63540 411304
rect 63217 411299 63283 411302
rect 63534 411300 63540 411302
rect 63604 411300 63610 411364
rect 63534 411164 63540 411228
rect 63604 411226 63610 411228
rect 63604 411166 64124 411226
rect 63604 411164 63610 411166
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 336917 409594 336983 409597
rect 533429 409594 533495 409597
rect 336917 409592 340124 409594
rect 336917 409536 336922 409592
rect 336978 409536 340124 409592
rect 336917 409534 340124 409536
rect 533140 409592 533495 409594
rect 533140 409536 533434 409592
rect 533490 409536 533495 409592
rect 533140 409534 533495 409536
rect 336917 409531 336983 409534
rect 533429 409531 533495 409534
rect 245837 409186 245903 409189
rect 243892 409184 245903 409186
rect 243892 409128 245842 409184
rect 245898 409128 245903 409184
rect 243892 409126 245903 409128
rect 245837 409123 245903 409126
rect 60733 407826 60799 407829
rect 60733 407824 64124 407826
rect 60733 407768 60738 407824
rect 60794 407768 64124 407824
rect 60733 407766 64124 407768
rect 60733 407763 60799 407766
rect 337653 407554 337719 407557
rect 534257 407554 534323 407557
rect 337653 407552 340124 407554
rect 337653 407496 337658 407552
rect 337714 407496 340124 407552
rect 337653 407494 340124 407496
rect 533140 407552 534323 407554
rect 533140 407496 534262 407552
rect 534318 407496 534323 407552
rect 533140 407494 534323 407496
rect 337653 407491 337719 407494
rect 534257 407491 534323 407494
rect 245837 405786 245903 405789
rect 243892 405784 245903 405786
rect 243892 405728 245842 405784
rect 245898 405728 245903 405784
rect 243892 405726 245903 405728
rect 245837 405723 245903 405726
rect 327349 405650 327415 405653
rect 327809 405650 327875 405653
rect 327349 405648 327875 405650
rect 327349 405592 327354 405648
rect 327410 405592 327814 405648
rect 327870 405592 327875 405648
rect 327349 405590 327875 405592
rect 327349 405587 327415 405590
rect 327809 405587 327875 405590
rect 63350 405044 63356 405108
rect 63420 405106 63426 405108
rect 140589 405106 140655 405109
rect 63420 405104 140655 405106
rect 63420 405048 140594 405104
rect 140650 405048 140655 405104
rect 63420 405046 140655 405048
rect 63420 405044 63426 405046
rect 140589 405043 140655 405046
rect 63166 404908 63172 404972
rect 63236 404970 63242 404972
rect 327349 404970 327415 404973
rect 63236 404968 327415 404970
rect 63236 404912 327354 404968
rect 327410 404912 327415 404968
rect 63236 404910 327415 404912
rect 63236 404908 63242 404910
rect 327349 404907 327415 404910
rect 579705 404970 579771 404973
rect 583520 404970 584960 405060
rect 579705 404968 584960 404970
rect 579705 404912 579710 404968
rect 579766 404912 584960 404968
rect 579705 404910 584960 404912
rect 579705 404907 579771 404910
rect 337745 404834 337811 404837
rect 535453 404834 535519 404837
rect 337745 404832 340124 404834
rect 337745 404776 337750 404832
rect 337806 404776 340124 404832
rect 337745 404774 340124 404776
rect 533140 404832 535519 404834
rect 533140 404776 535458 404832
rect 535514 404776 535519 404832
rect 583520 404820 584960 404910
rect 533140 404774 535519 404776
rect 337745 404771 337811 404774
rect 535453 404771 535519 404774
rect 61878 404364 61884 404428
rect 61948 404426 61954 404428
rect 64873 404426 64939 404429
rect 61948 404424 64939 404426
rect 61948 404368 64878 404424
rect 64934 404368 64939 404424
rect 61948 404366 64939 404368
rect 61948 404364 61954 404366
rect 64873 404363 64939 404366
rect 59118 403548 59124 403612
rect 59188 403610 59194 403612
rect 104985 403610 105051 403613
rect 59188 403608 105051 403610
rect 59188 403552 104990 403608
rect 105046 403552 105051 403608
rect 59188 403550 105051 403552
rect 59188 403548 59194 403550
rect 104985 403547 105051 403550
rect 50838 402188 50844 402252
rect 50908 402250 50914 402252
rect 80697 402250 80763 402253
rect 50908 402248 80763 402250
rect 50908 402192 80702 402248
rect 80758 402192 80763 402248
rect 50908 402190 80763 402192
rect 50908 402188 50914 402190
rect 80697 402187 80763 402190
rect 108481 402250 108547 402253
rect 125726 402250 125732 402252
rect 108481 402248 125732 402250
rect 108481 402192 108486 402248
rect 108542 402192 125732 402248
rect 108481 402190 125732 402192
rect 108481 402187 108547 402190
rect 125726 402188 125732 402190
rect 125796 402188 125802 402252
rect 166758 402188 166764 402252
rect 166828 402250 166834 402252
rect 225689 402250 225755 402253
rect 166828 402248 225755 402250
rect 166828 402192 225694 402248
rect 225750 402192 225755 402248
rect 166828 402190 225755 402192
rect 166828 402188 166834 402190
rect 225689 402187 225755 402190
rect 535821 402114 535887 402117
rect 533140 402112 535887 402114
rect 138606 401644 138612 401708
rect 138676 401706 138682 401708
rect 140037 401706 140103 401709
rect 138676 401704 140103 401706
rect 138676 401648 140042 401704
rect 140098 401648 140103 401704
rect 138676 401646 140103 401648
rect 138676 401644 138682 401646
rect 140037 401643 140103 401646
rect 337469 401706 337535 401709
rect 338021 401706 338087 401709
rect 340094 401706 340154 402084
rect 533140 402056 535826 402112
rect 535882 402056 535887 402112
rect 533140 402054 535887 402056
rect 535821 402051 535887 402054
rect 337469 401704 340154 401706
rect 337469 401648 337474 401704
rect 337530 401648 338026 401704
rect 338082 401648 340154 401704
rect 337469 401646 340154 401648
rect 337469 401643 337535 401646
rect 338021 401643 338087 401646
rect 84837 400890 84903 400893
rect 98821 400890 98887 400893
rect 340270 400890 340276 400892
rect 84837 400888 340276 400890
rect 84837 400832 84842 400888
rect 84898 400832 98826 400888
rect 98882 400832 340276 400888
rect 84837 400830 340276 400832
rect 84837 400827 84903 400830
rect 98821 400827 98887 400830
rect 340270 400828 340276 400830
rect 340340 400828 340346 400892
rect 533429 400074 533495 400077
rect 533140 400072 533495 400074
rect 533140 400016 533434 400072
rect 533490 400016 533495 400072
rect 533140 400014 533495 400016
rect 533429 400011 533495 400014
rect 246246 399876 246252 399940
rect 246316 399938 246322 399940
rect 246573 399938 246639 399941
rect 550725 399938 550791 399941
rect 246316 399936 550791 399938
rect 246316 399880 246578 399936
rect 246634 399880 550730 399936
rect 550786 399880 550791 399936
rect 246316 399878 550791 399880
rect 246316 399876 246322 399878
rect 246573 399875 246639 399878
rect 550725 399875 550791 399878
rect 246430 399740 246436 399804
rect 246500 399802 246506 399804
rect 550633 399802 550699 399805
rect 246500 399800 550699 399802
rect 246500 399744 550638 399800
rect 550694 399744 550699 399800
rect 246500 399742 550699 399744
rect 246500 399740 246506 399742
rect 550633 399739 550699 399742
rect 55070 399468 55076 399532
rect 55140 399530 55146 399532
rect 88977 399530 89043 399533
rect 55140 399528 89043 399530
rect 55140 399472 88982 399528
rect 89038 399472 89043 399528
rect 55140 399470 89043 399472
rect 55140 399468 55146 399470
rect 88977 399467 89043 399470
rect 339166 398788 339172 398852
rect 339236 398850 339242 398852
rect 339401 398850 339467 398853
rect 339236 398848 339467 398850
rect 339236 398792 339406 398848
rect 339462 398792 339467 398848
rect 339236 398790 339467 398792
rect 339236 398788 339242 398790
rect 339401 398787 339467 398790
rect 242934 398652 242940 398716
rect 243004 398714 243010 398716
rect 244181 398714 244247 398717
rect 547965 398714 548031 398717
rect 243004 398712 548031 398714
rect 243004 398656 244186 398712
rect 244242 398656 547970 398712
rect 548026 398656 548031 398712
rect 243004 398654 548031 398656
rect 243004 398652 243010 398654
rect 244181 398651 244247 398654
rect 547965 398651 548031 398654
rect 546493 398578 546559 398581
rect 287010 398576 546559 398578
rect 287010 398520 546498 398576
rect 546554 398520 546559 398576
rect 287010 398518 546559 398520
rect 280797 398306 280863 398309
rect 281441 398306 281507 398309
rect 287010 398306 287070 398518
rect 546493 398515 546559 398518
rect 340270 398380 340276 398444
rect 340340 398442 340346 398444
rect 376753 398442 376819 398445
rect 377949 398442 378015 398445
rect 340340 398440 378015 398442
rect 340340 398384 376758 398440
rect 376814 398384 377954 398440
rect 378010 398384 378015 398440
rect 340340 398382 378015 398384
rect 340340 398380 340346 398382
rect 376753 398379 376819 398382
rect 377949 398379 378015 398382
rect 280797 398304 287070 398306
rect 280797 398248 280802 398304
rect 280858 398248 281446 398304
rect 281502 398248 287070 398304
rect 280797 398246 287070 398248
rect 280797 398243 280863 398246
rect 281441 398243 281507 398246
rect -960 397490 480 397580
rect 3969 397490 4035 397493
rect -960 397488 4035 397490
rect -960 397432 3974 397488
rect 4030 397432 4035 397488
rect -960 397430 4035 397432
rect -960 397340 480 397430
rect 3969 397427 4035 397430
rect 331121 396810 331187 396813
rect 343633 396810 343699 396813
rect 331121 396808 343699 396810
rect 331121 396752 331126 396808
rect 331182 396752 343638 396808
rect 343694 396752 343699 396808
rect 331121 396750 343699 396752
rect 331121 396747 331187 396750
rect 343633 396747 343699 396750
rect 328361 396674 328427 396677
rect 354673 396674 354739 396677
rect 328361 396672 354739 396674
rect 328361 396616 328366 396672
rect 328422 396616 354678 396672
rect 354734 396616 354739 396672
rect 328361 396614 354739 396616
rect 328361 396611 328427 396614
rect 354673 396611 354739 396614
rect 498837 396674 498903 396677
rect 539542 396674 539548 396676
rect 498837 396672 539548 396674
rect 498837 396616 498842 396672
rect 498898 396616 539548 396672
rect 498837 396614 539548 396616
rect 498837 396611 498903 396614
rect 539542 396612 539548 396614
rect 539612 396612 539618 396676
rect 338982 395388 338988 395452
rect 339052 395450 339058 395452
rect 421005 395450 421071 395453
rect 339052 395448 421071 395450
rect 339052 395392 421010 395448
rect 421066 395392 421071 395448
rect 339052 395390 421071 395392
rect 339052 395388 339058 395390
rect 421005 395387 421071 395390
rect 508497 395450 508563 395453
rect 541014 395450 541020 395452
rect 508497 395448 541020 395450
rect 508497 395392 508502 395448
rect 508558 395392 541020 395448
rect 508497 395390 541020 395392
rect 508497 395387 508563 395390
rect 541014 395388 541020 395390
rect 541084 395388 541090 395452
rect 177062 395252 177068 395316
rect 177132 395314 177138 395316
rect 536782 395314 536788 395316
rect 177132 395254 536788 395314
rect 177132 395252 177138 395254
rect 536782 395252 536788 395254
rect 536852 395252 536858 395316
rect 59077 393274 59143 393277
rect 543774 393274 543780 393276
rect 59077 393272 543780 393274
rect 59077 393216 59082 393272
rect 59138 393216 543780 393272
rect 59077 393214 543780 393216
rect 59077 393211 59143 393214
rect 543774 393212 543780 393214
rect 543844 393212 543850 393276
rect 58617 392050 58683 392053
rect 59077 392050 59143 392053
rect 58617 392048 59143 392050
rect 58617 391992 58622 392048
rect 58678 391992 59082 392048
rect 59138 391992 59143 392048
rect 58617 391990 59143 391992
rect 58617 391987 58683 391990
rect 59077 391987 59143 391990
rect 583520 391628 584960 391868
rect 53598 391308 53604 391372
rect 53668 391370 53674 391372
rect 120022 391370 120028 391372
rect 53668 391310 120028 391370
rect 53668 391308 53674 391310
rect 120022 391308 120028 391310
rect 120092 391308 120098 391372
rect 46606 391172 46612 391236
rect 46676 391234 46682 391236
rect 116577 391234 116643 391237
rect 46676 391232 116643 391234
rect 46676 391176 116582 391232
rect 116638 391176 116643 391232
rect 46676 391174 116643 391176
rect 46676 391172 46682 391174
rect 116577 391171 116643 391174
rect 130377 389874 130443 389877
rect 246430 389874 246436 389876
rect 130377 389872 246436 389874
rect 130377 389816 130382 389872
rect 130438 389816 246436 389872
rect 130377 389814 246436 389816
rect 130377 389811 130443 389814
rect 246430 389812 246436 389814
rect 246500 389812 246506 389876
rect 238017 389194 238083 389197
rect 238661 389194 238727 389197
rect 295558 389194 295564 389196
rect 238017 389192 295564 389194
rect 238017 389136 238022 389192
rect 238078 389136 238666 389192
rect 238722 389136 295564 389192
rect 238017 389134 295564 389136
rect 238017 389131 238083 389134
rect 238661 389131 238727 389134
rect 295558 389132 295564 389134
rect 295628 389132 295634 389196
rect 434805 387698 434871 387701
rect 439078 387698 439084 387700
rect 434805 387696 439084 387698
rect 434805 387640 434810 387696
rect 434866 387640 439084 387696
rect 434805 387638 439084 387640
rect 434805 387635 434871 387638
rect 439078 387636 439084 387638
rect 439148 387636 439154 387700
rect 63534 386956 63540 387020
rect 63604 387018 63610 387020
rect 125593 387018 125659 387021
rect 63604 387016 125659 387018
rect 63604 386960 125598 387016
rect 125654 386960 125659 387016
rect 63604 386958 125659 386960
rect 63604 386956 63610 386958
rect 125593 386955 125659 386958
rect -960 384284 480 384524
rect 345749 382938 345815 382941
rect 542670 382938 542676 382940
rect 345749 382936 542676 382938
rect 345749 382880 345754 382936
rect 345810 382880 542676 382936
rect 345749 382878 542676 382880
rect 345749 382875 345815 382878
rect 542670 382876 542676 382878
rect 542740 382876 542746 382940
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 176377 373282 176443 373285
rect 337326 373282 337332 373284
rect 176377 373280 337332 373282
rect 176377 373224 176382 373280
rect 176438 373224 337332 373280
rect 176377 373222 337332 373224
rect 176377 373219 176443 373222
rect 337326 373220 337332 373222
rect 337396 373220 337402 373284
rect 176285 371922 176351 371925
rect 337510 371922 337516 371924
rect 176285 371920 337516 371922
rect 176285 371864 176290 371920
rect 176346 371864 337516 371920
rect 176285 371862 337516 371864
rect 176285 371859 176351 371862
rect 337510 371860 337516 371862
rect 337580 371860 337586 371924
rect -960 371378 480 371468
rect 2957 371378 3023 371381
rect -960 371376 3023 371378
rect -960 371320 2962 371376
rect 3018 371320 3023 371376
rect -960 371318 3023 371320
rect -960 371228 480 371318
rect 2957 371315 3023 371318
rect 57646 370500 57652 370564
rect 57716 370562 57722 370564
rect 113817 370562 113883 370565
rect 57716 370560 113883 370562
rect 57716 370504 113822 370560
rect 113878 370504 113883 370560
rect 57716 370502 113883 370504
rect 57716 370500 57722 370502
rect 113817 370499 113883 370502
rect 309225 369884 309291 369885
rect 309174 369882 309180 369884
rect 309134 369822 309180 369882
rect 309244 369880 309291 369884
rect 309286 369824 309291 369880
rect 309174 369820 309180 369822
rect 309244 369820 309291 369824
rect 309225 369819 309291 369820
rect 135989 368658 136055 368661
rect 295374 368658 295380 368660
rect 135989 368656 295380 368658
rect 135989 368600 135994 368656
rect 136050 368600 295380 368656
rect 135989 368598 295380 368600
rect 135989 368595 136055 368598
rect 295374 368596 295380 368598
rect 295444 368596 295450 368660
rect 180793 368522 180859 368525
rect 342846 368522 342852 368524
rect 180793 368520 342852 368522
rect 180793 368464 180798 368520
rect 180854 368464 342852 368520
rect 180793 368462 342852 368464
rect 180793 368459 180859 368462
rect 342846 368460 342852 368462
rect 342916 368460 342922 368524
rect 148174 366284 148180 366348
rect 148244 366346 148250 366348
rect 228357 366346 228423 366349
rect 148244 366344 228423 366346
rect 148244 366288 228362 366344
rect 228418 366288 228423 366344
rect 148244 366286 228423 366288
rect 148244 366284 148250 366286
rect 228357 366283 228423 366286
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 58934 364924 58940 364988
rect 59004 364986 59010 364988
rect 98729 364986 98795 364989
rect 59004 364984 98795 364986
rect 59004 364928 98734 364984
rect 98790 364928 98795 364984
rect 583520 364972 584960 365062
rect 59004 364926 98795 364928
rect 59004 364924 59010 364926
rect 98729 364923 98795 364926
rect 340137 362812 340203 362813
rect 340086 362810 340092 362812
rect 340046 362750 340092 362810
rect 340156 362808 340203 362812
rect 340198 362752 340203 362808
rect 340086 362748 340092 362750
rect 340156 362748 340203 362752
rect 340137 362747 340203 362748
rect 175181 362266 175247 362269
rect 340137 362266 340203 362269
rect 175181 362264 340203 362266
rect 175181 362208 175186 362264
rect 175242 362208 340142 362264
rect 340198 362208 340203 362264
rect 175181 362206 340203 362208
rect 175181 362203 175247 362206
rect 340137 362203 340203 362206
rect 260741 360906 260807 360909
rect 299606 360906 299612 360908
rect 260741 360904 299612 360906
rect 260741 360848 260746 360904
rect 260802 360848 299612 360904
rect 260741 360846 299612 360848
rect 260741 360843 260807 360846
rect 299606 360844 299612 360846
rect 299676 360844 299682 360908
rect 340086 360906 340092 360908
rect 335310 360846 340092 360906
rect 191741 360226 191807 360229
rect 335310 360226 335370 360846
rect 340086 360844 340092 360846
rect 340156 360906 340162 360908
rect 538438 360906 538444 360908
rect 340156 360846 538444 360906
rect 340156 360844 340162 360846
rect 538438 360844 538444 360846
rect 538508 360844 538514 360908
rect 191741 360224 335370 360226
rect 191741 360168 191746 360224
rect 191802 360168 335370 360224
rect 191741 360166 335370 360168
rect 191741 360163 191807 360166
rect 233785 358866 233851 358869
rect 336774 358866 336780 358868
rect 233785 358864 336780 358866
rect 233785 358808 233790 358864
rect 233846 358808 336780 358864
rect 233785 358806 336780 358808
rect 233785 358803 233851 358806
rect 336774 358804 336780 358806
rect 336844 358804 336850 358868
rect 282085 358730 282151 358733
rect 282821 358730 282887 358733
rect 282085 358728 282887 358730
rect 282085 358672 282090 358728
rect 282146 358672 282826 358728
rect 282882 358672 282887 358728
rect 282085 358670 282887 358672
rect 282085 358667 282151 358670
rect 282821 358667 282887 358670
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 297950 357988 297956 358052
rect 298020 358050 298026 358052
rect 530669 358050 530735 358053
rect 298020 358048 530735 358050
rect 298020 357992 530674 358048
rect 530730 357992 530735 358048
rect 298020 357990 530735 357992
rect 298020 357988 298026 357990
rect 530669 357987 530735 357990
rect 298001 357914 298067 357917
rect 305494 357914 305500 357916
rect 298001 357912 305500 357914
rect 298001 357856 298006 357912
rect 298062 357856 305500 357912
rect 298001 357854 305500 357856
rect 298001 357851 298067 357854
rect 305494 357852 305500 357854
rect 305564 357852 305570 357916
rect 282085 357642 282151 357645
rect 291694 357642 291700 357644
rect 282085 357640 291700 357642
rect 282085 357584 282090 357640
rect 282146 357584 291700 357640
rect 282085 357582 291700 357584
rect 282085 357579 282151 357582
rect 291694 357580 291700 357582
rect 291764 357580 291770 357644
rect 157190 357444 157196 357508
rect 157260 357506 157266 357508
rect 184933 357506 184999 357509
rect 157260 357504 184999 357506
rect 157260 357448 184938 357504
rect 184994 357448 184999 357504
rect 157260 357446 184999 357448
rect 157260 357444 157266 357446
rect 184933 357443 184999 357446
rect 252461 357506 252527 357509
rect 353293 357506 353359 357509
rect 252461 357504 353359 357506
rect 252461 357448 252466 357504
rect 252522 357448 353298 357504
rect 353354 357448 353359 357504
rect 252461 357446 353359 357448
rect 252461 357443 252527 357446
rect 353293 357443 353359 357446
rect 168189 356146 168255 356149
rect 320817 356146 320883 356149
rect 168189 356144 320883 356146
rect 168189 356088 168194 356144
rect 168250 356088 320822 356144
rect 320878 356088 320883 356144
rect 168189 356086 320883 356088
rect 168189 356083 168255 356086
rect 320817 356083 320883 356086
rect 291101 356010 291167 356013
rect 294086 356010 294092 356012
rect 291101 356008 294092 356010
rect 291101 355952 291106 356008
rect 291162 355952 294092 356008
rect 291101 355950 294092 355952
rect 291101 355947 291167 355950
rect 294086 355948 294092 355950
rect 294156 355948 294162 356012
rect 179137 355330 179203 355333
rect 186957 355330 187023 355333
rect 179137 355328 187023 355330
rect 179137 355272 179142 355328
rect 179198 355272 186962 355328
rect 187018 355272 187023 355328
rect 179137 355270 187023 355272
rect 179137 355267 179203 355270
rect 186957 355267 187023 355270
rect 291837 355058 291903 355061
rect 297398 355058 297404 355060
rect 291837 355056 297404 355058
rect 291837 355000 291842 355056
rect 291898 355000 297404 355056
rect 291837 354998 297404 355000
rect 291837 354995 291903 354998
rect 297398 354996 297404 354998
rect 297468 355058 297474 355060
rect 297950 355058 297956 355060
rect 297468 354998 297956 355058
rect 297468 354996 297474 354998
rect 297950 354996 297956 354998
rect 298020 354996 298026 355060
rect 178677 354922 178743 354925
rect 305085 354922 305151 354925
rect 178677 354920 305151 354922
rect 178677 354864 178682 354920
rect 178738 354864 305090 354920
rect 305146 354864 305151 354920
rect 178677 354862 305151 354864
rect 178677 354859 178743 354862
rect 305085 354859 305151 354862
rect 200113 354786 200179 354789
rect 291837 354786 291903 354789
rect 200113 354784 291903 354786
rect 200113 354728 200118 354784
rect 200174 354728 291842 354784
rect 291898 354728 291903 354784
rect 200113 354726 291903 354728
rect 200113 354723 200179 354726
rect 291837 354723 291903 354726
rect 291193 354650 291259 354653
rect 292573 354650 292639 354653
rect 296713 354650 296779 354653
rect 291193 354648 292314 354650
rect 291193 354592 291198 354648
rect 291254 354592 292314 354648
rect 291193 354590 292314 354592
rect 291193 354587 291259 354590
rect 292254 354514 292314 354590
rect 292573 354648 296779 354650
rect 292573 354592 292578 354648
rect 292634 354592 296718 354648
rect 296774 354592 296779 354648
rect 292573 354590 296779 354592
rect 292573 354587 292639 354590
rect 296713 354587 296779 354590
rect 293309 354514 293375 354517
rect 292254 354454 292682 354514
rect 179229 354378 179295 354381
rect 292622 354378 292682 354454
rect 293309 354512 296730 354514
rect 293309 354456 293314 354512
rect 293370 354456 296730 354512
rect 293309 354454 296730 354456
rect 293309 354451 293375 354454
rect 295425 354378 295491 354381
rect 179229 354376 180044 354378
rect 179229 354320 179234 354376
rect 179290 354320 180044 354376
rect 292622 354376 295491 354378
rect 292622 354348 295430 354376
rect 179229 354318 180044 354320
rect 292652 354320 295430 354348
rect 295486 354320 295491 354376
rect 292652 354318 295491 354320
rect 179229 354315 179295 354318
rect 295425 354315 295491 354318
rect 296670 353426 296730 354454
rect 410517 353426 410583 353429
rect 296670 353424 410583 353426
rect 296670 353368 410522 353424
rect 410578 353368 410583 353424
rect 296670 353366 410583 353368
rect 410517 353363 410583 353366
rect 292614 353228 292620 353292
rect 292684 353290 292690 353292
rect 299473 353290 299539 353293
rect 292684 353288 299539 353290
rect 292684 353232 299478 353288
rect 299534 353232 299539 353288
rect 292684 353230 299539 353232
rect 292684 353228 292690 353230
rect 299473 353227 299539 353230
rect 295425 352338 295491 352341
rect 292836 352336 295491 352338
rect 292836 352280 295430 352336
rect 295486 352280 295491 352336
rect 292836 352278 295491 352280
rect 295425 352275 295491 352278
rect 179462 352210 180044 352270
rect 175038 352140 175044 352204
rect 175108 352202 175114 352204
rect 179462 352202 179522 352210
rect 175108 352142 179522 352202
rect 175108 352140 175114 352142
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 179830 350170 180044 350230
rect 179830 350029 179890 350170
rect 176510 349964 176516 350028
rect 176580 350026 176586 350028
rect 179830 350026 179939 350029
rect 176580 350024 179939 350026
rect 176580 349968 179878 350024
rect 179934 349968 179939 350024
rect 176580 349966 179939 349968
rect 176580 349964 176586 349966
rect 179873 349963 179939 349966
rect 295425 349618 295491 349621
rect 292836 349616 295491 349618
rect 292836 349560 295430 349616
rect 295486 349560 295491 349616
rect 292836 349558 295491 349560
rect 295425 349555 295491 349558
rect 179462 348130 180044 348190
rect 176653 348122 176719 348125
rect 179462 348122 179522 348130
rect 176653 348120 179522 348122
rect 176653 348064 176658 348120
rect 176714 348064 179522 348120
rect 176653 348062 179522 348064
rect 176653 348059 176719 348062
rect 295425 347578 295491 347581
rect 292836 347576 295491 347578
rect 292836 347520 295430 347576
rect 295486 347520 295491 347576
rect 292836 347518 295491 347520
rect 295425 347515 295491 347518
rect 176653 345538 176719 345541
rect 295609 345538 295675 345541
rect 176653 345536 179522 345538
rect -960 345402 480 345492
rect 176653 345480 176658 345536
rect 176714 345480 179522 345536
rect 176653 345478 179522 345480
rect 292836 345536 295675 345538
rect 292836 345480 295614 345536
rect 295670 345480 295675 345536
rect 292836 345478 295675 345480
rect 176653 345475 176719 345478
rect 179462 345470 179522 345478
rect 295609 345475 295675 345478
rect 179462 345410 180044 345470
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 177849 343498 177915 343501
rect 295425 343498 295491 343501
rect 177849 343496 179890 343498
rect 177849 343440 177854 343496
rect 177910 343440 179890 343496
rect 177849 343438 179890 343440
rect 292836 343496 295491 343498
rect 292836 343440 295430 343496
rect 295486 343440 295491 343496
rect 292836 343438 295491 343440
rect 177849 343435 177915 343438
rect 179830 343430 179890 343438
rect 295425 343435 295491 343438
rect 179830 343370 180044 343430
rect 177665 342274 177731 342277
rect 177849 342274 177915 342277
rect 177665 342272 177915 342274
rect 177665 342216 177670 342272
rect 177726 342216 177854 342272
rect 177910 342216 177915 342272
rect 177665 342214 177915 342216
rect 177665 342211 177731 342214
rect 177849 342211 177915 342214
rect 179830 341330 180044 341390
rect 176653 341322 176719 341325
rect 179830 341322 179890 341330
rect 176653 341320 179890 341322
rect 176653 341264 176658 341320
rect 176714 341264 179890 341320
rect 176653 341262 179890 341264
rect 176653 341259 176719 341262
rect 295425 340778 295491 340781
rect 292836 340776 295491 340778
rect 292836 340720 295430 340776
rect 295486 340720 295491 340776
rect 292836 340718 295491 340720
rect 295425 340715 295491 340718
rect 179462 339290 180044 339350
rect 176653 339282 176719 339285
rect 179462 339282 179522 339290
rect 176653 339280 179522 339282
rect 176653 339224 176658 339280
rect 176714 339224 179522 339280
rect 176653 339222 179522 339224
rect 176653 339219 176719 339222
rect 295425 338738 295491 338741
rect 292836 338736 295491 338738
rect 292836 338680 295430 338736
rect 295486 338680 295491 338736
rect 292836 338678 295491 338680
rect 295425 338675 295491 338678
rect 583520 338452 584960 338692
rect 174854 336636 174860 336700
rect 174924 336698 174930 336700
rect 176561 336698 176627 336701
rect 295558 336698 295564 336700
rect 174924 336696 179890 336698
rect 174924 336640 176566 336696
rect 176622 336640 179890 336696
rect 174924 336638 179890 336640
rect 292836 336638 295564 336698
rect 174924 336636 174930 336638
rect 176561 336635 176627 336638
rect 179830 336630 179890 336638
rect 295558 336636 295564 336638
rect 295628 336698 295634 336700
rect 295701 336698 295767 336701
rect 295977 336700 296043 336701
rect 295926 336698 295932 336700
rect 295628 336696 295767 336698
rect 295628 336640 295706 336696
rect 295762 336640 295767 336696
rect 295628 336638 295767 336640
rect 295886 336638 295932 336698
rect 295996 336696 296043 336700
rect 296038 336640 296043 336696
rect 295628 336636 295634 336638
rect 295701 336635 295767 336638
rect 295926 336636 295932 336638
rect 295996 336636 296043 336640
rect 295977 336635 296043 336636
rect 179830 336570 180044 336630
rect 363597 336018 363663 336021
rect 535678 336018 535684 336020
rect 363597 336016 535684 336018
rect 363597 335960 363602 336016
rect 363658 335960 535684 336016
rect 363597 335958 535684 335960
rect 363597 335955 363663 335958
rect 535678 335956 535684 335958
rect 535748 335956 535754 336020
rect 176653 334658 176719 334661
rect 176653 334656 179890 334658
rect 176653 334600 176658 334656
rect 176714 334600 179890 334656
rect 176653 334598 179890 334600
rect 176653 334595 176719 334598
rect 179830 334590 179890 334598
rect 179830 334530 180044 334590
rect 292806 334386 292866 334628
rect 295425 334388 295491 334389
rect 295374 334386 295380 334388
rect 292806 334326 295380 334386
rect 295444 334384 295491 334388
rect 295486 334328 295491 334384
rect 295374 334324 295380 334326
rect 295444 334324 295491 334328
rect 295425 334323 295491 334324
rect 176653 332618 176719 332621
rect 176653 332616 179890 332618
rect 176653 332560 176658 332616
rect 176714 332560 179890 332616
rect 176653 332558 179890 332560
rect 176653 332555 176719 332558
rect 179830 332550 179890 332558
rect 179830 332490 180044 332550
rect -960 332196 480 332436
rect 293125 331938 293191 331941
rect 293861 331938 293927 331941
rect 292836 331936 293927 331938
rect 292836 331880 293130 331936
rect 293186 331880 293866 331936
rect 293922 331880 293927 331936
rect 292836 331878 293927 331880
rect 293125 331875 293191 331878
rect 293861 331875 293927 331878
rect 179462 330450 180044 330510
rect 177849 330442 177915 330445
rect 179462 330442 179522 330450
rect 177849 330440 179522 330442
rect 177849 330384 177854 330440
rect 177910 330384 179522 330440
rect 177849 330382 179522 330384
rect 177849 330379 177915 330382
rect 295425 329898 295491 329901
rect 292836 329896 295491 329898
rect 292836 329840 295430 329896
rect 295486 329840 295491 329896
rect 292836 329838 295491 329840
rect 295425 329835 295491 329838
rect 295517 327858 295583 327861
rect 292836 327856 295583 327858
rect 292836 327800 295522 327856
rect 295578 327800 295583 327856
rect 292836 327798 295583 327800
rect 295517 327795 295583 327798
rect 179462 327730 180044 327790
rect 176561 327722 176627 327725
rect 179462 327722 179522 327730
rect 176561 327720 179522 327722
rect 176561 327664 176566 327720
rect 176622 327664 179522 327720
rect 176561 327662 179522 327664
rect 176561 327659 176627 327662
rect 296110 327660 296116 327724
rect 296180 327722 296186 327724
rect 537017 327722 537083 327725
rect 296180 327720 537083 327722
rect 296180 327664 537022 327720
rect 537078 327664 537083 327720
rect 296180 327662 537083 327664
rect 296180 327660 296186 327662
rect 537017 327659 537083 327662
rect 176653 325818 176719 325821
rect 293125 325818 293191 325821
rect 176653 325816 179522 325818
rect 176653 325760 176658 325816
rect 176714 325760 179522 325816
rect 176653 325758 179522 325760
rect 292836 325816 293191 325818
rect 292836 325760 293130 325816
rect 293186 325760 293191 325816
rect 292836 325758 293191 325760
rect 176653 325755 176719 325758
rect 179462 325750 179522 325758
rect 293125 325755 293191 325758
rect 179462 325690 180044 325750
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect 179462 323650 180044 323710
rect 176326 323580 176332 323644
rect 176396 323642 176402 323644
rect 179462 323642 179522 323650
rect 176396 323582 179522 323642
rect 176396 323580 176402 323582
rect 294321 323098 294387 323101
rect 292836 323096 294387 323098
rect 292836 323040 294326 323096
rect 294382 323040 294387 323096
rect 292836 323038 294387 323040
rect 294321 323035 294387 323038
rect 146293 322962 146359 322965
rect 149646 322962 149652 322964
rect 146293 322960 149652 322962
rect 146293 322904 146298 322960
rect 146354 322904 149652 322960
rect 146293 322902 149652 322904
rect 146293 322899 146359 322902
rect 149646 322900 149652 322902
rect 149716 322900 149722 322964
rect 179830 321610 180044 321670
rect 177573 321602 177639 321605
rect 179830 321602 179890 321610
rect 177573 321600 179890 321602
rect 177573 321544 177578 321600
rect 177634 321544 179890 321600
rect 177573 321542 179890 321544
rect 177573 321539 177639 321542
rect 295333 321058 295399 321061
rect 292836 321056 295399 321058
rect 292836 321000 295338 321056
rect 295394 321000 295399 321056
rect 292836 320998 295399 321000
rect 295333 320995 295399 320998
rect -960 319290 480 319380
rect 3141 319290 3207 319293
rect -960 319288 3207 319290
rect -960 319232 3146 319288
rect 3202 319232 3207 319288
rect -960 319230 3207 319232
rect -960 319140 480 319230
rect 3141 319227 3207 319230
rect 179137 319018 179203 319021
rect 179270 319018 179276 319020
rect 179137 319016 179276 319018
rect 179137 318960 179142 319016
rect 179198 318960 179276 319016
rect 179137 318958 179276 318960
rect 179137 318955 179203 318958
rect 179270 318956 179276 318958
rect 179340 319018 179346 319020
rect 295333 319018 295399 319021
rect 179340 318958 179890 319018
rect 292836 319016 295399 319018
rect 292836 318960 295338 319016
rect 295394 318960 295399 319016
rect 292836 318958 295399 318960
rect 179340 318956 179346 318958
rect 179830 318950 179890 318958
rect 295333 318955 295399 318958
rect 179830 318890 180044 318950
rect 295333 316978 295399 316981
rect 292836 316976 295399 316978
rect 292836 316920 295338 316976
rect 295394 316920 295399 316976
rect 292836 316918 295399 316920
rect 295333 316915 295399 316918
rect 179830 316850 180044 316910
rect 179137 316842 179203 316845
rect 179830 316842 179890 316850
rect 179137 316840 179890 316842
rect 179137 316784 179142 316840
rect 179198 316784 179890 316840
rect 179137 316782 179890 316784
rect 179137 316779 179203 316782
rect 179505 314870 179571 314873
rect 179505 314868 180044 314870
rect 179505 314812 179510 314868
rect 179566 314812 180044 314868
rect 179505 314810 180044 314812
rect 179505 314807 179571 314810
rect 295333 314258 295399 314261
rect 292836 314256 295399 314258
rect 292836 314200 295338 314256
rect 295394 314200 295399 314256
rect 292836 314198 295399 314200
rect 295333 314195 295399 314198
rect 179462 312770 180044 312830
rect 176653 312762 176719 312765
rect 179462 312762 179522 312770
rect 176653 312760 179522 312762
rect 176653 312704 176658 312760
rect 176714 312704 179522 312760
rect 176653 312702 179522 312704
rect 176653 312699 176719 312702
rect 295333 312218 295399 312221
rect 292836 312216 295399 312218
rect 292836 312160 295338 312216
rect 295394 312160 295399 312216
rect 292836 312158 295399 312160
rect 295333 312155 295399 312158
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect 176653 310178 176719 310181
rect 295333 310178 295399 310181
rect 176653 310176 179890 310178
rect 176653 310120 176658 310176
rect 176714 310120 179890 310176
rect 176653 310118 179890 310120
rect 292836 310176 295399 310178
rect 292836 310120 295338 310176
rect 295394 310120 295399 310176
rect 292836 310118 295399 310120
rect 176653 310115 176719 310118
rect 179830 310110 179890 310118
rect 295333 310115 295399 310118
rect 179830 310050 180044 310110
rect 77937 309090 78003 309093
rect 78581 309090 78647 309093
rect 77937 309088 78647 309090
rect 77937 309032 77942 309088
rect 77998 309032 78586 309088
rect 78642 309032 78647 309088
rect 77937 309030 78647 309032
rect 77937 309027 78003 309030
rect 78581 309027 78647 309030
rect 292614 308620 292620 308684
rect 292684 308620 292690 308684
rect 179505 308070 179571 308073
rect 179505 308068 180044 308070
rect 179505 308012 179510 308068
rect 179566 308012 180044 308068
rect 179505 308010 180044 308012
rect 179505 308007 179571 308010
rect 77937 307866 78003 307869
rect 142654 307866 142660 307868
rect 77937 307864 142660 307866
rect 77937 307808 77942 307864
rect 77998 307808 142660 307864
rect 77937 307806 142660 307808
rect 77937 307803 78003 307806
rect 142654 307804 142660 307806
rect 142724 307804 142730 307868
rect 292622 307866 292682 308620
rect 295333 307866 295399 307869
rect 292622 307864 295399 307866
rect 292622 307808 295338 307864
rect 295394 307808 295399 307864
rect 292622 307806 295399 307808
rect 295333 307803 295399 307806
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 176653 306098 176719 306101
rect 176653 306096 179522 306098
rect 176653 306040 176658 306096
rect 176714 306040 179522 306096
rect 176653 306038 179522 306040
rect 176653 306035 176719 306038
rect 179462 306030 179522 306038
rect 179462 305970 180044 306030
rect 294045 305418 294111 305421
rect 292836 305416 294111 305418
rect 292836 305360 294050 305416
rect 294106 305360 294111 305416
rect 292836 305358 294111 305360
rect 294045 305355 294111 305358
rect 179462 303930 180044 303990
rect 177941 303922 178007 303925
rect 179462 303922 179522 303930
rect 177941 303920 179522 303922
rect 177941 303864 177946 303920
rect 178002 303864 179522 303920
rect 177941 303862 179522 303864
rect 177941 303859 178007 303862
rect 295333 303378 295399 303381
rect 292836 303376 295399 303378
rect 292836 303320 295338 303376
rect 295394 303320 295399 303376
rect 292836 303318 295399 303320
rect 295333 303315 295399 303318
rect 109125 302290 109191 302293
rect 110321 302290 110387 302293
rect 161974 302290 161980 302292
rect 109125 302288 161980 302290
rect 109125 302232 109130 302288
rect 109186 302232 110326 302288
rect 110382 302232 161980 302288
rect 109125 302230 161980 302232
rect 109125 302227 109191 302230
rect 110321 302227 110387 302230
rect 161974 302228 161980 302230
rect 162044 302228 162050 302292
rect 295333 301338 295399 301341
rect 292836 301336 295399 301338
rect 292836 301280 295338 301336
rect 295394 301280 295399 301336
rect 292836 301278 295399 301280
rect 295333 301275 295399 301278
rect 179462 301210 180044 301270
rect 176469 301202 176535 301205
rect 179462 301202 179522 301210
rect 176469 301200 179522 301202
rect 176469 301144 176474 301200
rect 176530 301144 179522 301200
rect 176469 301142 179522 301144
rect 176469 301139 176535 301142
rect 70526 300868 70532 300932
rect 70596 300930 70602 300932
rect 142981 300930 143047 300933
rect 70596 300928 143047 300930
rect 70596 300872 142986 300928
rect 143042 300872 143047 300928
rect 70596 300870 143047 300872
rect 70596 300868 70602 300870
rect 142981 300867 143047 300870
rect 110873 299570 110939 299573
rect 111701 299570 111767 299573
rect 124806 299570 124812 299572
rect 110873 299568 124812 299570
rect 110873 299512 110878 299568
rect 110934 299512 111706 299568
rect 111762 299512 124812 299568
rect 110873 299510 124812 299512
rect 110873 299507 110939 299510
rect 111701 299507 111767 299510
rect 124806 299508 124812 299510
rect 124876 299508 124882 299572
rect 176653 299298 176719 299301
rect 294045 299298 294111 299301
rect 176653 299296 179522 299298
rect 176653 299240 176658 299296
rect 176714 299240 179522 299296
rect 176653 299238 179522 299240
rect 292836 299296 294111 299298
rect 292836 299240 294050 299296
rect 294106 299240 294111 299296
rect 292836 299238 294111 299240
rect 176653 299235 176719 299238
rect 179462 299230 179522 299238
rect 294045 299235 294111 299238
rect 377949 299298 378015 299301
rect 379605 299298 379671 299301
rect 377949 299296 380052 299298
rect 377949 299240 377954 299296
rect 378010 299240 379610 299296
rect 379666 299240 380052 299296
rect 377949 299238 380052 299240
rect 377949 299235 378015 299238
rect 379605 299235 379671 299238
rect 179462 299170 180044 299230
rect 60038 298692 60044 298756
rect 60108 298754 60114 298756
rect 121494 298754 121500 298756
rect 60108 298694 121500 298754
rect 60108 298692 60114 298694
rect 121494 298692 121500 298694
rect 121564 298692 121570 298756
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect 104157 298210 104223 298213
rect 156597 298210 156663 298213
rect 104157 298208 156663 298210
rect 104157 298152 104162 298208
rect 104218 298152 156602 298208
rect 156658 298152 156663 298208
rect 104157 298150 156663 298152
rect 104157 298147 104223 298150
rect 156597 298147 156663 298150
rect 112437 297666 112503 297669
rect 117221 297666 117287 297669
rect 112437 297664 117287 297666
rect 112437 297608 112442 297664
rect 112498 297608 117226 297664
rect 117282 297608 117287 297664
rect 112437 297606 117287 297608
rect 112437 297603 112503 297606
rect 117221 297603 117287 297606
rect 65977 297394 66043 297397
rect 164877 297394 164943 297397
rect 65977 297392 164943 297394
rect 65977 297336 65982 297392
rect 66038 297336 164882 297392
rect 164938 297336 164943 297392
rect 65977 297334 164943 297336
rect 65977 297331 66043 297334
rect 164877 297331 164943 297334
rect 179462 297130 180044 297190
rect 176653 297122 176719 297125
rect 179462 297122 179522 297130
rect 176653 297120 179522 297122
rect 176653 297064 176658 297120
rect 176714 297064 179522 297120
rect 176653 297062 179522 297064
rect 376937 297122 377003 297125
rect 442809 297122 442875 297125
rect 376937 297120 380052 297122
rect 376937 297064 376942 297120
rect 376998 297064 380052 297120
rect 376937 297062 380052 297064
rect 439852 297120 442875 297122
rect 439852 297064 442814 297120
rect 442870 297064 442875 297120
rect 439852 297062 442875 297064
rect 176653 297059 176719 297062
rect 376937 297059 377003 297062
rect 442809 297059 442875 297062
rect 116669 296850 116735 296853
rect 124305 296850 124371 296853
rect 116669 296848 124371 296850
rect 116669 296792 116674 296848
rect 116730 296792 124310 296848
rect 124366 296792 124371 296848
rect 116669 296790 124371 296792
rect 116669 296787 116735 296790
rect 124305 296787 124371 296790
rect 295333 296578 295399 296581
rect 292836 296576 295399 296578
rect 292836 296520 295338 296576
rect 295394 296520 295399 296576
rect 292836 296518 295399 296520
rect 295333 296515 295399 296518
rect 80697 296034 80763 296037
rect 97717 296034 97783 296037
rect 80697 296032 97783 296034
rect 80697 295976 80702 296032
rect 80758 295976 97722 296032
rect 97778 295976 97783 296032
rect 80697 295974 97783 295976
rect 80697 295971 80763 295974
rect 97717 295971 97783 295974
rect 106733 295626 106799 295629
rect 119705 295626 119771 295629
rect 106733 295624 119771 295626
rect 106733 295568 106738 295624
rect 106794 295568 119710 295624
rect 119766 295568 119771 295624
rect 106733 295566 119771 295568
rect 106733 295563 106799 295566
rect 119705 295563 119771 295566
rect 97717 295490 97783 295493
rect 165061 295490 165127 295493
rect 97717 295488 165127 295490
rect 97717 295432 97722 295488
rect 97778 295432 165066 295488
rect 165122 295432 165127 295488
rect 97717 295430 165127 295432
rect 97717 295427 97783 295430
rect 165061 295427 165127 295430
rect 71957 295354 72023 295357
rect 73061 295354 73127 295357
rect 146886 295354 146892 295356
rect 71957 295352 146892 295354
rect 71957 295296 71962 295352
rect 72018 295296 73066 295352
rect 73122 295296 146892 295352
rect 71957 295294 146892 295296
rect 71957 295291 72023 295294
rect 73061 295291 73127 295294
rect 146886 295292 146892 295294
rect 146956 295292 146962 295356
rect 379145 295218 379211 295221
rect 379145 295216 380052 295218
rect 379145 295160 379150 295216
rect 379206 295160 380052 295216
rect 379145 295158 380052 295160
rect 379145 295155 379211 295158
rect 179462 295090 180044 295150
rect 176653 295082 176719 295085
rect 179462 295082 179522 295090
rect 441705 295082 441771 295085
rect 442809 295082 442875 295085
rect 176653 295080 179522 295082
rect 176653 295024 176658 295080
rect 176714 295024 179522 295080
rect 176653 295022 179522 295024
rect 439852 295080 442875 295082
rect 439852 295024 441710 295080
rect 441766 295024 442814 295080
rect 442870 295024 442875 295080
rect 439852 295022 442875 295024
rect 176653 295019 176719 295022
rect 441705 295019 441771 295022
rect 442809 295019 442875 295022
rect 296621 294538 296687 294541
rect 292836 294536 296687 294538
rect 292836 294480 296626 294536
rect 296682 294480 296687 294536
rect 292836 294478 296687 294480
rect 296621 294475 296687 294478
rect 75269 294266 75335 294269
rect 75821 294266 75887 294269
rect 173566 294266 173572 294268
rect 75269 294264 173572 294266
rect 75269 294208 75274 294264
rect 75330 294208 75826 294264
rect 75882 294208 173572 294264
rect 75269 294206 173572 294208
rect 75269 294203 75335 294206
rect 75821 294203 75887 294206
rect 173566 294204 173572 294206
rect 173636 294204 173642 294268
rect 117681 294130 117747 294133
rect 171726 294130 171732 294132
rect 117681 294128 171732 294130
rect 117681 294072 117686 294128
rect 117742 294072 171732 294128
rect 117681 294070 171732 294072
rect 117681 294067 117747 294070
rect 171726 294068 171732 294070
rect 171796 294068 171802 294132
rect 117221 293994 117287 293997
rect 118969 293994 119035 293997
rect 119654 293994 119660 293996
rect 117221 293992 119660 293994
rect 117221 293936 117226 293992
rect 117282 293936 118974 293992
rect 119030 293936 119660 293992
rect 117221 293934 119660 293936
rect 117221 293931 117287 293934
rect 118969 293931 119035 293934
rect 119654 293932 119660 293934
rect 119724 293932 119730 293996
rect 168281 293994 168347 293997
rect 170254 293994 170260 293996
rect 168281 293992 170260 293994
rect 168281 293936 168286 293992
rect 168342 293936 170260 293992
rect 168281 293934 170260 293936
rect 168281 293931 168347 293934
rect 170254 293932 170260 293934
rect 170324 293932 170330 293996
rect -960 293178 480 293268
rect 3233 293178 3299 293181
rect -960 293176 3299 293178
rect -960 293120 3238 293176
rect 3294 293120 3299 293176
rect -960 293118 3299 293120
rect -960 293028 480 293118
rect 3233 293115 3299 293118
rect 377397 293042 377463 293045
rect 443177 293042 443243 293045
rect 377397 293040 380052 293042
rect 377397 292984 377402 293040
rect 377458 292984 380052 293040
rect 377397 292982 380052 292984
rect 439852 293040 443243 293042
rect 439852 292984 443182 293040
rect 443238 292984 443243 293040
rect 439852 292982 443243 292984
rect 377397 292979 377463 292982
rect 443177 292979 443243 292982
rect 77753 292770 77819 292773
rect 126094 292770 126100 292772
rect 77753 292768 126100 292770
rect 77753 292712 77758 292768
rect 77814 292712 126100 292768
rect 77753 292710 126100 292712
rect 77753 292707 77819 292710
rect 126094 292708 126100 292710
rect 126164 292708 126170 292772
rect 92565 292634 92631 292637
rect 166257 292634 166323 292637
rect 92565 292632 166323 292634
rect 92565 292576 92570 292632
rect 92626 292576 166262 292632
rect 166318 292576 166323 292632
rect 92565 292574 166323 292576
rect 92565 292571 92631 292574
rect 166257 292571 166323 292574
rect 295333 292498 295399 292501
rect 292836 292496 295399 292498
rect 292836 292440 295338 292496
rect 295394 292440 295399 292496
rect 292836 292438 295399 292440
rect 295333 292435 295399 292438
rect 179462 292370 180044 292430
rect 179229 292362 179295 292365
rect 179462 292362 179522 292370
rect 179229 292360 179522 292362
rect 179229 292304 179234 292360
rect 179290 292304 179522 292360
rect 179229 292302 179522 292304
rect 179229 292299 179295 292302
rect 117221 292090 117287 292093
rect 160686 292090 160692 292092
rect 117221 292088 160692 292090
rect 117221 292032 117226 292088
rect 117282 292032 160692 292088
rect 117221 292030 160692 292032
rect 117221 292027 117287 292030
rect 160686 292028 160692 292030
rect 160756 292028 160762 292092
rect 118601 291954 118667 291957
rect 118601 291952 119354 291954
rect 118601 291896 118606 291952
rect 118662 291896 119354 291952
rect 118601 291894 119354 291896
rect 118601 291891 118667 291894
rect 68277 291818 68343 291821
rect 68277 291816 70196 291818
rect 68277 291760 68282 291816
rect 68338 291760 70196 291816
rect 119294 291788 119354 291894
rect 120022 291892 120028 291956
rect 120092 291954 120098 291956
rect 120165 291954 120231 291957
rect 120092 291952 120231 291954
rect 120092 291896 120170 291952
rect 120226 291896 120231 291952
rect 120092 291894 120231 291896
rect 120092 291892 120098 291894
rect 120165 291891 120231 291894
rect 305545 291818 305611 291821
rect 376150 291818 376156 291820
rect 305545 291816 376156 291818
rect 68277 291758 70196 291760
rect 305545 291760 305550 291816
rect 305606 291760 376156 291816
rect 305545 291758 376156 291760
rect 68277 291755 68343 291758
rect 305545 291755 305611 291758
rect 376150 291756 376156 291758
rect 376220 291756 376226 291820
rect 67725 291138 67791 291141
rect 121545 291138 121611 291141
rect 440325 291138 440391 291141
rect 67725 291136 70196 291138
rect 67725 291080 67730 291136
rect 67786 291080 70196 291136
rect 67725 291078 70196 291080
rect 119876 291136 121611 291138
rect 119876 291080 121550 291136
rect 121606 291080 121611 291136
rect 119876 291078 121611 291080
rect 439852 291136 440391 291138
rect 439852 291080 440330 291136
rect 440386 291080 440391 291136
rect 439852 291078 440391 291080
rect 67725 291075 67791 291078
rect 121545 291075 121611 291078
rect 440325 291075 440391 291078
rect 376937 291002 377003 291005
rect 376937 291000 380052 291002
rect 376937 290944 376942 291000
rect 376998 290944 380052 291000
rect 376937 290942 380052 290944
rect 376937 290939 377003 290942
rect 68921 290866 68987 290869
rect 70526 290866 70532 290868
rect 68921 290864 70532 290866
rect 68921 290808 68926 290864
rect 68982 290808 70532 290864
rect 68921 290806 70532 290808
rect 68921 290803 68987 290806
rect 70526 290804 70532 290806
rect 70596 290804 70602 290868
rect 67633 290458 67699 290461
rect 121637 290458 121703 290461
rect 67633 290456 70196 290458
rect 67633 290400 67638 290456
rect 67694 290400 70196 290456
rect 67633 290398 70196 290400
rect 119876 290456 121703 290458
rect 119876 290400 121642 290456
rect 121698 290400 121703 290456
rect 119876 290398 121703 290400
rect 67633 290395 67699 290398
rect 121637 290395 121703 290398
rect 176653 290458 176719 290461
rect 295333 290458 295399 290461
rect 176653 290456 179522 290458
rect 176653 290400 176658 290456
rect 176714 290400 179522 290456
rect 176653 290398 179522 290400
rect 292836 290456 295399 290458
rect 292836 290400 295338 290456
rect 295394 290400 295399 290456
rect 292836 290398 295399 290400
rect 176653 290395 176719 290398
rect 179462 290390 179522 290398
rect 295333 290395 295399 290398
rect 179462 290330 180044 290390
rect 67725 289778 67791 289781
rect 121545 289778 121611 289781
rect 67725 289776 70196 289778
rect 67725 289720 67730 289776
rect 67786 289720 70196 289776
rect 67725 289718 70196 289720
rect 119876 289776 121611 289778
rect 119876 289720 121550 289776
rect 121606 289720 121611 289776
rect 119876 289718 121611 289720
rect 67725 289715 67791 289718
rect 121545 289715 121611 289718
rect 439446 289580 439452 289644
rect 439516 289580 439522 289644
rect 67633 289098 67699 289101
rect 121637 289098 121703 289101
rect 67633 289096 70196 289098
rect 67633 289040 67638 289096
rect 67694 289040 70196 289096
rect 67633 289038 70196 289040
rect 119876 289096 121703 289098
rect 119876 289040 121642 289096
rect 121698 289040 121703 289096
rect 119876 289038 121703 289040
rect 67633 289035 67699 289038
rect 121637 289035 121703 289038
rect 135161 289098 135227 289101
rect 167678 289098 167684 289100
rect 135161 289096 167684 289098
rect 135161 289040 135166 289096
rect 135222 289040 167684 289096
rect 135161 289038 167684 289040
rect 135161 289035 135227 289038
rect 167678 289036 167684 289038
rect 167748 289036 167754 289100
rect 376937 288962 377003 288965
rect 376937 288960 380052 288962
rect 376937 288904 376942 288960
rect 376998 288904 380052 288960
rect 376937 288902 380052 288904
rect 376937 288899 377003 288902
rect 439454 288826 439514 289580
rect 440417 288826 440483 288829
rect 439454 288824 440483 288826
rect 439454 288768 440422 288824
rect 440478 288768 440483 288824
rect 439454 288766 440483 288768
rect 440417 288763 440483 288766
rect 69105 288418 69171 288421
rect 69105 288416 70196 288418
rect 69105 288360 69110 288416
rect 69166 288360 70196 288416
rect 69105 288358 70196 288360
rect 69105 288355 69171 288358
rect 119846 287874 119906 288388
rect 179462 288290 180044 288350
rect 176653 288282 176719 288285
rect 179462 288282 179522 288290
rect 176653 288280 179522 288282
rect 176653 288224 176658 288280
rect 176714 288224 179522 288280
rect 176653 288222 179522 288224
rect 176653 288219 176719 288222
rect 119846 287814 122850 287874
rect 67633 287738 67699 287741
rect 121545 287738 121611 287741
rect 67633 287736 70196 287738
rect 67633 287680 67638 287736
rect 67694 287680 70196 287736
rect 67633 287678 70196 287680
rect 119876 287736 121611 287738
rect 119876 287680 121550 287736
rect 121606 287680 121611 287736
rect 119876 287678 121611 287680
rect 67633 287675 67699 287678
rect 121545 287675 121611 287678
rect 122790 287194 122850 287814
rect 157374 287194 157380 287196
rect 122790 287134 157380 287194
rect 157374 287132 157380 287134
rect 157444 287132 157450 287196
rect 292806 287194 292866 287708
rect 296161 287196 296227 287197
rect 293902 287194 293908 287196
rect 292806 287134 293908 287194
rect 293902 287132 293908 287134
rect 293972 287194 293978 287196
rect 296110 287194 296116 287196
rect 293972 287134 296116 287194
rect 296180 287194 296227 287196
rect 296180 287192 296272 287194
rect 296222 287136 296272 287192
rect 293972 287132 293978 287134
rect 296110 287132 296116 287134
rect 296180 287134 296272 287136
rect 296180 287132 296227 287134
rect 296161 287131 296227 287132
rect 67725 287058 67791 287061
rect 121729 287058 121795 287061
rect 440969 287058 441035 287061
rect 441521 287058 441587 287061
rect 67725 287056 70196 287058
rect 67725 287000 67730 287056
rect 67786 287000 70196 287056
rect 67725 286998 70196 287000
rect 119876 287056 121795 287058
rect 119876 287000 121734 287056
rect 121790 287000 121795 287056
rect 119876 286998 121795 287000
rect 439852 287056 441587 287058
rect 439852 287000 440974 287056
rect 441030 287000 441526 287056
rect 441582 287000 441587 287056
rect 439852 286998 441587 287000
rect 67725 286995 67791 286998
rect 121729 286995 121795 286998
rect 440969 286995 441035 286998
rect 441521 286995 441587 286998
rect 376937 286922 377003 286925
rect 376937 286920 380052 286922
rect 376937 286864 376942 286920
rect 376998 286864 380052 286920
rect 376937 286862 380052 286864
rect 376937 286859 377003 286862
rect 68921 286378 68987 286381
rect 120257 286378 120323 286381
rect 295926 286378 295932 286380
rect 68921 286376 70196 286378
rect 68921 286320 68926 286376
rect 68982 286320 70196 286376
rect 68921 286318 70196 286320
rect 119876 286376 120323 286378
rect 119876 286320 120262 286376
rect 120318 286320 120323 286376
rect 119876 286318 120323 286320
rect 68921 286315 68987 286318
rect 120257 286315 120323 286318
rect 292806 286318 295932 286378
rect 179462 286250 180044 286310
rect 177297 286242 177363 286245
rect 179462 286242 179522 286250
rect 177297 286240 179522 286242
rect 177297 286184 177302 286240
rect 177358 286184 179522 286240
rect 177297 286182 179522 286184
rect 177297 286179 177363 286182
rect 68737 285698 68803 285701
rect 122741 285698 122807 285701
rect 68737 285696 70196 285698
rect 68737 285640 68742 285696
rect 68798 285640 70196 285696
rect 68737 285638 70196 285640
rect 119876 285696 122807 285698
rect 119876 285640 122746 285696
rect 122802 285640 122807 285696
rect 292806 285668 292866 286318
rect 295926 286316 295932 286318
rect 295996 286378 296002 286380
rect 373206 286378 373212 286380
rect 295996 286318 373212 286378
rect 295996 286316 296002 286318
rect 373206 286316 373212 286318
rect 373276 286316 373282 286380
rect 119876 285638 122807 285640
rect 68737 285635 68803 285638
rect 122741 285635 122807 285638
rect 583520 285276 584960 285516
rect 68645 285018 68711 285021
rect 122465 285018 122531 285021
rect 442165 285018 442231 285021
rect 68645 285016 70196 285018
rect 68645 284960 68650 285016
rect 68706 284960 70196 285016
rect 68645 284958 70196 284960
rect 119876 285016 122531 285018
rect 119876 284960 122470 285016
rect 122526 284960 122531 285016
rect 119876 284958 122531 284960
rect 439852 285016 442231 285018
rect 439852 284960 442170 285016
rect 442226 284960 442231 285016
rect 439852 284958 442231 284960
rect 68645 284955 68711 284958
rect 122465 284955 122531 284958
rect 442165 284955 442231 284958
rect 55622 284820 55628 284884
rect 55692 284882 55698 284884
rect 68001 284882 68067 284885
rect 55692 284880 68067 284882
rect 55692 284824 68006 284880
rect 68062 284824 68067 284880
rect 55692 284822 68067 284824
rect 55692 284820 55698 284822
rect 68001 284819 68067 284822
rect 120574 284820 120580 284884
rect 120644 284882 120650 284884
rect 138606 284882 138612 284884
rect 120644 284822 138612 284882
rect 120644 284820 120650 284822
rect 138606 284820 138612 284822
rect 138676 284820 138682 284884
rect 67633 284338 67699 284341
rect 121453 284338 121519 284341
rect 67633 284336 70196 284338
rect 67633 284280 67638 284336
rect 67694 284280 70196 284336
rect 67633 284278 70196 284280
rect 119876 284336 121519 284338
rect 119876 284280 121458 284336
rect 121514 284280 121519 284336
rect 119876 284278 121519 284280
rect 67633 284275 67699 284278
rect 121453 284275 121519 284278
rect 377305 284202 377371 284205
rect 377305 284200 380052 284202
rect 377305 284144 377310 284200
rect 377366 284144 380052 284200
rect 377305 284142 380052 284144
rect 377305 284139 377371 284142
rect 68001 283658 68067 283661
rect 68921 283658 68987 283661
rect 121453 283658 121519 283661
rect 68001 283656 70196 283658
rect 68001 283600 68006 283656
rect 68062 283600 68926 283656
rect 68982 283600 70196 283656
rect 68001 283598 70196 283600
rect 119876 283656 121519 283658
rect 119876 283600 121458 283656
rect 121514 283600 121519 283656
rect 119876 283598 121519 283600
rect 68001 283595 68067 283598
rect 68921 283595 68987 283598
rect 121453 283595 121519 283598
rect 176653 283658 176719 283661
rect 294781 283658 294847 283661
rect 295241 283658 295307 283661
rect 176653 283656 179522 283658
rect 176653 283600 176658 283656
rect 176714 283600 179522 283656
rect 176653 283598 179522 283600
rect 292836 283656 295307 283658
rect 292836 283600 294786 283656
rect 294842 283600 295246 283656
rect 295302 283600 295307 283656
rect 292836 283598 295307 283600
rect 176653 283595 176719 283598
rect 179462 283590 179522 283598
rect 294781 283595 294847 283598
rect 295241 283595 295307 283598
rect 179462 283530 180044 283590
rect 126094 283460 126100 283524
rect 126164 283522 126170 283524
rect 154389 283522 154455 283525
rect 158621 283522 158687 283525
rect 126164 283520 158687 283522
rect 126164 283464 154394 283520
rect 154450 283464 158626 283520
rect 158682 283464 158687 283520
rect 126164 283462 158687 283464
rect 126164 283460 126170 283462
rect 154389 283459 154455 283462
rect 158621 283459 158687 283462
rect 67725 282978 67791 282981
rect 122741 282978 122807 282981
rect 67725 282976 70196 282978
rect 67725 282920 67730 282976
rect 67786 282920 70196 282976
rect 67725 282918 70196 282920
rect 119876 282976 122807 282978
rect 119876 282920 122746 282976
rect 122802 282920 122807 282976
rect 119876 282918 122807 282920
rect 67725 282915 67791 282918
rect 122741 282915 122807 282918
rect 121545 282298 121611 282301
rect 119876 282296 121611 282298
rect 119876 282240 121550 282296
rect 121606 282240 121611 282296
rect 119876 282238 121611 282240
rect 121545 282235 121611 282238
rect 376937 282162 377003 282165
rect 442717 282162 442783 282165
rect 376937 282160 380052 282162
rect 376937 282104 376942 282160
rect 376998 282104 380052 282160
rect 376937 282102 380052 282104
rect 439852 282160 442783 282162
rect 439852 282104 442722 282160
rect 442778 282104 442783 282160
rect 439852 282102 442783 282104
rect 376937 282099 377003 282102
rect 442717 282099 442783 282102
rect 68553 281618 68619 281621
rect 121453 281618 121519 281621
rect 68553 281616 70196 281618
rect 68553 281560 68558 281616
rect 68614 281560 70196 281616
rect 68553 281558 70196 281560
rect 119876 281616 121519 281618
rect 119876 281560 121458 281616
rect 121514 281560 121519 281616
rect 119876 281558 121519 281560
rect 68553 281555 68619 281558
rect 121453 281555 121519 281558
rect 176653 281618 176719 281621
rect 295333 281618 295399 281621
rect 176653 281616 179522 281618
rect 176653 281560 176658 281616
rect 176714 281560 179522 281616
rect 176653 281558 179522 281560
rect 292836 281616 295399 281618
rect 292836 281560 295338 281616
rect 295394 281560 295399 281616
rect 292836 281558 295399 281560
rect 176653 281555 176719 281558
rect 179462 281550 179522 281558
rect 295333 281555 295399 281558
rect 179462 281490 180044 281550
rect 67633 280938 67699 280941
rect 121361 280938 121427 280941
rect 121494 280938 121500 280940
rect 67633 280936 70196 280938
rect 67633 280880 67638 280936
rect 67694 280880 70196 280936
rect 67633 280878 70196 280880
rect 119876 280936 121500 280938
rect 119876 280880 121366 280936
rect 121422 280880 121500 280936
rect 119876 280878 121500 280880
rect 67633 280875 67699 280878
rect 121361 280875 121427 280878
rect 121494 280876 121500 280878
rect 121564 280876 121570 280940
rect 67633 280258 67699 280261
rect 121453 280258 121519 280261
rect 67633 280256 70196 280258
rect -960 279972 480 280212
rect 67633 280200 67638 280256
rect 67694 280200 70196 280256
rect 67633 280198 70196 280200
rect 119876 280256 121519 280258
rect 119876 280200 121458 280256
rect 121514 280200 121519 280256
rect 119876 280198 121519 280200
rect 67633 280195 67699 280198
rect 121453 280195 121519 280198
rect 376937 280258 377003 280261
rect 442809 280258 442875 280261
rect 376937 280256 380052 280258
rect 376937 280200 376942 280256
rect 376998 280200 380052 280256
rect 376937 280198 380052 280200
rect 439852 280256 442875 280258
rect 439852 280200 442814 280256
rect 442870 280200 442875 280256
rect 439852 280198 442875 280200
rect 376937 280195 377003 280198
rect 442809 280195 442875 280198
rect 67633 279578 67699 279581
rect 122649 279578 122715 279581
rect 67633 279576 70196 279578
rect 67633 279520 67638 279576
rect 67694 279520 70196 279576
rect 67633 279518 70196 279520
rect 119876 279576 122715 279578
rect 119876 279520 122654 279576
rect 122710 279520 122715 279576
rect 119876 279518 122715 279520
rect 67633 279515 67699 279518
rect 122649 279515 122715 279518
rect 176653 279578 176719 279581
rect 176653 279576 179522 279578
rect 176653 279520 176658 279576
rect 176714 279520 179522 279576
rect 176653 279518 179522 279520
rect 176653 279515 176719 279518
rect 179462 279510 179522 279518
rect 179462 279450 180044 279510
rect 67357 278898 67423 278901
rect 121453 278898 121519 278901
rect 296529 278898 296595 278901
rect 297214 278898 297220 278900
rect 67357 278896 70196 278898
rect 67357 278840 67362 278896
rect 67418 278840 70196 278896
rect 67357 278838 70196 278840
rect 119876 278896 121519 278898
rect 119876 278840 121458 278896
rect 121514 278840 121519 278896
rect 119876 278838 121519 278840
rect 292836 278896 297220 278898
rect 292836 278840 296534 278896
rect 296590 278840 297220 278896
rect 292836 278838 297220 278840
rect 67357 278835 67423 278838
rect 121453 278835 121519 278838
rect 296529 278835 296595 278838
rect 297214 278836 297220 278838
rect 297284 278836 297290 278900
rect 67633 278218 67699 278221
rect 120073 278218 120139 278221
rect 122465 278218 122531 278221
rect 67633 278216 70196 278218
rect 67633 278160 67638 278216
rect 67694 278160 70196 278216
rect 67633 278158 70196 278160
rect 119876 278216 122531 278218
rect 119876 278160 120078 278216
rect 120134 278160 122470 278216
rect 122526 278160 122531 278216
rect 119876 278158 122531 278160
rect 67633 278155 67699 278158
rect 120073 278155 120139 278158
rect 122465 278155 122531 278158
rect 376753 278082 376819 278085
rect 442625 278082 442691 278085
rect 376753 278080 380052 278082
rect 376753 278024 376758 278080
rect 376814 278024 380052 278080
rect 376753 278022 380052 278024
rect 439852 278080 442691 278082
rect 439852 278024 442630 278080
rect 442686 278024 442691 278080
rect 439852 278022 442691 278024
rect 376753 278019 376819 278022
rect 442625 278019 442691 278022
rect 67633 277538 67699 277541
rect 121545 277538 121611 277541
rect 67633 277536 70196 277538
rect 67633 277480 67638 277536
rect 67694 277480 70196 277536
rect 67633 277478 70196 277480
rect 119876 277536 121611 277538
rect 119876 277480 121550 277536
rect 121606 277480 121611 277536
rect 119876 277478 121611 277480
rect 67633 277475 67699 277478
rect 121545 277475 121611 277478
rect 176653 277538 176719 277541
rect 176653 277536 179522 277538
rect 176653 277480 176658 277536
rect 176714 277480 179522 277536
rect 176653 277478 179522 277480
rect 176653 277475 176719 277478
rect 179462 277470 179522 277478
rect 179462 277410 180044 277470
rect 293033 276994 293099 276997
rect 292806 276992 293099 276994
rect 292806 276936 293038 276992
rect 293094 276936 293099 276992
rect 292806 276934 293099 276936
rect 67725 276858 67791 276861
rect 121453 276858 121519 276861
rect 67725 276856 70196 276858
rect 67725 276800 67730 276856
rect 67786 276800 70196 276856
rect 67725 276798 70196 276800
rect 119876 276856 121519 276858
rect 119876 276800 121458 276856
rect 121514 276800 121519 276856
rect 292806 276828 292866 276934
rect 293033 276931 293099 276934
rect 119876 276798 121519 276800
rect 67725 276795 67791 276798
rect 121453 276795 121519 276798
rect 67633 276178 67699 276181
rect 121453 276178 121519 276181
rect 67633 276176 70196 276178
rect 67633 276120 67638 276176
rect 67694 276120 70196 276176
rect 67633 276118 70196 276120
rect 119876 276176 121519 276178
rect 119876 276120 121458 276176
rect 121514 276120 121519 276176
rect 119876 276118 121519 276120
rect 67633 276115 67699 276118
rect 121453 276115 121519 276118
rect 377765 276042 377831 276045
rect 379513 276042 379579 276045
rect 440325 276042 440391 276045
rect 440877 276042 440943 276045
rect 377765 276040 380052 276042
rect 377765 275984 377770 276040
rect 377826 275984 379518 276040
rect 379574 275984 380052 276040
rect 377765 275982 380052 275984
rect 439852 276040 440943 276042
rect 439852 275984 440330 276040
rect 440386 275984 440882 276040
rect 440938 275984 440943 276040
rect 439852 275982 440943 275984
rect 377765 275979 377831 275982
rect 379513 275979 379579 275982
rect 440325 275979 440391 275982
rect 440877 275979 440943 275982
rect 54334 275844 54340 275908
rect 54404 275906 54410 275908
rect 54845 275906 54911 275909
rect 54404 275904 54911 275906
rect 54404 275848 54850 275904
rect 54906 275848 54911 275904
rect 54404 275846 54911 275848
rect 54404 275844 54410 275846
rect 54845 275843 54911 275846
rect 67633 275498 67699 275501
rect 121453 275498 121519 275501
rect 67633 275496 70196 275498
rect 67633 275440 67638 275496
rect 67694 275440 70196 275496
rect 67633 275438 70196 275440
rect 119876 275496 121519 275498
rect 119876 275440 121458 275496
rect 121514 275440 121519 275496
rect 119876 275438 121519 275440
rect 67633 275435 67699 275438
rect 121453 275435 121519 275438
rect 68277 274818 68343 274821
rect 121545 274818 121611 274821
rect 68277 274816 70196 274818
rect 68277 274760 68282 274816
rect 68338 274760 70196 274816
rect 68277 274758 70196 274760
rect 119876 274816 121611 274818
rect 119876 274760 121550 274816
rect 121606 274760 121611 274816
rect 119876 274758 121611 274760
rect 68277 274755 68343 274758
rect 121545 274755 121611 274758
rect 176653 274818 176719 274821
rect 295333 274818 295399 274821
rect 176653 274816 179522 274818
rect 176653 274760 176658 274816
rect 176714 274760 179522 274816
rect 176653 274758 179522 274760
rect 292836 274816 295399 274818
rect 292836 274760 295338 274816
rect 295394 274760 295399 274816
rect 292836 274758 295399 274760
rect 176653 274755 176719 274758
rect 179462 274750 179522 274758
rect 295333 274755 295399 274758
rect 179462 274690 180044 274750
rect 67633 274138 67699 274141
rect 121453 274138 121519 274141
rect 67633 274136 70196 274138
rect 67633 274080 67638 274136
rect 67694 274080 70196 274136
rect 67633 274078 70196 274080
rect 119876 274136 121519 274138
rect 119876 274080 121458 274136
rect 121514 274080 121519 274136
rect 119876 274078 121519 274080
rect 67633 274075 67699 274078
rect 121453 274075 121519 274078
rect 377765 274002 377831 274005
rect 379421 274002 379487 274005
rect 442717 274002 442783 274005
rect 377765 274000 380052 274002
rect 377765 273944 377770 274000
rect 377826 273944 379426 274000
rect 379482 273944 380052 274000
rect 377765 273942 380052 273944
rect 439852 274000 442783 274002
rect 439852 273944 442722 274000
rect 442778 273944 442783 274000
rect 439852 273942 442783 273944
rect 377765 273939 377831 273942
rect 379421 273939 379487 273942
rect 442717 273939 442783 273942
rect 67817 273458 67883 273461
rect 121453 273458 121519 273461
rect 67817 273456 70196 273458
rect 67817 273400 67822 273456
rect 67878 273400 70196 273456
rect 67817 273398 70196 273400
rect 119876 273456 121519 273458
rect 119876 273400 121458 273456
rect 121514 273400 121519 273456
rect 119876 273398 121519 273400
rect 67817 273395 67883 273398
rect 121453 273395 121519 273398
rect 67633 272778 67699 272781
rect 121453 272778 121519 272781
rect 295333 272778 295399 272781
rect 67633 272776 70196 272778
rect 67633 272720 67638 272776
rect 67694 272720 70196 272776
rect 67633 272718 70196 272720
rect 119876 272776 121519 272778
rect 119876 272720 121458 272776
rect 121514 272720 121519 272776
rect 119876 272718 121519 272720
rect 292836 272776 295399 272778
rect 292836 272720 295338 272776
rect 295394 272720 295399 272776
rect 292836 272718 295399 272720
rect 67633 272715 67699 272718
rect 121453 272715 121519 272718
rect 295333 272715 295399 272718
rect 179462 272650 180044 272710
rect 176653 272642 176719 272645
rect 179462 272642 179522 272650
rect 176653 272640 179522 272642
rect 176653 272584 176658 272640
rect 176714 272584 179522 272640
rect 176653 272582 179522 272584
rect 176653 272579 176719 272582
rect 582373 272234 582439 272237
rect 583520 272234 584960 272324
rect 582373 272232 584960 272234
rect 582373 272176 582378 272232
rect 582434 272176 584960 272232
rect 582373 272174 584960 272176
rect 582373 272171 582439 272174
rect 67449 272098 67515 272101
rect 122189 272098 122255 272101
rect 67449 272096 70196 272098
rect 67449 272040 67454 272096
rect 67510 272040 70196 272096
rect 67449 272038 70196 272040
rect 119876 272096 122255 272098
rect 119876 272040 122194 272096
rect 122250 272040 122255 272096
rect 119876 272038 122255 272040
rect 67449 272035 67515 272038
rect 122189 272035 122255 272038
rect 378869 272098 378935 272101
rect 379237 272098 379303 272101
rect 442809 272098 442875 272101
rect 378869 272096 380052 272098
rect 378869 272040 378874 272096
rect 378930 272040 379242 272096
rect 379298 272040 380052 272096
rect 378869 272038 380052 272040
rect 439852 272096 442875 272098
rect 439852 272040 442814 272096
rect 442870 272040 442875 272096
rect 583520 272084 584960 272174
rect 439852 272038 442875 272040
rect 378869 272035 378935 272038
rect 379237 272035 379303 272038
rect 442809 272035 442875 272038
rect 67725 271418 67791 271421
rect 121453 271418 121519 271421
rect 67725 271416 70196 271418
rect 67725 271360 67730 271416
rect 67786 271360 70196 271416
rect 67725 271358 70196 271360
rect 119876 271416 121519 271418
rect 119876 271360 121458 271416
rect 121514 271360 121519 271416
rect 119876 271358 121519 271360
rect 67725 271355 67791 271358
rect 121453 271355 121519 271358
rect 67633 270738 67699 270741
rect 67633 270736 70196 270738
rect 67633 270680 67638 270736
rect 67694 270680 70196 270736
rect 67633 270678 70196 270680
rect 67633 270675 67699 270678
rect 179689 270670 179755 270673
rect 179462 270668 180044 270670
rect 179462 270612 179694 270668
rect 179750 270612 180044 270668
rect 179462 270610 180044 270612
rect 179462 270605 179522 270610
rect 179689 270607 179755 270610
rect 179413 270600 179522 270605
rect 179413 270544 179418 270600
rect 179474 270544 179522 270600
rect 179413 270542 179522 270544
rect 179413 270539 179479 270542
rect 295926 270466 295932 270468
rect 292806 270406 295932 270466
rect 67633 270058 67699 270061
rect 121453 270058 121519 270061
rect 67633 270056 70196 270058
rect 67633 270000 67638 270056
rect 67694 270000 70196 270056
rect 67633 269998 70196 270000
rect 119876 270056 121519 270058
rect 119876 270000 121458 270056
rect 121514 270000 121519 270056
rect 292806 270028 292866 270406
rect 295926 270404 295932 270406
rect 295996 270466 296002 270468
rect 296069 270466 296135 270469
rect 295996 270464 296135 270466
rect 295996 270408 296074 270464
rect 296130 270408 296135 270464
rect 295996 270406 296135 270408
rect 295996 270404 296002 270406
rect 296069 270403 296135 270406
rect 119876 269998 121519 270000
rect 67633 269995 67699 269998
rect 121453 269995 121519 269998
rect 442257 269922 442323 269925
rect 439852 269920 442323 269922
rect 439852 269864 442262 269920
rect 442318 269864 442323 269920
rect 439852 269862 442323 269864
rect 442257 269859 442323 269862
rect 67725 269378 67791 269381
rect 121545 269378 121611 269381
rect 67725 269376 70196 269378
rect 67725 269320 67730 269376
rect 67786 269320 70196 269376
rect 67725 269318 70196 269320
rect 119876 269376 121611 269378
rect 119876 269320 121550 269376
rect 121606 269320 121611 269376
rect 119876 269318 121611 269320
rect 67725 269315 67791 269318
rect 121545 269315 121611 269318
rect 120758 269180 120764 269244
rect 120828 269242 120834 269244
rect 165521 269242 165587 269245
rect 120828 269240 165587 269242
rect 120828 269184 165526 269240
rect 165582 269184 165587 269240
rect 120828 269182 165587 269184
rect 120828 269180 120834 269182
rect 165521 269179 165587 269182
rect 378726 269180 378732 269244
rect 378796 269242 378802 269244
rect 378796 269182 380052 269242
rect 378796 269180 378802 269182
rect 67725 268698 67791 268701
rect 121453 268698 121519 268701
rect 67725 268696 70196 268698
rect 67725 268640 67730 268696
rect 67786 268640 70196 268696
rect 67725 268638 70196 268640
rect 119876 268696 121519 268698
rect 119876 268640 121458 268696
rect 121514 268640 121519 268696
rect 119876 268638 121519 268640
rect 67725 268635 67791 268638
rect 121453 268635 121519 268638
rect 179462 268570 180044 268630
rect 176653 268562 176719 268565
rect 179462 268562 179522 268570
rect 176653 268560 179522 268562
rect 176653 268504 176658 268560
rect 176714 268504 179522 268560
rect 176653 268502 179522 268504
rect 176653 268499 176719 268502
rect 67633 268018 67699 268021
rect 121453 268018 121519 268021
rect 294229 268018 294295 268021
rect 67633 268016 70196 268018
rect 67633 267960 67638 268016
rect 67694 267960 70196 268016
rect 67633 267958 70196 267960
rect 119876 268016 121519 268018
rect 119876 267960 121458 268016
rect 121514 267960 121519 268016
rect 119876 267958 121519 267960
rect 292836 268016 294295 268018
rect 292836 267960 294234 268016
rect 294290 267960 294295 268016
rect 292836 267958 294295 267960
rect 67633 267955 67699 267958
rect 121453 267955 121519 267958
rect 294229 267955 294295 267958
rect 67633 267338 67699 267341
rect 122281 267338 122347 267341
rect 67633 267336 70196 267338
rect -960 267202 480 267292
rect 67633 267280 67638 267336
rect 67694 267280 70196 267336
rect 67633 267278 70196 267280
rect 119876 267336 122347 267338
rect 119876 267280 122286 267336
rect 122342 267280 122347 267336
rect 119876 267278 122347 267280
rect 67633 267275 67699 267278
rect 122281 267275 122347 267278
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 379237 267202 379303 267205
rect 442809 267202 442875 267205
rect 379237 267200 380052 267202
rect 379237 267144 379242 267200
rect 379298 267144 380052 267200
rect 379237 267142 380052 267144
rect 439852 267200 442875 267202
rect 439852 267144 442814 267200
rect 442870 267144 442875 267200
rect 439852 267142 442875 267144
rect 379237 267139 379303 267142
rect 442809 267139 442875 267142
rect 67725 266658 67791 266661
rect 122097 266658 122163 266661
rect 67725 266656 70196 266658
rect 67725 266600 67730 266656
rect 67786 266600 70196 266656
rect 67725 266598 70196 266600
rect 119876 266656 122163 266658
rect 119876 266600 122102 266656
rect 122158 266600 122163 266656
rect 119876 266598 122163 266600
rect 67725 266595 67791 266598
rect 122097 266595 122163 266598
rect 121637 265978 121703 265981
rect 119876 265976 121703 265978
rect 69013 265434 69079 265437
rect 70166 265434 70226 265948
rect 119876 265920 121642 265976
rect 121698 265920 121703 265976
rect 119876 265918 121703 265920
rect 121637 265915 121703 265918
rect 176653 265978 176719 265981
rect 176653 265976 179522 265978
rect 176653 265920 176658 265976
rect 176714 265920 179522 265976
rect 176653 265918 179522 265920
rect 176653 265915 176719 265918
rect 179462 265910 179522 265918
rect 179462 265850 180044 265910
rect 64830 265432 70226 265434
rect 64830 265376 69018 265432
rect 69074 265376 70226 265432
rect 64830 265374 70226 265376
rect 63166 265100 63172 265164
rect 63236 265162 63242 265164
rect 64830 265162 64890 265374
rect 69013 265371 69079 265374
rect 67633 265298 67699 265301
rect 121453 265298 121519 265301
rect 67633 265296 70196 265298
rect 67633 265240 67638 265296
rect 67694 265240 70196 265296
rect 67633 265238 70196 265240
rect 119876 265296 121519 265298
rect 119876 265240 121458 265296
rect 121514 265240 121519 265296
rect 119876 265238 121519 265240
rect 292806 265298 292866 265948
rect 292806 265238 296730 265298
rect 67633 265235 67699 265238
rect 121453 265235 121519 265238
rect 63236 265102 64890 265162
rect 63236 265100 63242 265102
rect 296670 265026 296730 265238
rect 376937 265162 377003 265165
rect 442349 265162 442415 265165
rect 376937 265160 380052 265162
rect 376937 265104 376942 265160
rect 376998 265104 380052 265160
rect 376937 265102 380052 265104
rect 439852 265160 442415 265162
rect 439852 265104 442354 265160
rect 442410 265104 442415 265160
rect 439852 265102 442415 265104
rect 376937 265099 377003 265102
rect 442349 265099 442415 265102
rect 341374 265026 341380 265028
rect 296670 264966 341380 265026
rect 341374 264964 341380 264966
rect 341444 264964 341450 265028
rect 67725 264618 67791 264621
rect 122465 264618 122531 264621
rect 67725 264616 70196 264618
rect 67725 264560 67730 264616
rect 67786 264560 70196 264616
rect 67725 264558 70196 264560
rect 119876 264616 122531 264618
rect 119876 264560 122470 264616
rect 122526 264560 122531 264616
rect 119876 264558 122531 264560
rect 67725 264555 67791 264558
rect 122465 264555 122531 264558
rect 67633 263938 67699 263941
rect 121453 263938 121519 263941
rect 67633 263936 70196 263938
rect 67633 263880 67638 263936
rect 67694 263880 70196 263936
rect 67633 263878 70196 263880
rect 119876 263936 121519 263938
rect 119876 263880 121458 263936
rect 121514 263880 121519 263936
rect 119876 263878 121519 263880
rect 67633 263875 67699 263878
rect 121453 263875 121519 263878
rect 176377 263938 176443 263941
rect 179086 263938 179092 263940
rect 176377 263936 179092 263938
rect 176377 263880 176382 263936
rect 176438 263880 179092 263936
rect 176377 263878 179092 263880
rect 176377 263875 176443 263878
rect 179086 263876 179092 263878
rect 179156 263938 179162 263940
rect 179156 263878 179890 263938
rect 179156 263876 179162 263878
rect 179830 263870 179890 263878
rect 179830 263810 180044 263870
rect 292806 263666 292866 263908
rect 292806 263606 295442 263666
rect 295382 263532 295442 263606
rect 295374 263468 295380 263532
rect 295444 263530 295450 263532
rect 296345 263530 296411 263533
rect 295444 263528 296411 263530
rect 295444 263472 296350 263528
rect 296406 263472 296411 263528
rect 295444 263470 296411 263472
rect 295444 263468 295450 263470
rect 296345 263467 296411 263470
rect 67725 263258 67791 263261
rect 121453 263258 121519 263261
rect 67725 263256 70196 263258
rect 67725 263200 67730 263256
rect 67786 263200 70196 263256
rect 67725 263198 70196 263200
rect 119876 263256 121519 263258
rect 119876 263200 121458 263256
rect 121514 263200 121519 263256
rect 119876 263198 121519 263200
rect 67725 263195 67791 263198
rect 121453 263195 121519 263198
rect 377305 263258 377371 263261
rect 377990 263258 377996 263260
rect 377305 263256 377996 263258
rect 377305 263200 377310 263256
rect 377366 263200 377996 263256
rect 377305 263198 377996 263200
rect 377305 263195 377371 263198
rect 377990 263196 377996 263198
rect 378060 263258 378066 263260
rect 378060 263198 380052 263258
rect 378060 263196 378066 263198
rect 442717 263122 442783 263125
rect 439852 263120 442783 263122
rect 439852 263064 442722 263120
rect 442778 263064 442783 263120
rect 439852 263062 442783 263064
rect 442717 263059 442783 263062
rect 133781 262850 133847 262853
rect 171910 262850 171916 262852
rect 133781 262848 171916 262850
rect 133781 262792 133786 262848
rect 133842 262792 171916 262848
rect 133781 262790 171916 262792
rect 133781 262787 133847 262790
rect 171910 262788 171916 262790
rect 171980 262788 171986 262852
rect 67633 262578 67699 262581
rect 121545 262578 121611 262581
rect 67633 262576 70196 262578
rect 67633 262520 67638 262576
rect 67694 262520 70196 262576
rect 67633 262518 70196 262520
rect 119876 262576 121611 262578
rect 119876 262520 121550 262576
rect 121606 262520 121611 262576
rect 119876 262518 121611 262520
rect 67633 262515 67699 262518
rect 121545 262515 121611 262518
rect 67725 261898 67791 261901
rect 120165 261898 120231 261901
rect 120901 261898 120967 261901
rect 67725 261896 70196 261898
rect 67725 261840 67730 261896
rect 67786 261840 70196 261896
rect 67725 261838 70196 261840
rect 119876 261896 120967 261898
rect 119876 261840 120170 261896
rect 120226 261840 120906 261896
rect 120962 261840 120967 261896
rect 119876 261838 120967 261840
rect 67725 261835 67791 261838
rect 120165 261835 120231 261838
rect 120901 261835 120967 261838
rect 179462 261770 180044 261830
rect 176653 261762 176719 261765
rect 179462 261762 179522 261770
rect 176653 261760 179522 261762
rect 176653 261704 176658 261760
rect 176714 261704 179522 261760
rect 176653 261702 179522 261704
rect 176653 261699 176719 261702
rect 67633 261218 67699 261221
rect 121453 261218 121519 261221
rect 295333 261218 295399 261221
rect 67633 261216 70196 261218
rect 67633 261160 67638 261216
rect 67694 261160 70196 261216
rect 67633 261158 70196 261160
rect 119876 261216 121519 261218
rect 119876 261160 121458 261216
rect 121514 261160 121519 261216
rect 119876 261158 121519 261160
rect 292836 261216 295399 261218
rect 292836 261160 295338 261216
rect 295394 261160 295399 261216
rect 292836 261158 295399 261160
rect 67633 261155 67699 261158
rect 121453 261155 121519 261158
rect 295333 261155 295399 261158
rect 379329 261218 379395 261221
rect 441705 261218 441771 261221
rect 442809 261218 442875 261221
rect 379329 261216 380052 261218
rect 379329 261160 379334 261216
rect 379390 261160 380052 261216
rect 379329 261158 380052 261160
rect 439852 261216 442875 261218
rect 439852 261160 441710 261216
rect 441766 261160 442814 261216
rect 442870 261160 442875 261216
rect 439852 261158 442875 261160
rect 379329 261155 379395 261158
rect 441705 261155 441771 261158
rect 442809 261155 442875 261158
rect 67633 260538 67699 260541
rect 121453 260538 121519 260541
rect 67633 260536 70196 260538
rect 67633 260480 67638 260536
rect 67694 260480 70196 260536
rect 67633 260478 70196 260480
rect 119876 260536 121519 260538
rect 119876 260480 121458 260536
rect 121514 260480 121519 260536
rect 119876 260478 121519 260480
rect 67633 260475 67699 260478
rect 121453 260475 121519 260478
rect 67725 259858 67791 259861
rect 121453 259858 121519 259861
rect 67725 259856 70196 259858
rect 67725 259800 67730 259856
rect 67786 259800 70196 259856
rect 67725 259798 70196 259800
rect 119876 259856 121519 259858
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 67725 259795 67791 259798
rect 121453 259795 121519 259798
rect 179462 259730 180044 259790
rect 177757 259722 177823 259725
rect 179462 259722 179522 259730
rect 177757 259720 179522 259722
rect 177757 259664 177762 259720
rect 177818 259664 179522 259720
rect 177757 259662 179522 259664
rect 177757 259659 177823 259662
rect 67725 259178 67791 259181
rect 122097 259178 122163 259181
rect 293861 259178 293927 259181
rect 440233 259178 440299 259181
rect 67725 259176 70196 259178
rect 67725 259120 67730 259176
rect 67786 259120 70196 259176
rect 67725 259118 70196 259120
rect 119876 259176 122163 259178
rect 119876 259120 122102 259176
rect 122158 259120 122163 259176
rect 292836 259176 293927 259178
rect 292836 259148 293866 259176
rect 119876 259118 122163 259120
rect 67725 259115 67791 259118
rect 122097 259115 122163 259118
rect 292806 259120 293866 259148
rect 293922 259120 293927 259176
rect 292806 259118 293927 259120
rect 439852 259176 440299 259178
rect 439852 259120 440238 259176
rect 440294 259120 440299 259176
rect 439852 259118 440299 259120
rect 292806 258906 292866 259118
rect 293861 259115 293927 259118
rect 440233 259115 440299 259118
rect 376937 259042 377003 259045
rect 376937 259040 380052 259042
rect 376937 258984 376942 259040
rect 376998 258984 380052 259040
rect 376937 258982 380052 258984
rect 376937 258979 377003 258982
rect 293033 258906 293099 258909
rect 292806 258904 293099 258906
rect 292806 258848 293038 258904
rect 293094 258848 293099 258904
rect 292806 258846 293099 258848
rect 293033 258843 293099 258846
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 69013 258498 69079 258501
rect 121453 258498 121519 258501
rect 69013 258496 70196 258498
rect 69013 258440 69018 258496
rect 69074 258440 70196 258496
rect 69013 258438 70196 258440
rect 119876 258496 121519 258498
rect 119876 258440 121458 258496
rect 121514 258440 121519 258496
rect 119876 258438 121519 258440
rect 69013 258435 69079 258438
rect 121453 258435 121519 258438
rect 67633 257818 67699 257821
rect 121545 257818 121611 257821
rect 67633 257816 70196 257818
rect 67633 257760 67638 257816
rect 67694 257760 70196 257816
rect 67633 257758 70196 257760
rect 119876 257816 121611 257818
rect 119876 257760 121550 257816
rect 121606 257760 121611 257816
rect 119876 257758 121611 257760
rect 67633 257755 67699 257758
rect 121545 257755 121611 257758
rect 121453 257138 121519 257141
rect 295333 257138 295399 257141
rect 440509 257138 440575 257141
rect 119876 257136 121519 257138
rect 59118 256804 59124 256868
rect 59188 256866 59194 256868
rect 70166 256866 70226 257108
rect 119876 257080 121458 257136
rect 121514 257080 121519 257136
rect 119876 257078 121519 257080
rect 292836 257136 295399 257138
rect 292836 257080 295338 257136
rect 295394 257080 295399 257136
rect 292836 257078 295399 257080
rect 439852 257136 440575 257138
rect 439852 257080 440514 257136
rect 440570 257080 440575 257136
rect 439852 257078 440575 257080
rect 121453 257075 121519 257078
rect 295333 257075 295399 257078
rect 440509 257075 440575 257078
rect 179462 257010 180044 257070
rect 176653 257002 176719 257005
rect 179462 257002 179522 257010
rect 176653 257000 179522 257002
rect 176653 256944 176658 257000
rect 176714 256944 179522 257000
rect 176653 256942 179522 256944
rect 176653 256939 176719 256942
rect 378910 256940 378916 257004
rect 378980 257002 378986 257004
rect 378980 256942 380052 257002
rect 378980 256940 378986 256942
rect 59188 256806 70226 256866
rect 59188 256804 59194 256806
rect 67725 256458 67791 256461
rect 121453 256458 121519 256461
rect 67725 256456 70196 256458
rect 67725 256400 67730 256456
rect 67786 256400 70196 256456
rect 67725 256398 70196 256400
rect 119876 256456 121519 256458
rect 119876 256400 121458 256456
rect 121514 256400 121519 256456
rect 119876 256398 121519 256400
rect 67725 256395 67791 256398
rect 121453 256395 121519 256398
rect 67633 255778 67699 255781
rect 121453 255778 121519 255781
rect 67633 255776 70196 255778
rect 67633 255720 67638 255776
rect 67694 255720 70196 255776
rect 67633 255718 70196 255720
rect 119876 255776 121519 255778
rect 119876 255720 121458 255776
rect 121514 255720 121519 255776
rect 119876 255718 121519 255720
rect 67633 255715 67699 255718
rect 121453 255715 121519 255718
rect 67633 255098 67699 255101
rect 122189 255098 122255 255101
rect 67633 255096 70196 255098
rect 67633 255040 67638 255096
rect 67694 255040 70196 255096
rect 67633 255038 70196 255040
rect 119876 255096 122255 255098
rect 119876 255040 122194 255096
rect 122250 255040 122255 255096
rect 119876 255038 122255 255040
rect 67633 255035 67699 255038
rect 122189 255035 122255 255038
rect 176653 255098 176719 255101
rect 295333 255098 295399 255101
rect 443085 255098 443151 255101
rect 176653 255096 179522 255098
rect 176653 255040 176658 255096
rect 176714 255040 179522 255096
rect 176653 255038 179522 255040
rect 292836 255096 295399 255098
rect 292836 255040 295338 255096
rect 295394 255040 295399 255096
rect 292836 255038 295399 255040
rect 439852 255096 443151 255098
rect 439852 255040 443090 255096
rect 443146 255040 443151 255096
rect 439852 255038 443151 255040
rect 176653 255035 176719 255038
rect 179462 255030 179522 255038
rect 295333 255035 295399 255038
rect 443085 255035 443151 255038
rect 179462 254970 180044 255030
rect 67725 254418 67791 254421
rect 121453 254418 121519 254421
rect 67725 254416 70196 254418
rect 67725 254360 67730 254416
rect 67786 254360 70196 254416
rect 67725 254358 70196 254360
rect 119876 254416 121519 254418
rect 119876 254360 121458 254416
rect 121514 254360 121519 254416
rect 119876 254358 121519 254360
rect 67725 254355 67791 254358
rect 121453 254355 121519 254358
rect 377305 254418 377371 254421
rect 378041 254418 378107 254421
rect 377305 254416 380052 254418
rect 377305 254360 377310 254416
rect 377366 254360 378046 254416
rect 378102 254360 380052 254416
rect 377305 254358 380052 254360
rect 377305 254355 377371 254358
rect 378041 254355 378107 254358
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 67633 253738 67699 253741
rect 121453 253738 121519 253741
rect 67633 253736 70196 253738
rect 67633 253680 67638 253736
rect 67694 253680 70196 253736
rect 67633 253678 70196 253680
rect 119876 253736 121519 253738
rect 119876 253680 121458 253736
rect 121514 253680 121519 253736
rect 119876 253678 121519 253680
rect 67633 253675 67699 253678
rect 121453 253675 121519 253678
rect 121545 253058 121611 253061
rect 119876 253056 121611 253058
rect 70166 252650 70226 253028
rect 119876 253000 121550 253056
rect 121606 253000 121611 253056
rect 119876 252998 121611 253000
rect 121545 252995 121611 252998
rect 179462 252930 180044 252990
rect 179321 252922 179387 252925
rect 179462 252922 179522 252930
rect 179321 252920 179522 252922
rect 179321 252864 179326 252920
rect 179382 252864 179522 252920
rect 179321 252862 179522 252864
rect 179321 252859 179387 252862
rect 67590 252590 70226 252650
rect 38561 252514 38627 252517
rect 66846 252514 66852 252516
rect 38561 252512 66852 252514
rect 38561 252456 38566 252512
rect 38622 252456 66852 252512
rect 38561 252454 66852 252456
rect 38561 252451 38627 252454
rect 66846 252452 66852 252454
rect 66916 252514 66922 252516
rect 67590 252514 67650 252590
rect 66916 252454 67650 252514
rect 66916 252452 66922 252454
rect 67541 252378 67607 252381
rect 121545 252378 121611 252381
rect 295333 252378 295399 252381
rect 442901 252378 442967 252381
rect 67541 252376 70196 252378
rect 67541 252320 67546 252376
rect 67602 252320 70196 252376
rect 67541 252318 70196 252320
rect 119876 252376 121611 252378
rect 119876 252320 121550 252376
rect 121606 252320 121611 252376
rect 119876 252318 121611 252320
rect 292836 252376 295399 252378
rect 292836 252320 295338 252376
rect 295394 252320 295399 252376
rect 292836 252318 295399 252320
rect 439852 252376 442967 252378
rect 439852 252320 442906 252376
rect 442962 252320 442967 252376
rect 439852 252318 442967 252320
rect 67541 252315 67607 252318
rect 121545 252315 121611 252318
rect 295333 252315 295399 252318
rect 442901 252315 442967 252318
rect 376937 252242 377003 252245
rect 376937 252240 380052 252242
rect 376937 252184 376942 252240
rect 376998 252184 380052 252240
rect 376937 252182 380052 252184
rect 376937 252179 377003 252182
rect 67633 251698 67699 251701
rect 121453 251698 121519 251701
rect 67633 251696 70196 251698
rect 67633 251640 67638 251696
rect 67694 251640 70196 251696
rect 67633 251638 70196 251640
rect 119876 251696 121519 251698
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 67633 251635 67699 251638
rect 121453 251635 121519 251638
rect 57697 251154 57763 251157
rect 57830 251154 57836 251156
rect 57697 251152 57836 251154
rect 57697 251096 57702 251152
rect 57758 251096 57836 251152
rect 57697 251094 57836 251096
rect 57697 251091 57763 251094
rect 57830 251092 57836 251094
rect 57900 251092 57906 251156
rect 67633 251018 67699 251021
rect 120165 251018 120231 251021
rect 120625 251018 120691 251021
rect 67633 251016 70196 251018
rect 67633 250960 67638 251016
rect 67694 250960 70196 251016
rect 67633 250958 70196 250960
rect 119876 251016 120691 251018
rect 119876 250960 120170 251016
rect 120226 250960 120630 251016
rect 120686 250960 120691 251016
rect 119876 250958 120691 250960
rect 67633 250955 67699 250958
rect 120165 250955 120231 250958
rect 120625 250955 120691 250958
rect 179462 250890 180044 250950
rect 176377 250882 176443 250885
rect 179462 250882 179522 250890
rect 176377 250880 179522 250882
rect 176377 250824 176382 250880
rect 176438 250824 179522 250880
rect 176377 250822 179522 250824
rect 176377 250819 176443 250822
rect 67357 250338 67423 250341
rect 121453 250338 121519 250341
rect 295333 250338 295399 250341
rect 442717 250338 442783 250341
rect 67357 250336 70196 250338
rect 67357 250280 67362 250336
rect 67418 250280 70196 250336
rect 67357 250278 70196 250280
rect 119876 250336 121519 250338
rect 119876 250280 121458 250336
rect 121514 250280 121519 250336
rect 119876 250278 121519 250280
rect 292836 250336 295399 250338
rect 292836 250280 295338 250336
rect 295394 250280 295399 250336
rect 292836 250278 295399 250280
rect 439852 250336 442783 250338
rect 439852 250280 442722 250336
rect 442778 250280 442783 250336
rect 439852 250278 442783 250280
rect 67357 250275 67423 250278
rect 121453 250275 121519 250278
rect 295333 250275 295399 250278
rect 442717 250275 442783 250278
rect 376109 250202 376175 250205
rect 376109 250200 380052 250202
rect 376109 250144 376114 250200
rect 376170 250144 380052 250200
rect 376109 250142 380052 250144
rect 376109 250139 376175 250142
rect 67633 249658 67699 249661
rect 121453 249658 121519 249661
rect 67633 249656 70196 249658
rect 67633 249600 67638 249656
rect 67694 249600 70196 249656
rect 67633 249598 70196 249600
rect 119876 249656 121519 249658
rect 119876 249600 121458 249656
rect 121514 249600 121519 249656
rect 119876 249598 121519 249600
rect 67633 249595 67699 249598
rect 121453 249595 121519 249598
rect 120901 249114 120967 249117
rect 166206 249114 166212 249116
rect 120901 249112 166212 249114
rect 120901 249056 120906 249112
rect 120962 249056 166212 249112
rect 120901 249054 166212 249056
rect 120901 249051 120967 249054
rect 166206 249052 166212 249054
rect 166276 249052 166282 249116
rect 68001 248978 68067 248981
rect 121545 248978 121611 248981
rect 68001 248976 70196 248978
rect 68001 248920 68006 248976
rect 68062 248920 70196 248976
rect 68001 248918 70196 248920
rect 119876 248976 121611 248978
rect 119876 248920 121550 248976
rect 121606 248920 121611 248976
rect 119876 248918 121611 248920
rect 68001 248915 68067 248918
rect 121545 248915 121611 248918
rect 119654 248644 119660 248708
rect 119724 248706 119730 248708
rect 119981 248706 120047 248709
rect 119724 248704 120047 248706
rect 119724 248648 119986 248704
rect 120042 248648 120047 248704
rect 119724 248646 120047 248648
rect 119724 248644 119730 248646
rect 119981 248643 120047 248646
rect 67633 248298 67699 248301
rect 121545 248298 121611 248301
rect 67633 248296 70196 248298
rect 67633 248240 67638 248296
rect 67694 248240 70196 248296
rect 67633 248238 70196 248240
rect 119876 248296 121611 248298
rect 119876 248240 121550 248296
rect 121606 248240 121611 248296
rect 119876 248238 121611 248240
rect 67633 248235 67699 248238
rect 121545 248235 121611 248238
rect 177062 248236 177068 248300
rect 177132 248298 177138 248300
rect 295333 248298 295399 248301
rect 177132 248238 179890 248298
rect 292836 248296 295399 248298
rect 292836 248240 295338 248296
rect 295394 248240 295399 248296
rect 292836 248238 295399 248240
rect 177132 248236 177138 248238
rect 179830 248230 179890 248238
rect 295333 248235 295399 248238
rect 179830 248170 180044 248230
rect 376937 248162 377003 248165
rect 441613 248162 441679 248165
rect 376937 248160 380052 248162
rect 376937 248104 376942 248160
rect 376998 248104 380052 248160
rect 376937 248102 380052 248104
rect 439852 248160 441679 248162
rect 439852 248104 441618 248160
rect 441674 248104 441679 248160
rect 439852 248102 441679 248104
rect 376937 248099 377003 248102
rect 441613 248099 441679 248102
rect 67725 247618 67791 247621
rect 121453 247618 121519 247621
rect 67725 247616 70196 247618
rect 67725 247560 67730 247616
rect 67786 247560 70196 247616
rect 67725 247558 70196 247560
rect 119876 247616 121519 247618
rect 119876 247560 121458 247616
rect 121514 247560 121519 247616
rect 119876 247558 121519 247560
rect 67725 247555 67791 247558
rect 121453 247555 121519 247558
rect 441613 247074 441679 247077
rect 441797 247074 441863 247077
rect 441613 247072 441863 247074
rect 441613 247016 441618 247072
rect 441674 247016 441802 247072
rect 441858 247016 441863 247072
rect 441613 247014 441863 247016
rect 441613 247011 441679 247014
rect 441797 247011 441863 247014
rect 67633 246938 67699 246941
rect 121545 246938 121611 246941
rect 67633 246936 70196 246938
rect 67633 246880 67638 246936
rect 67694 246880 70196 246936
rect 67633 246878 70196 246880
rect 119876 246936 121611 246938
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 67633 246875 67699 246878
rect 121545 246875 121611 246878
rect 120022 246332 120028 246396
rect 120092 246394 120098 246396
rect 166942 246394 166948 246396
rect 120092 246334 166948 246394
rect 120092 246332 120098 246334
rect 166942 246332 166948 246334
rect 167012 246332 167018 246396
rect 68093 246258 68159 246261
rect 121453 246258 121519 246261
rect 293953 246258 294019 246261
rect 294321 246258 294387 246261
rect 68093 246256 70196 246258
rect 68093 246200 68098 246256
rect 68154 246200 70196 246256
rect 68093 246198 70196 246200
rect 119876 246256 121519 246258
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 292836 246256 294387 246258
rect 292836 246200 293958 246256
rect 294014 246200 294326 246256
rect 294382 246200 294387 246256
rect 292836 246198 294387 246200
rect 68093 246195 68159 246198
rect 121453 246195 121519 246198
rect 293953 246195 294019 246198
rect 294321 246195 294387 246198
rect 297398 246196 297404 246260
rect 297468 246258 297474 246260
rect 364701 246258 364767 246261
rect 441613 246258 441679 246261
rect 442901 246258 442967 246261
rect 297468 246256 364767 246258
rect 297468 246200 364706 246256
rect 364762 246200 364767 246256
rect 297468 246198 364767 246200
rect 439852 246256 442967 246258
rect 439852 246200 441618 246256
rect 441674 246200 442906 246256
rect 442962 246200 442967 246256
rect 439852 246198 442967 246200
rect 297468 246196 297474 246198
rect 364701 246195 364767 246198
rect 441613 246195 441679 246198
rect 442901 246195 442967 246198
rect 179462 246130 180044 246190
rect 176653 246122 176719 246125
rect 179462 246122 179522 246130
rect 176653 246120 179522 246122
rect 176653 246064 176658 246120
rect 176714 246064 179522 246120
rect 176653 246062 179522 246064
rect 376937 246122 377003 246125
rect 376937 246120 380052 246122
rect 376937 246064 376942 246120
rect 376998 246064 380052 246120
rect 376937 246062 380052 246064
rect 176653 246059 176719 246062
rect 376937 246059 377003 246062
rect 67633 245578 67699 245581
rect 121545 245578 121611 245581
rect 67633 245576 70196 245578
rect 67633 245520 67638 245576
rect 67694 245520 70196 245576
rect 67633 245518 70196 245520
rect 119876 245576 121611 245578
rect 119876 245520 121550 245576
rect 121606 245520 121611 245576
rect 119876 245518 121611 245520
rect 67633 245515 67699 245518
rect 121545 245515 121611 245518
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 67541 244898 67607 244901
rect 121453 244898 121519 244901
rect 67541 244896 70196 244898
rect 67541 244840 67546 244896
rect 67602 244840 70196 244896
rect 67541 244838 70196 244840
rect 119876 244896 121519 244898
rect 119876 244840 121458 244896
rect 121514 244840 121519 244896
rect 119876 244838 121519 244840
rect 67541 244835 67607 244838
rect 121453 244835 121519 244838
rect 147489 244354 147555 244357
rect 148174 244354 148180 244356
rect 147489 244352 148180 244354
rect 147489 244296 147494 244352
rect 147550 244296 148180 244352
rect 147489 244294 148180 244296
rect 147489 244291 147555 244294
rect 148174 244292 148180 244294
rect 148244 244292 148250 244356
rect 67633 244218 67699 244221
rect 121453 244218 121519 244221
rect 67633 244216 70196 244218
rect 67633 244160 67638 244216
rect 67694 244160 70196 244216
rect 67633 244158 70196 244160
rect 119876 244216 121519 244218
rect 119876 244160 121458 244216
rect 121514 244160 121519 244216
rect 119876 244158 121519 244160
rect 67633 244155 67699 244158
rect 121453 244155 121519 244158
rect 179454 244088 179460 244152
rect 179524 244150 179530 244152
rect 179524 244090 180044 244150
rect 179524 244088 179530 244090
rect 377949 244082 378015 244085
rect 442165 244082 442231 244085
rect 377949 244080 380052 244082
rect 377949 244024 377954 244080
rect 378010 244024 380052 244080
rect 377949 244022 380052 244024
rect 439852 244080 442231 244082
rect 439852 244024 442170 244080
rect 442226 244024 442231 244080
rect 439852 244022 442231 244024
rect 377949 244019 378015 244022
rect 442165 244019 442231 244022
rect 67725 243538 67791 243541
rect 121637 243538 121703 243541
rect 67725 243536 70196 243538
rect 67725 243480 67730 243536
rect 67786 243480 70196 243536
rect 67725 243478 70196 243480
rect 119876 243536 121703 243538
rect 119876 243480 121642 243536
rect 121698 243480 121703 243536
rect 119876 243478 121703 243480
rect 67725 243475 67791 243478
rect 121637 243475 121703 243478
rect 179505 243538 179571 243541
rect 179822 243538 179828 243540
rect 179505 243536 179828 243538
rect 179505 243480 179510 243536
rect 179566 243480 179828 243536
rect 179505 243478 179828 243480
rect 179505 243475 179571 243478
rect 179822 243476 179828 243478
rect 179892 243476 179898 243540
rect 296253 243538 296319 243541
rect 313917 243538 313983 243541
rect 292836 243536 296319 243538
rect 292836 243480 296258 243536
rect 296314 243480 296319 243536
rect 292836 243478 296319 243480
rect 296253 243475 296319 243478
rect 302190 243536 313983 243538
rect 302190 243480 313922 243536
rect 313978 243480 313983 243536
rect 302190 243478 313983 243480
rect 293166 243340 293172 243404
rect 293236 243402 293242 243404
rect 302190 243402 302250 243478
rect 313917 243475 313983 243478
rect 293236 243342 302250 243402
rect 293236 243340 293242 243342
rect 67725 242858 67791 242861
rect 121453 242858 121519 242861
rect 67725 242856 70196 242858
rect 67725 242800 67730 242856
rect 67786 242800 70196 242856
rect 67725 242798 70196 242800
rect 119876 242856 121519 242858
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 67725 242795 67791 242798
rect 121453 242795 121519 242798
rect 292614 242388 292620 242452
rect 292684 242450 292690 242452
rect 294086 242450 294092 242452
rect 292684 242390 294092 242450
rect 292684 242388 292690 242390
rect 294086 242388 294092 242390
rect 294156 242388 294162 242452
rect 379697 242314 379763 242317
rect 373950 242312 379763 242314
rect 373950 242256 379702 242312
rect 379758 242256 379763 242312
rect 373950 242254 379763 242256
rect 67633 242178 67699 242181
rect 121545 242178 121611 242181
rect 67633 242176 70196 242178
rect 67633 242120 67638 242176
rect 67694 242120 70196 242176
rect 67633 242118 70196 242120
rect 119876 242176 121611 242178
rect 119876 242120 121550 242176
rect 121606 242120 121611 242176
rect 119876 242118 121611 242120
rect 67633 242115 67699 242118
rect 121545 242115 121611 242118
rect 349889 242178 349955 242181
rect 373950 242178 374010 242254
rect 379697 242251 379763 242254
rect 442901 242178 442967 242181
rect 349889 242176 374010 242178
rect 349889 242120 349894 242176
rect 349950 242120 374010 242176
rect 349889 242118 374010 242120
rect 439852 242176 442967 242178
rect 439852 242120 442906 242176
rect 442962 242120 442967 242176
rect 439852 242118 442967 242120
rect 349889 242115 349955 242118
rect 442901 242115 442967 242118
rect 179462 242050 180044 242110
rect 176653 242042 176719 242045
rect 179462 242042 179522 242050
rect 176653 242040 179522 242042
rect 176653 241984 176658 242040
rect 176714 241984 179522 242040
rect 176653 241982 179522 241984
rect 376661 242042 376727 242045
rect 376661 242040 380052 242042
rect 376661 241984 376666 242040
rect 376722 241984 380052 242040
rect 376661 241982 380052 241984
rect 176653 241979 176719 241982
rect 376661 241979 376727 241982
rect 293309 241906 293375 241909
rect 302233 241906 302299 241909
rect 293309 241904 302299 241906
rect 293309 241848 293314 241904
rect 293370 241848 302238 241904
rect 302294 241848 302299 241904
rect 293309 241846 302299 241848
rect 293309 241843 293375 241846
rect 302233 241843 302299 241846
rect 373717 241906 373783 241909
rect 373717 241904 374010 241906
rect 373717 241848 373722 241904
rect 373778 241848 374010 241904
rect 373717 241846 374010 241848
rect 373717 241843 373783 241846
rect 373950 241770 374010 241846
rect 382774 241770 382780 241772
rect 373950 241710 382780 241770
rect 382774 241708 382780 241710
rect 382844 241708 382850 241772
rect 67265 241634 67331 241637
rect 70526 241634 70532 241636
rect 67265 241632 70532 241634
rect 67265 241576 67270 241632
rect 67326 241576 70532 241632
rect 67265 241574 70532 241576
rect 67265 241571 67331 241574
rect 70526 241572 70532 241574
rect 70596 241572 70602 241636
rect 67633 241498 67699 241501
rect 120073 241498 120139 241501
rect 296437 241498 296503 241501
rect 67633 241496 70196 241498
rect 67633 241440 67638 241496
rect 67694 241440 70196 241496
rect 67633 241438 70196 241440
rect 119876 241496 120139 241498
rect 119876 241440 120078 241496
rect 120134 241440 120139 241496
rect 119876 241438 120139 241440
rect 292836 241496 296503 241498
rect 292836 241440 296442 241496
rect 296498 241440 296503 241496
rect 292836 241438 296503 241440
rect 67633 241435 67699 241438
rect 120073 241435 120139 241438
rect 296437 241435 296503 241438
rect 119889 241226 119955 241229
rect 120022 241226 120028 241228
rect 119889 241224 120028 241226
rect -960 241090 480 241180
rect 119889 241168 119894 241224
rect 119950 241168 120028 241224
rect 119889 241166 120028 241168
rect 119889 241163 119955 241166
rect 120022 241164 120028 241166
rect 120092 241164 120098 241228
rect 291694 241164 291700 241228
rect 291764 241226 291770 241228
rect 293309 241226 293375 241229
rect 291764 241224 293375 241226
rect 291764 241168 293314 241224
rect 293370 241168 293375 241224
rect 291764 241166 293375 241168
rect 291764 241164 291770 241166
rect 293309 241163 293375 241166
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 67633 240818 67699 240821
rect 121453 240818 121519 240821
rect 67633 240816 70196 240818
rect 67633 240760 67638 240816
rect 67694 240760 70196 240816
rect 67633 240758 70196 240760
rect 119876 240816 121519 240818
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 67633 240755 67699 240758
rect 121453 240755 121519 240758
rect 163589 240818 163655 240821
rect 163589 240816 258090 240818
rect 163589 240760 163594 240816
rect 163650 240760 258090 240816
rect 163589 240758 258090 240760
rect 163589 240755 163655 240758
rect 258030 240682 258090 240758
rect 289486 240756 289492 240820
rect 289556 240818 289562 240820
rect 298185 240818 298251 240821
rect 289556 240816 298251 240818
rect 289556 240760 298190 240816
rect 298246 240760 298251 240816
rect 289556 240758 298251 240760
rect 289556 240756 289562 240758
rect 298185 240755 298251 240758
rect 351177 240818 351243 240821
rect 351177 240816 374010 240818
rect 351177 240760 351182 240816
rect 351238 240760 374010 240816
rect 351177 240758 374010 240760
rect 351177 240755 351243 240758
rect 271137 240682 271203 240685
rect 258030 240680 271203 240682
rect 258030 240624 271142 240680
rect 271198 240624 271203 240680
rect 258030 240622 271203 240624
rect 373950 240682 374010 240758
rect 381629 240682 381695 240685
rect 373950 240680 381695 240682
rect 373950 240624 381634 240680
rect 381690 240624 381695 240680
rect 373950 240622 381695 240624
rect 271137 240619 271203 240622
rect 381629 240619 381695 240622
rect 292614 240484 292620 240548
rect 292684 240546 292690 240548
rect 292941 240546 293007 240549
rect 293166 240546 293172 240548
rect 292684 240544 293172 240546
rect 292684 240488 292946 240544
rect 293002 240488 293172 240544
rect 292684 240486 293172 240488
rect 292684 240484 292690 240486
rect 292941 240483 293007 240486
rect 293166 240484 293172 240486
rect 293236 240484 293242 240548
rect 176377 240274 176443 240277
rect 182817 240274 182883 240277
rect 176377 240272 182883 240274
rect 176377 240216 176382 240272
rect 176438 240216 182822 240272
rect 182878 240216 182883 240272
rect 176377 240214 182883 240216
rect 176377 240211 176443 240214
rect 182817 240211 182883 240214
rect 305085 240274 305151 240277
rect 305637 240274 305703 240277
rect 382273 240274 382339 240277
rect 305085 240272 382339 240274
rect 305085 240216 305090 240272
rect 305146 240216 305642 240272
rect 305698 240216 382278 240272
rect 382334 240216 382339 240272
rect 305085 240214 382339 240216
rect 305085 240211 305151 240214
rect 305637 240211 305703 240214
rect 382273 240211 382339 240214
rect 121637 240138 121703 240141
rect 119876 240136 121703 240138
rect 119876 240080 121642 240136
rect 121698 240080 121703 240136
rect 119876 240078 121703 240080
rect 121637 240075 121703 240078
rect 157374 240076 157380 240140
rect 157444 240138 157450 240140
rect 158253 240138 158319 240141
rect 157444 240136 158319 240138
rect 157444 240080 158258 240136
rect 158314 240080 158319 240136
rect 157444 240078 158319 240080
rect 157444 240076 157450 240078
rect 158253 240075 158319 240078
rect 70526 239804 70532 239868
rect 70596 239866 70602 239868
rect 70669 239866 70735 239869
rect 70596 239864 70735 239866
rect 70596 239808 70674 239864
rect 70730 239808 70735 239864
rect 70596 239806 70735 239808
rect 70596 239804 70602 239806
rect 70669 239803 70735 239806
rect 170673 239594 170739 239597
rect 185577 239594 185643 239597
rect 170673 239592 185643 239594
rect 170673 239536 170678 239592
rect 170734 239536 185582 239592
rect 185638 239536 185643 239592
rect 170673 239534 185643 239536
rect 170673 239531 170739 239534
rect 185577 239531 185643 239534
rect 157241 239458 157307 239461
rect 214557 239458 214623 239461
rect 157241 239456 214623 239458
rect 157241 239400 157246 239456
rect 157302 239400 214562 239456
rect 214618 239400 214623 239456
rect 157241 239398 214623 239400
rect 157241 239395 157307 239398
rect 214557 239395 214623 239398
rect 438853 239458 438919 239461
rect 439270 239458 439330 239972
rect 438853 239456 439330 239458
rect 438853 239400 438858 239456
rect 438914 239400 439330 239456
rect 438853 239398 439330 239400
rect 438853 239395 438919 239398
rect 273989 238778 274055 238781
rect 305085 238778 305151 238781
rect 273989 238776 305151 238778
rect 273989 238720 273994 238776
rect 274050 238720 305090 238776
rect 305146 238720 305151 238776
rect 273989 238718 305151 238720
rect 273989 238715 274055 238718
rect 305085 238715 305151 238718
rect 376150 238716 376156 238780
rect 376220 238778 376226 238780
rect 427905 238778 427971 238781
rect 376220 238776 427971 238778
rect 376220 238720 427910 238776
rect 427966 238720 427971 238776
rect 376220 238718 427971 238720
rect 376220 238716 376226 238718
rect 427905 238715 427971 238718
rect 63350 238580 63356 238644
rect 63420 238642 63426 238644
rect 73889 238642 73955 238645
rect 63420 238640 73955 238642
rect 63420 238584 73894 238640
rect 73950 238584 73955 238640
rect 63420 238582 73955 238584
rect 63420 238580 63426 238582
rect 73889 238579 73955 238582
rect 60641 238506 60707 238509
rect 72601 238506 72667 238509
rect 81617 238506 81683 238509
rect 264973 238506 265039 238509
rect 60641 238504 74550 238506
rect 60641 238448 60646 238504
rect 60702 238448 72606 238504
rect 72662 238448 74550 238504
rect 60641 238446 74550 238448
rect 60641 238443 60707 238446
rect 72601 238443 72667 238446
rect 54334 238308 54340 238372
rect 54404 238370 54410 238372
rect 54753 238370 54819 238373
rect 54404 238368 54819 238370
rect 54404 238312 54758 238368
rect 54814 238312 54819 238368
rect 54404 238310 54819 238312
rect 74490 238370 74550 238446
rect 81617 238504 265039 238506
rect 81617 238448 81622 238504
rect 81678 238448 264978 238504
rect 265034 238448 265039 238504
rect 81617 238446 265039 238448
rect 81617 238443 81683 238446
rect 264973 238443 265039 238446
rect 271781 238506 271847 238509
rect 293217 238506 293283 238509
rect 271781 238504 293283 238506
rect 271781 238448 271786 238504
rect 271842 238448 293222 238504
rect 293278 238448 293283 238504
rect 271781 238446 293283 238448
rect 271781 238443 271847 238446
rect 293217 238443 293283 238446
rect 120758 238370 120764 238372
rect 74490 238310 120764 238370
rect 54404 238308 54410 238310
rect 54753 238307 54819 238310
rect 120758 238308 120764 238310
rect 120828 238308 120834 238372
rect 279417 238370 279483 238373
rect 417417 238370 417483 238373
rect 279417 238368 417483 238370
rect 279417 238312 279422 238368
rect 279478 238312 417422 238368
rect 417478 238312 417483 238368
rect 279417 238310 417483 238312
rect 279417 238307 279483 238310
rect 417417 238307 417483 238310
rect 62849 238234 62915 238237
rect 82261 238234 82327 238237
rect 277945 238234 278011 238237
rect 62849 238232 278011 238234
rect 62849 238176 62854 238232
rect 62910 238176 82266 238232
rect 82322 238176 277950 238232
rect 278006 238176 278011 238232
rect 62849 238174 278011 238176
rect 62849 238171 62915 238174
rect 82261 238171 82327 238174
rect 277945 238171 278011 238174
rect 242249 237962 242315 237965
rect 389817 237962 389883 237965
rect 242249 237960 389883 237962
rect 242249 237904 242254 237960
rect 242310 237904 389822 237960
rect 389878 237904 389883 237960
rect 242249 237902 389883 237904
rect 242249 237899 242315 237902
rect 389817 237899 389883 237902
rect 63166 237220 63172 237284
rect 63236 237282 63242 237284
rect 333329 237282 333395 237285
rect 63236 237280 333395 237282
rect 63236 237224 333334 237280
rect 333390 237224 333395 237280
rect 63236 237222 333395 237224
rect 63236 237220 63242 237222
rect 333329 237219 333395 237222
rect 174997 237146 175063 237149
rect 377949 237146 378015 237149
rect 174997 237144 378015 237146
rect 174997 237088 175002 237144
rect 175058 237088 377954 237144
rect 378010 237088 378015 237144
rect 174997 237086 378015 237088
rect 174997 237083 175063 237086
rect 377949 237083 378015 237086
rect 265525 237010 265591 237013
rect 299606 237010 299612 237012
rect 265525 237008 299612 237010
rect 265525 236952 265530 237008
rect 265586 236952 299612 237008
rect 265525 236950 299612 236952
rect 265525 236947 265591 236950
rect 299606 236948 299612 236950
rect 299676 237010 299682 237012
rect 443177 237010 443243 237013
rect 299676 237008 443243 237010
rect 299676 236952 443182 237008
rect 443238 236952 443243 237008
rect 299676 236950 443243 236952
rect 299676 236948 299682 236950
rect 443177 236947 443243 236950
rect 377949 236194 378015 236197
rect 380566 236194 380572 236196
rect 377949 236192 380572 236194
rect 377949 236136 377954 236192
rect 378010 236136 380572 236192
rect 377949 236134 380572 236136
rect 377949 236131 378015 236134
rect 380566 236132 380572 236134
rect 380636 236132 380642 236196
rect 264053 236058 264119 236061
rect 265525 236058 265591 236061
rect 264053 236056 265591 236058
rect 264053 236000 264058 236056
rect 264114 236000 265530 236056
rect 265586 236000 265591 236056
rect 264053 235998 265591 236000
rect 264053 235995 264119 235998
rect 265525 235995 265591 235998
rect 332593 236058 332659 236061
rect 333329 236058 333395 236061
rect 332593 236056 333395 236058
rect 332593 236000 332598 236056
rect 332654 236000 333334 236056
rect 333390 236000 333395 236056
rect 332593 235998 333395 236000
rect 332593 235995 332659 235998
rect 333329 235995 333395 235998
rect 377990 235996 377996 236060
rect 378060 236058 378066 236060
rect 383009 236058 383075 236061
rect 378060 236056 383075 236058
rect 378060 236000 383014 236056
rect 383070 236000 383075 236056
rect 378060 235998 383075 236000
rect 378060 235996 378066 235998
rect 383009 235995 383075 235998
rect 93209 235922 93275 235925
rect 93761 235922 93827 235925
rect 120574 235922 120580 235924
rect 93209 235920 120580 235922
rect 93209 235864 93214 235920
rect 93270 235864 93766 235920
rect 93822 235864 120580 235920
rect 93209 235862 120580 235864
rect 93209 235859 93275 235862
rect 93761 235859 93827 235862
rect 120574 235860 120580 235862
rect 120644 235860 120650 235924
rect 121637 235922 121703 235925
rect 318149 235922 318215 235925
rect 121637 235920 318215 235922
rect 121637 235864 121642 235920
rect 121698 235864 318154 235920
rect 318210 235864 318215 235920
rect 121637 235862 318215 235864
rect 121637 235859 121703 235862
rect 318149 235859 318215 235862
rect 171910 235180 171916 235244
rect 171980 235242 171986 235244
rect 239397 235242 239463 235245
rect 171980 235240 239463 235242
rect 171980 235184 239402 235240
rect 239458 235184 239463 235240
rect 171980 235182 239463 235184
rect 171980 235180 171986 235182
rect 239397 235179 239463 235182
rect 65793 233882 65859 233885
rect 259494 233882 259500 233884
rect 65793 233880 259500 233882
rect 65793 233824 65798 233880
rect 65854 233824 259500 233880
rect 65793 233822 259500 233824
rect 65793 233819 65859 233822
rect 259494 233820 259500 233822
rect 259564 233820 259570 233884
rect 380934 233276 380940 233340
rect 381004 233338 381010 233340
rect 485773 233338 485839 233341
rect 381004 233336 485839 233338
rect 381004 233280 485778 233336
rect 485834 233280 485839 233336
rect 381004 233278 485839 233280
rect 381004 233276 381010 233278
rect 485773 233275 485839 233278
rect 259361 233204 259427 233205
rect 259310 233202 259316 233204
rect 259270 233142 259316 233202
rect 259380 233202 259427 233204
rect 288525 233202 288591 233205
rect 378726 233202 378732 233204
rect 259380 233200 267750 233202
rect 259422 233144 267750 233200
rect 259310 233140 259316 233142
rect 259380 233142 267750 233144
rect 259380 233140 259427 233142
rect 259361 233139 259427 233140
rect 267690 233066 267750 233142
rect 288525 233200 378732 233202
rect 288525 233144 288530 233200
rect 288586 233144 378732 233200
rect 288525 233142 378732 233144
rect 288525 233139 288591 233142
rect 378726 233140 378732 233142
rect 378796 233140 378802 233204
rect 311014 233066 311020 233068
rect 267690 233006 311020 233066
rect 311014 233004 311020 233006
rect 311084 233004 311090 233068
rect 262121 232522 262187 232525
rect 278681 232522 278747 232525
rect 318006 232522 318012 232524
rect 262121 232520 318012 232522
rect 262121 232464 262126 232520
rect 262182 232464 278686 232520
rect 278742 232464 318012 232520
rect 262121 232462 318012 232464
rect 262121 232459 262187 232462
rect 278681 232459 278747 232462
rect 318006 232460 318012 232462
rect 318076 232460 318082 232524
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect 271086 232052 271092 232116
rect 271156 232114 271162 232116
rect 271229 232114 271295 232117
rect 271156 232112 271295 232114
rect 271156 232056 271234 232112
rect 271290 232056 271295 232112
rect 271156 232054 271295 232056
rect 271156 232052 271162 232054
rect 271229 232051 271295 232054
rect 362953 231842 363019 231845
rect 364149 231842 364215 231845
rect 380934 231842 380940 231844
rect 362953 231840 380940 231842
rect 362953 231784 362958 231840
rect 363014 231784 364154 231840
rect 364210 231784 380940 231840
rect 362953 231782 380940 231784
rect 362953 231779 363019 231782
rect 364149 231779 364215 231782
rect 380934 231780 380940 231782
rect 381004 231780 381010 231844
rect 288198 231236 288204 231300
rect 288268 231298 288274 231300
rect 296713 231298 296779 231301
rect 288268 231296 296779 231298
rect 288268 231240 296718 231296
rect 296774 231240 296779 231296
rect 288268 231238 296779 231240
rect 288268 231236 288274 231238
rect 296713 231235 296779 231238
rect 270401 231162 270467 231165
rect 291878 231162 291884 231164
rect 270401 231160 291884 231162
rect 270401 231104 270406 231160
rect 270462 231104 291884 231160
rect 270401 231102 291884 231104
rect 270401 231099 270467 231102
rect 291878 231100 291884 231102
rect 291948 231100 291954 231164
rect 122189 230482 122255 230485
rect 322749 230482 322815 230485
rect 322974 230482 322980 230484
rect 122189 230480 322980 230482
rect 122189 230424 122194 230480
rect 122250 230424 322754 230480
rect 322810 230424 322980 230480
rect 122189 230422 322980 230424
rect 122189 230419 122255 230422
rect 322749 230419 322815 230422
rect 322974 230420 322980 230422
rect 323044 230420 323050 230484
rect 165521 228306 165587 228309
rect 378041 228306 378107 228309
rect 165521 228304 378107 228306
rect 165521 228248 165526 228304
rect 165582 228248 378046 228304
rect 378102 228248 378107 228304
rect 165521 228246 378107 228248
rect 165521 228243 165587 228246
rect 378041 228243 378107 228246
rect -960 227884 480 228124
rect 378041 227762 378107 227765
rect 378910 227762 378916 227764
rect 378041 227760 378916 227762
rect 378041 227704 378046 227760
rect 378102 227704 378916 227760
rect 378041 227702 378916 227704
rect 378041 227699 378107 227702
rect 378910 227700 378916 227702
rect 378980 227700 378986 227764
rect 161974 227020 161980 227084
rect 162044 227082 162050 227084
rect 211797 227082 211863 227085
rect 162044 227080 211863 227082
rect 162044 227024 211802 227080
rect 211858 227024 211863 227080
rect 162044 227022 211863 227024
rect 162044 227020 162050 227022
rect 211797 227019 211863 227022
rect 59118 226884 59124 226948
rect 59188 226946 59194 226948
rect 318701 226946 318767 226949
rect 323117 226946 323183 226949
rect 59188 226944 323183 226946
rect 59188 226888 318706 226944
rect 318762 226888 323122 226944
rect 323178 226888 323183 226944
rect 59188 226886 323183 226888
rect 59188 226884 59194 226886
rect 318701 226883 318767 226886
rect 323117 226883 323183 226886
rect 378726 226884 378732 226948
rect 378796 226946 378802 226948
rect 414289 226946 414355 226949
rect 378796 226944 414355 226946
rect 378796 226888 414294 226944
rect 414350 226888 414355 226944
rect 378796 226886 414355 226888
rect 378796 226884 378802 226886
rect 414289 226883 414355 226886
rect 298001 225586 298067 225589
rect 313774 225586 313780 225588
rect 298001 225584 313780 225586
rect 298001 225528 298006 225584
rect 298062 225528 313780 225584
rect 298001 225526 313780 225528
rect 298001 225523 298067 225526
rect 313774 225524 313780 225526
rect 313844 225524 313850 225588
rect 253933 224906 253999 224909
rect 454125 224908 454191 224909
rect 454125 224906 454172 224908
rect 253933 224904 454172 224906
rect 253933 224848 253938 224904
rect 253994 224848 454130 224904
rect 253933 224846 454172 224848
rect 253933 224843 253999 224846
rect 454125 224844 454172 224846
rect 454236 224844 454242 224908
rect 454125 224843 454191 224844
rect 342294 224436 342300 224500
rect 342364 224498 342370 224500
rect 342989 224498 343055 224501
rect 342364 224496 343055 224498
rect 342364 224440 342994 224496
rect 343050 224440 343055 224496
rect 342364 224438 343055 224440
rect 342364 224436 342370 224438
rect 342989 224435 343055 224438
rect 187693 222186 187759 222189
rect 188981 222186 189047 222189
rect 187693 222184 189047 222186
rect 187693 222128 187698 222184
rect 187754 222128 188986 222184
rect 189042 222128 189047 222184
rect 187693 222126 189047 222128
rect 187693 222123 187759 222126
rect 188981 222123 189047 222126
rect 167678 221444 167684 221508
rect 167748 221506 167754 221508
rect 185577 221506 185643 221509
rect 167748 221504 185643 221506
rect 167748 221448 185582 221504
rect 185638 221448 185643 221504
rect 167748 221446 185643 221448
rect 167748 221444 167754 221446
rect 185577 221443 185643 221446
rect 188981 220962 189047 220965
rect 448462 220962 448468 220964
rect 188981 220960 448468 220962
rect 188981 220904 188986 220960
rect 189042 220904 448468 220960
rect 188981 220902 448468 220904
rect 188981 220899 189047 220902
rect 448462 220900 448468 220902
rect 448532 220900 448538 220964
rect 208393 220826 208459 220829
rect 209681 220826 209747 220829
rect 301446 220826 301452 220828
rect 208393 220824 301452 220826
rect 208393 220768 208398 220824
rect 208454 220768 209686 220824
rect 209742 220768 301452 220824
rect 208393 220766 301452 220768
rect 208393 220763 208459 220766
rect 209681 220763 209747 220766
rect 301446 220764 301452 220766
rect 301516 220764 301522 220828
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 286961 218650 287027 218653
rect 309174 218650 309180 218652
rect 286961 218648 309180 218650
rect 286961 218592 286966 218648
rect 287022 218592 309180 218648
rect 286961 218590 309180 218592
rect 286961 218587 287027 218590
rect 309174 218588 309180 218590
rect 309244 218588 309250 218652
rect 152457 217970 152523 217973
rect 324814 217970 324820 217972
rect 152457 217968 324820 217970
rect 152457 217912 152462 217968
rect 152518 217912 324820 217968
rect 152457 217910 324820 217912
rect 152457 217907 152523 217910
rect 324814 217908 324820 217910
rect 324884 217908 324890 217972
rect 160686 217364 160692 217428
rect 160756 217426 160762 217428
rect 313181 217426 313247 217429
rect 160756 217424 313247 217426
rect 160756 217368 313186 217424
rect 313242 217368 313247 217424
rect 160756 217366 313247 217368
rect 160756 217364 160762 217366
rect 313181 217363 313247 217366
rect 53465 217290 53531 217293
rect 256734 217290 256740 217292
rect 53465 217288 256740 217290
rect 53465 217232 53470 217288
rect 53526 217232 256740 217288
rect 53465 217230 256740 217232
rect 53465 217227 53531 217230
rect 256734 217228 256740 217230
rect 256804 217228 256810 217292
rect 313181 216746 313247 216749
rect 314653 216746 314719 216749
rect 313181 216744 314719 216746
rect 313181 216688 313186 216744
rect 313242 216688 314658 216744
rect 314714 216688 314719 216744
rect 313181 216686 314719 216688
rect 313181 216683 313247 216686
rect 314653 216683 314719 216686
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 164969 214570 165035 214573
rect 255262 214570 255268 214572
rect 164969 214568 255268 214570
rect 164969 214512 164974 214568
rect 165030 214512 255268 214568
rect 164969 214510 255268 214512
rect 164969 214507 165035 214510
rect 255262 214508 255268 214510
rect 255332 214508 255338 214572
rect 180793 214434 180859 214437
rect 182081 214434 182147 214437
rect 180793 214432 182147 214434
rect 180793 214376 180798 214432
rect 180854 214376 182086 214432
rect 182142 214376 182147 214432
rect 180793 214374 182147 214376
rect 180793 214371 180859 214374
rect 182081 214371 182147 214374
rect 182081 214026 182147 214029
rect 451038 214026 451044 214028
rect 182081 214024 451044 214026
rect 182081 213968 182086 214024
rect 182142 213968 451044 214024
rect 182081 213966 451044 213968
rect 182081 213963 182147 213966
rect 451038 213964 451044 213966
rect 451108 213964 451114 214028
rect 68921 210354 68987 210357
rect 261334 210354 261340 210356
rect 68921 210352 261340 210354
rect 68921 210296 68926 210352
rect 68982 210296 261340 210352
rect 68921 210294 261340 210296
rect 68921 210291 68987 210294
rect 261334 210292 261340 210294
rect 261404 210292 261410 210356
rect 322841 209810 322907 209813
rect 329782 209810 329788 209812
rect 322841 209808 329788 209810
rect 322841 209752 322846 209808
rect 322902 209752 329788 209808
rect 322841 209750 329788 209752
rect 322841 209747 322907 209750
rect 329782 209748 329788 209750
rect 329852 209748 329858 209812
rect 322933 207090 322999 207093
rect 323158 207090 323164 207092
rect 322933 207088 323164 207090
rect 322933 207032 322938 207088
rect 322994 207032 323164 207088
rect 322933 207030 323164 207032
rect 322933 207027 322999 207030
rect 323158 207028 323164 207030
rect 323228 207028 323234 207092
rect 142654 206892 142660 206956
rect 142724 206954 142730 206956
rect 334617 206954 334683 206957
rect 142724 206952 334683 206954
rect 142724 206896 334622 206952
rect 334678 206896 334683 206952
rect 142724 206894 334683 206896
rect 142724 206892 142730 206894
rect 334617 206891 334683 206894
rect 334014 205668 334020 205732
rect 334084 205730 334090 205732
rect 334617 205730 334683 205733
rect 334084 205728 334683 205730
rect 334084 205672 334622 205728
rect 334678 205672 334683 205728
rect 334084 205670 334683 205672
rect 334084 205668 334090 205670
rect 334617 205667 334683 205670
rect 579981 205730 580047 205733
rect 583520 205730 584960 205820
rect 579981 205728 584960 205730
rect 579981 205672 579986 205728
rect 580042 205672 584960 205728
rect 579981 205670 584960 205672
rect 579981 205667 580047 205670
rect 125777 205596 125843 205597
rect 125726 205594 125732 205596
rect 125686 205534 125732 205594
rect 125796 205592 125843 205596
rect 125838 205536 125843 205592
rect 583520 205580 584960 205670
rect 125726 205532 125732 205534
rect 125796 205532 125843 205536
rect 125777 205531 125843 205532
rect 295926 202132 295932 202196
rect 295996 202194 296002 202196
rect 349245 202194 349311 202197
rect 295996 202192 349311 202194
rect 295996 202136 349250 202192
rect 349306 202136 349311 202192
rect 295996 202134 349311 202136
rect 295996 202132 296002 202134
rect 349245 202131 349311 202134
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 349245 201514 349311 201517
rect 446581 201514 446647 201517
rect 349245 201512 446647 201514
rect 349245 201456 349250 201512
rect 349306 201456 446586 201512
rect 446642 201456 446647 201512
rect 349245 201454 446647 201456
rect 349245 201451 349311 201454
rect 446581 201451 446647 201454
rect 158161 200018 158227 200021
rect 331806 200018 331812 200020
rect 158161 200016 331812 200018
rect 158161 199960 158166 200016
rect 158222 199960 331812 200016
rect 158161 199958 331812 199960
rect 158161 199955 158227 199958
rect 331806 199956 331812 199958
rect 331876 199956 331882 200020
rect 157190 199276 157196 199340
rect 157260 199338 157266 199340
rect 210417 199338 210483 199341
rect 157260 199336 210483 199338
rect 157260 199280 210422 199336
rect 210478 199280 210483 199336
rect 157260 199278 210483 199280
rect 157260 199276 157266 199278
rect 210417 199275 210483 199278
rect 331397 198794 331463 198797
rect 331806 198794 331812 198796
rect 331397 198792 331812 198794
rect 331397 198736 331402 198792
rect 331458 198736 331812 198792
rect 331397 198734 331812 198736
rect 331397 198731 331463 198734
rect 331806 198732 331812 198734
rect 331876 198732 331882 198796
rect 292665 198116 292731 198117
rect 292614 198052 292620 198116
rect 292684 198114 292731 198116
rect 292684 198112 292776 198114
rect 292726 198056 292776 198112
rect 292684 198054 292776 198056
rect 292684 198052 292731 198054
rect 292665 198051 292731 198052
rect 43897 197298 43963 197301
rect 333237 197298 333303 197301
rect 43897 197296 333303 197298
rect 43897 197240 43902 197296
rect 43958 197240 333242 197296
rect 333298 197240 333303 197296
rect 43897 197238 333303 197240
rect 43897 197235 43963 197238
rect 333237 197235 333303 197238
rect 324814 196556 324820 196620
rect 324884 196618 324890 196620
rect 347773 196618 347839 196621
rect 324884 196616 347839 196618
rect 324884 196560 347778 196616
rect 347834 196560 347839 196616
rect 324884 196558 347839 196560
rect 324884 196556 324890 196558
rect 347773 196555 347839 196558
rect 332542 196012 332548 196076
rect 332612 196074 332618 196076
rect 333237 196074 333303 196077
rect 332612 196072 333303 196074
rect 332612 196016 333242 196072
rect 333298 196016 333303 196072
rect 332612 196014 333303 196016
rect 332612 196012 332618 196014
rect 333237 196011 333303 196014
rect 335445 196074 335511 196077
rect 335670 196074 335676 196076
rect 335445 196072 335676 196074
rect 335445 196016 335450 196072
rect 335506 196016 335676 196072
rect 335445 196014 335676 196016
rect 335445 196011 335511 196014
rect 335670 196012 335676 196014
rect 335740 196012 335746 196076
rect 56409 195258 56475 195261
rect 259678 195258 259684 195260
rect 56409 195256 259684 195258
rect 56409 195200 56414 195256
rect 56470 195200 259684 195256
rect 56409 195198 259684 195200
rect 56409 195195 56475 195198
rect 259678 195196 259684 195198
rect 259748 195196 259754 195260
rect 115841 192674 115907 192677
rect 322054 192674 322060 192676
rect 115841 192672 322060 192674
rect 115841 192616 115846 192672
rect 115902 192616 322060 192672
rect 115841 192614 322060 192616
rect 115841 192611 115907 192614
rect 322054 192612 322060 192614
rect 322124 192612 322130 192676
rect 56501 192538 56567 192541
rect 320214 192538 320220 192540
rect 56501 192536 320220 192538
rect 56501 192480 56506 192536
rect 56562 192480 320220 192536
rect 56501 192478 320220 192480
rect 56501 192475 56567 192478
rect 320214 192476 320220 192478
rect 320284 192476 320290 192540
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 113081 191178 113147 191181
rect 346342 191178 346348 191180
rect 113081 191176 346348 191178
rect 113081 191120 113086 191176
rect 113142 191120 346348 191176
rect 113081 191118 346348 191120
rect 113081 191115 113147 191118
rect 346342 191116 346348 191118
rect 346412 191116 346418 191180
rect 66846 190980 66852 191044
rect 66916 191042 66922 191044
rect 324405 191042 324471 191045
rect 66916 191040 324471 191042
rect 66916 190984 324410 191040
rect 324466 190984 324471 191040
rect 66916 190982 324471 190984
rect 66916 190980 66922 190982
rect 324405 190979 324471 190982
rect 138749 189682 138815 189685
rect 263542 189682 263548 189684
rect 138749 189680 263548 189682
rect 138749 189624 138754 189680
rect 138810 189624 263548 189680
rect 138749 189622 263548 189624
rect 138749 189619 138815 189622
rect 263542 189620 263548 189622
rect 263612 189620 263618 189684
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 166206 187172 166212 187236
rect 166276 187234 166282 187236
rect 313917 187234 313983 187237
rect 166276 187232 313983 187234
rect 166276 187176 313922 187232
rect 313978 187176 313983 187232
rect 166276 187174 313983 187176
rect 166276 187172 166282 187174
rect 313917 187171 313983 187174
rect 146886 187036 146892 187100
rect 146956 187098 146962 187100
rect 342437 187098 342503 187101
rect 146956 187096 342503 187098
rect 146956 187040 342442 187096
rect 342498 187040 342503 187096
rect 146956 187038 342503 187040
rect 146956 187036 146962 187038
rect 342437 187035 342503 187038
rect 50981 186962 51047 186965
rect 262254 186962 262260 186964
rect 50981 186960 262260 186962
rect 50981 186904 50986 186960
rect 51042 186904 262260 186960
rect 50981 186902 262260 186904
rect 50981 186899 51047 186902
rect 262254 186900 262260 186902
rect 262324 186900 262330 186964
rect 159357 185738 159423 185741
rect 252502 185738 252508 185740
rect 159357 185736 252508 185738
rect 159357 185680 159362 185736
rect 159418 185680 252508 185736
rect 159357 185678 252508 185680
rect 159357 185675 159423 185678
rect 252502 185676 252508 185678
rect 252572 185676 252578 185740
rect 124806 185540 124812 185604
rect 124876 185602 124882 185604
rect 335629 185602 335695 185605
rect 124876 185600 335695 185602
rect 124876 185544 335634 185600
rect 335690 185544 335695 185600
rect 124876 185542 335695 185544
rect 124876 185540 124882 185542
rect 335629 185539 335695 185542
rect 155217 184378 155283 184381
rect 255446 184378 255452 184380
rect 155217 184376 255452 184378
rect 155217 184320 155222 184376
rect 155278 184320 255452 184376
rect 155217 184318 255452 184320
rect 155217 184315 155283 184318
rect 255446 184316 255452 184318
rect 255516 184316 255522 184380
rect 130377 184242 130443 184245
rect 169702 184242 169708 184244
rect 130377 184240 169708 184242
rect 130377 184184 130382 184240
rect 130438 184184 169708 184240
rect 130377 184182 169708 184184
rect 130377 184179 130443 184182
rect 169702 184180 169708 184182
rect 169772 184180 169778 184244
rect 211797 184242 211863 184245
rect 328678 184242 328684 184244
rect 211797 184240 328684 184242
rect 211797 184184 211802 184240
rect 211858 184184 328684 184240
rect 211797 184182 328684 184184
rect 211797 184179 211863 184182
rect 328678 184180 328684 184182
rect 328748 184180 328754 184244
rect 171501 182882 171567 182885
rect 327022 182882 327028 182884
rect 171501 182880 327028 182882
rect 171501 182824 171506 182880
rect 171562 182824 327028 182880
rect 171501 182822 327028 182824
rect 171501 182819 171567 182822
rect 327022 182820 327028 182822
rect 327092 182820 327098 182884
rect 114369 182202 114435 182205
rect 166206 182202 166212 182204
rect 114369 182200 166212 182202
rect 114369 182144 114374 182200
rect 114430 182144 166212 182200
rect 114369 182142 166212 182144
rect 114369 182139 114435 182142
rect 166206 182140 166212 182142
rect 166276 182140 166282 182204
rect 149789 181658 149855 181661
rect 263726 181658 263732 181660
rect 149789 181656 263732 181658
rect 149789 181600 149794 181656
rect 149850 181600 263732 181656
rect 149789 181598 263732 181600
rect 149789 181595 149855 181598
rect 263726 181596 263732 181598
rect 263796 181596 263802 181660
rect 149646 181460 149652 181524
rect 149716 181522 149722 181524
rect 332777 181522 332843 181525
rect 149716 181520 332843 181522
rect 149716 181464 332782 181520
rect 332838 181464 332843 181520
rect 149716 181462 332843 181464
rect 149716 181460 149722 181462
rect 332777 181459 332843 181462
rect 66161 181386 66227 181389
rect 251214 181386 251220 181388
rect 66161 181384 251220 181386
rect 66161 181328 66166 181384
rect 66222 181328 251220 181384
rect 66161 181326 251220 181328
rect 66161 181323 66227 181326
rect 251214 181324 251220 181326
rect 251284 181324 251290 181388
rect 273897 181386 273963 181389
rect 331254 181386 331260 181388
rect 273897 181384 331260 181386
rect 273897 181328 273902 181384
rect 273958 181328 331260 181384
rect 273897 181326 331260 181328
rect 273897 181323 273963 181326
rect 331254 181324 331260 181326
rect 331324 181324 331330 181388
rect 134517 180162 134583 180165
rect 256918 180162 256924 180164
rect 134517 180160 256924 180162
rect 134517 180104 134522 180160
rect 134578 180104 256924 180160
rect 134517 180102 256924 180104
rect 134517 180099 134583 180102
rect 256918 180100 256924 180102
rect 256988 180100 256994 180164
rect 170489 180026 170555 180029
rect 347865 180026 347931 180029
rect 170489 180024 347931 180026
rect 170489 179968 170494 180024
rect 170550 179968 347870 180024
rect 347926 179968 347931 180024
rect 170489 179966 347931 179968
rect 170489 179963 170555 179966
rect 347865 179963 347931 179966
rect 398741 180026 398807 180029
rect 534206 180026 534212 180028
rect 398741 180024 534212 180026
rect 398741 179968 398746 180024
rect 398802 179968 534212 180024
rect 398741 179966 534212 179968
rect 398741 179963 398807 179966
rect 534206 179964 534212 179966
rect 534276 179964 534282 180028
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 232497 178938 232563 178941
rect 249006 178938 249012 178940
rect 232497 178936 249012 178938
rect 232497 178880 232502 178936
rect 232558 178880 249012 178936
rect 232497 178878 249012 178880
rect 232497 178875 232563 178878
rect 249006 178876 249012 178878
rect 249076 178876 249082 178940
rect 314469 178938 314535 178941
rect 328494 178938 328500 178940
rect 314469 178936 328500 178938
rect 314469 178880 314474 178936
rect 314530 178880 328500 178936
rect 314469 178878 328500 178880
rect 314469 178875 314535 178878
rect 328494 178876 328500 178878
rect 328564 178876 328570 178940
rect 246297 178802 246363 178805
rect 326654 178802 326660 178804
rect 246297 178800 326660 178802
rect 246297 178744 246302 178800
rect 246358 178744 326660 178800
rect 246297 178742 326660 178744
rect 246297 178739 246363 178742
rect 326654 178740 326660 178742
rect 326724 178740 326730 178804
rect 336825 178802 336891 178805
rect 337878 178802 337884 178804
rect 336825 178800 337884 178802
rect 336825 178744 336830 178800
rect 336886 178744 337884 178800
rect 336825 178742 337884 178744
rect 336825 178739 336891 178742
rect 337878 178740 337884 178742
rect 337948 178740 337954 178804
rect 167494 178604 167500 178668
rect 167564 178666 167570 178668
rect 343725 178666 343791 178669
rect 167564 178664 343791 178666
rect 167564 178608 343730 178664
rect 343786 178608 343791 178664
rect 167564 178606 343791 178608
rect 167564 178604 167570 178606
rect 343725 178603 343791 178606
rect 166390 178122 166396 178124
rect 110646 178062 166396 178122
rect 110646 177988 110706 178062
rect 166390 178060 166396 178062
rect 166460 178060 166466 178124
rect 110638 177924 110644 177988
rect 110708 177924 110714 177988
rect 247861 177850 247927 177853
rect 249742 177850 249748 177852
rect 247861 177848 249748 177850
rect 247861 177792 247866 177848
rect 247922 177792 249748 177848
rect 247861 177790 249748 177792
rect 247861 177787 247927 177790
rect 249742 177788 249748 177790
rect 249812 177788 249818 177852
rect 99414 177516 99420 177580
rect 99484 177578 99490 177580
rect 100661 177578 100727 177581
rect 99484 177576 100727 177578
rect 99484 177520 100666 177576
rect 100722 177520 100727 177576
rect 99484 177518 100727 177520
rect 99484 177516 99490 177518
rect 100661 177515 100727 177518
rect 106038 177516 106044 177580
rect 106108 177578 106114 177580
rect 106181 177578 106247 177581
rect 106108 177576 106247 177578
rect 106108 177520 106186 177576
rect 106242 177520 106247 177576
rect 106108 177518 106247 177520
rect 106108 177516 106114 177518
rect 106181 177515 106247 177518
rect 106958 177516 106964 177580
rect 107028 177578 107034 177580
rect 107561 177578 107627 177581
rect 107028 177576 107627 177578
rect 107028 177520 107566 177576
rect 107622 177520 107627 177576
rect 107028 177518 107627 177520
rect 107028 177516 107034 177518
rect 107561 177515 107627 177518
rect 112110 177516 112116 177580
rect 112180 177578 112186 177580
rect 112621 177578 112687 177581
rect 112180 177576 112687 177578
rect 112180 177520 112626 177576
rect 112682 177520 112687 177576
rect 112180 177518 112687 177520
rect 112180 177516 112186 177518
rect 112621 177515 112687 177518
rect 114134 177516 114140 177580
rect 114204 177578 114210 177580
rect 114369 177578 114435 177581
rect 114204 177576 114435 177578
rect 114204 177520 114374 177576
rect 114430 177520 114435 177576
rect 114204 177518 114435 177520
rect 114204 177516 114210 177518
rect 114369 177515 114435 177518
rect 120758 177516 120764 177580
rect 120828 177578 120834 177580
rect 121177 177578 121243 177581
rect 120828 177576 121243 177578
rect 120828 177520 121182 177576
rect 121238 177520 121243 177576
rect 120828 177518 121243 177520
rect 120828 177516 120834 177518
rect 121177 177515 121243 177518
rect 122966 177516 122972 177580
rect 123036 177578 123042 177580
rect 124121 177578 124187 177581
rect 123036 177576 124187 177578
rect 123036 177520 124126 177576
rect 124182 177520 124187 177576
rect 123036 177518 124187 177520
rect 123036 177516 123042 177518
rect 124121 177515 124187 177518
rect 127014 177516 127020 177580
rect 127084 177578 127090 177580
rect 127801 177578 127867 177581
rect 127084 177576 127867 177578
rect 127084 177520 127806 177576
rect 127862 177520 127867 177576
rect 127084 177518 127867 177520
rect 127084 177516 127090 177518
rect 127801 177515 127867 177518
rect 245653 177578 245719 177581
rect 249190 177578 249196 177580
rect 245653 177576 249196 177578
rect 245653 177520 245658 177576
rect 245714 177520 249196 177576
rect 245653 177518 249196 177520
rect 245653 177515 245719 177518
rect 249190 177516 249196 177518
rect 249260 177516 249266 177580
rect 315941 177442 316007 177445
rect 331438 177442 331444 177444
rect 315941 177440 331444 177442
rect 315941 177384 315946 177440
rect 316002 177384 331444 177440
rect 315941 177382 331444 177384
rect 315941 177379 316007 177382
rect 331438 177380 331444 177382
rect 331508 177380 331514 177444
rect 113214 177244 113220 177308
rect 113284 177306 113290 177308
rect 114461 177306 114527 177309
rect 113284 177304 114527 177306
rect 113284 177248 114466 177304
rect 114522 177248 114527 177304
rect 113284 177246 114527 177248
rect 113284 177244 113290 177246
rect 114461 177243 114527 177246
rect 156597 177306 156663 177309
rect 325969 177306 326035 177309
rect 156597 177304 326035 177306
rect 156597 177248 156602 177304
rect 156658 177248 325974 177304
rect 326030 177248 326035 177304
rect 156597 177246 326035 177248
rect 156597 177243 156663 177246
rect 325969 177243 326035 177246
rect 115841 177172 115907 177173
rect 116945 177172 117011 177173
rect 115790 177170 115796 177172
rect 115750 177110 115796 177170
rect 115860 177168 115907 177172
rect 116894 177170 116900 177172
rect 115902 177112 115907 177168
rect 115790 177108 115796 177110
rect 115860 177108 115907 177112
rect 116854 177110 116900 177170
rect 116964 177168 117011 177172
rect 117006 177112 117011 177168
rect 116894 177108 116900 177110
rect 116964 177108 117011 177112
rect 124438 177108 124444 177172
rect 124508 177170 124514 177172
rect 124949 177170 125015 177173
rect 148225 177172 148291 177173
rect 148174 177170 148180 177172
rect 124508 177168 125015 177170
rect 124508 177112 124954 177168
rect 125010 177112 125015 177168
rect 124508 177110 125015 177112
rect 148134 177110 148180 177170
rect 148244 177168 148291 177172
rect 148286 177112 148291 177168
rect 124508 177108 124514 177110
rect 115841 177107 115907 177108
rect 116945 177107 117011 177108
rect 124949 177107 125015 177110
rect 148174 177108 148180 177110
rect 148244 177108 148291 177112
rect 148225 177107 148291 177108
rect 101990 176972 101996 177036
rect 102060 177034 102066 177036
rect 167678 177034 167684 177036
rect 102060 176974 167684 177034
rect 102060 176972 102066 176974
rect 167678 176972 167684 176974
rect 167748 176972 167754 177036
rect 103278 176836 103284 176900
rect 103348 176898 103354 176900
rect 167494 176898 167500 176900
rect 103348 176838 167500 176898
rect 103348 176836 103354 176838
rect 167494 176836 167500 176838
rect 167564 176836 167570 176900
rect 97022 176700 97028 176764
rect 97092 176762 97098 176764
rect 97809 176762 97875 176765
rect 97092 176760 97875 176762
rect 97092 176704 97814 176760
rect 97870 176704 97875 176760
rect 97092 176702 97875 176704
rect 97092 176700 97098 176702
rect 97809 176699 97875 176702
rect 98310 176700 98316 176764
rect 98380 176762 98386 176764
rect 99189 176762 99255 176765
rect 100753 176764 100819 176765
rect 108113 176764 108179 176765
rect 100702 176762 100708 176764
rect 98380 176760 99255 176762
rect 98380 176704 99194 176760
rect 99250 176704 99255 176760
rect 98380 176702 99255 176704
rect 100662 176702 100708 176762
rect 100772 176760 100819 176764
rect 108062 176762 108068 176764
rect 100814 176704 100819 176760
rect 98380 176700 98386 176702
rect 99189 176699 99255 176702
rect 100702 176700 100708 176702
rect 100772 176700 100819 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 110045 176762 110111 176765
rect 118417 176764 118483 176765
rect 125777 176764 125843 176765
rect 118366 176762 118372 176764
rect 109604 176760 110111 176762
rect 109604 176704 110050 176760
rect 110106 176704 110111 176760
rect 109604 176702 110111 176704
rect 118326 176702 118372 176762
rect 118436 176760 118483 176764
rect 125726 176762 125732 176764
rect 118478 176704 118483 176760
rect 109604 176700 109610 176702
rect 100753 176699 100819 176700
rect 108113 176699 108179 176700
rect 110045 176699 110111 176702
rect 118366 176700 118372 176702
rect 118436 176700 118483 176704
rect 125686 176702 125732 176762
rect 125796 176760 125843 176764
rect 128169 176762 128235 176765
rect 130745 176764 130811 176765
rect 132033 176764 132099 176765
rect 134425 176764 134491 176765
rect 135713 176764 135779 176765
rect 130694 176762 130700 176764
rect 125838 176704 125843 176760
rect 125726 176700 125732 176702
rect 125796 176700 125843 176704
rect 118417 176699 118483 176700
rect 125777 176699 125843 176700
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 130654 176702 130700 176762
rect 130764 176760 130811 176764
rect 131982 176762 131988 176764
rect 130806 176704 130811 176760
rect 130694 176700 130700 176702
rect 130764 176700 130811 176704
rect 131942 176702 131988 176762
rect 132052 176760 132099 176764
rect 134374 176762 134380 176764
rect 132094 176704 132099 176760
rect 131982 176700 131988 176702
rect 132052 176700 132099 176704
rect 134334 176702 134380 176762
rect 134444 176760 134491 176764
rect 135662 176762 135668 176764
rect 134486 176704 134491 176760
rect 134374 176700 134380 176702
rect 134444 176700 134491 176704
rect 135622 176702 135668 176762
rect 135732 176760 135779 176764
rect 135774 176704 135779 176760
rect 135662 176700 135668 176702
rect 135732 176700 135779 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 159265 176762 159331 176765
rect 158916 176760 159331 176762
rect 158916 176704 159270 176760
rect 159326 176704 159331 176760
rect 158916 176702 159331 176704
rect 158916 176700 158922 176702
rect 130745 176699 130811 176700
rect 132033 176699 132099 176700
rect 134425 176699 134491 176700
rect 135713 176699 135779 176700
rect 159265 176699 159331 176702
rect 128126 176492 128186 176699
rect 260966 176564 260972 176628
rect 261036 176626 261042 176628
rect 261201 176626 261267 176629
rect 261036 176624 261267 176626
rect 261036 176568 261206 176624
rect 261262 176568 261267 176624
rect 261036 176566 261267 176568
rect 261036 176564 261042 176566
rect 261201 176563 261267 176566
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 318149 176218 318215 176221
rect 327206 176218 327212 176220
rect 318149 176216 327212 176218
rect 318149 176160 318154 176216
rect 318210 176160 327212 176216
rect 318149 176158 327212 176160
rect 318149 176155 318215 176158
rect 327206 176156 327212 176158
rect 327276 176156 327282 176220
rect 162117 176082 162183 176085
rect 249977 176082 250043 176085
rect 162117 176080 250043 176082
rect -960 175796 480 176036
rect 162117 176024 162122 176080
rect 162178 176024 249982 176080
rect 250038 176024 250043 176080
rect 162117 176022 250043 176024
rect 162117 176019 162183 176022
rect 249977 176019 250043 176022
rect 321461 176082 321527 176085
rect 321461 176080 321570 176082
rect 321461 176024 321466 176080
rect 321522 176024 321570 176080
rect 321461 176019 321570 176024
rect 69013 175946 69079 175949
rect 254526 175946 254532 175948
rect 69013 175944 254532 175946
rect 69013 175888 69018 175944
rect 69074 175888 254532 175944
rect 69013 175886 254532 175888
rect 69013 175883 69079 175886
rect 254526 175884 254532 175886
rect 254596 175884 254602 175948
rect 265014 175884 265020 175948
rect 265084 175946 265090 175948
rect 266261 175946 266327 175949
rect 265084 175944 266327 175946
rect 265084 175888 266266 175944
rect 266322 175888 266327 175944
rect 265084 175886 266327 175888
rect 265084 175884 265090 175886
rect 266261 175883 266327 175886
rect 246941 175810 247007 175813
rect 246941 175808 248338 175810
rect 246941 175752 246946 175808
rect 247002 175752 248338 175808
rect 246941 175750 248338 175752
rect 246941 175747 247007 175750
rect 213913 175674 213979 175677
rect 213913 175672 217212 175674
rect 213913 175616 213918 175672
rect 213974 175616 217212 175672
rect 248278 175644 248338 175750
rect 307661 175674 307727 175677
rect 307661 175672 310132 175674
rect 213913 175614 217212 175616
rect 307661 175616 307666 175672
rect 307722 175616 310132 175672
rect 307661 175614 310132 175616
rect 213913 175611 213979 175614
rect 307661 175611 307727 175614
rect 321510 175508 321570 176019
rect 104617 175404 104683 175405
rect 121913 175404 121979 175405
rect 129457 175404 129523 175405
rect 133137 175404 133203 175405
rect 104566 175402 104572 175404
rect 104526 175342 104572 175402
rect 104636 175400 104683 175404
rect 121862 175402 121868 175404
rect 104678 175344 104683 175400
rect 104566 175340 104572 175342
rect 104636 175340 104683 175344
rect 121822 175342 121868 175402
rect 121932 175400 121979 175404
rect 129406 175402 129412 175404
rect 121974 175344 121979 175400
rect 121862 175340 121868 175342
rect 121932 175340 121979 175344
rect 129366 175342 129412 175402
rect 129476 175400 129523 175404
rect 133086 175402 133092 175404
rect 129518 175344 129523 175400
rect 129406 175340 129412 175342
rect 129476 175340 129523 175344
rect 133046 175342 133092 175402
rect 133156 175400 133203 175404
rect 133198 175344 133203 175400
rect 133086 175340 133092 175342
rect 133156 175340 133203 175344
rect 104617 175339 104683 175340
rect 121913 175339 121979 175340
rect 129457 175339 129523 175340
rect 133137 175339 133203 175340
rect 249241 175266 249307 175269
rect 248860 175264 249307 175266
rect 248860 175208 249246 175264
rect 249302 175208 249307 175264
rect 248860 175206 249307 175208
rect 249241 175203 249307 175206
rect 307017 175266 307083 175269
rect 307017 175264 310132 175266
rect 307017 175208 307022 175264
rect 307078 175208 310132 175264
rect 307017 175206 310132 175208
rect 307017 175203 307083 175206
rect 119429 174996 119495 174997
rect 119392 174994 119398 174996
rect 119338 174934 119398 174994
rect 119462 174992 119495 174996
rect 119490 174936 119495 174992
rect 119392 174932 119398 174934
rect 119462 174932 119495 174936
rect 119429 174931 119495 174932
rect 213913 174994 213979 174997
rect 213913 174992 217212 174994
rect 213913 174936 213918 174992
rect 213974 174936 217212 174992
rect 213913 174934 217212 174936
rect 213913 174931 213979 174934
rect 307477 174858 307543 174861
rect 307477 174856 310132 174858
rect 307477 174800 307482 174856
rect 307538 174800 310132 174856
rect 307477 174798 310132 174800
rect 307477 174795 307543 174798
rect 249190 174722 249196 174724
rect 248860 174662 249196 174722
rect 249190 174660 249196 174662
rect 249260 174660 249266 174724
rect 324589 174722 324655 174725
rect 321908 174720 324655 174722
rect 321908 174664 324594 174720
rect 324650 174664 324655 174720
rect 321908 174662 324655 174664
rect 324589 174659 324655 174662
rect 265566 174524 265572 174588
rect 265636 174586 265642 174588
rect 285581 174586 285647 174589
rect 265636 174584 285647 174586
rect 265636 174528 285586 174584
rect 285642 174528 285647 174584
rect 265636 174526 285647 174528
rect 265636 174524 265642 174526
rect 285581 174523 285647 174526
rect 342846 174524 342852 174588
rect 342916 174586 342922 174588
rect 398097 174586 398163 174589
rect 533654 174586 533660 174588
rect 342916 174584 533660 174586
rect 342916 174528 398102 174584
rect 398158 174528 533660 174584
rect 342916 174526 533660 174528
rect 342916 174524 342922 174526
rect 398097 174523 398163 174526
rect 533654 174524 533660 174526
rect 533724 174524 533730 174588
rect 307569 174450 307635 174453
rect 307569 174448 310132 174450
rect 307569 174392 307574 174448
rect 307630 174392 310132 174448
rect 307569 174390 310132 174392
rect 307569 174387 307635 174390
rect 321318 174388 321324 174452
rect 321388 174388 321394 174452
rect 214005 174314 214071 174317
rect 249742 174314 249748 174316
rect 214005 174312 217212 174314
rect 214005 174256 214010 174312
rect 214066 174256 217212 174312
rect 214005 174254 217212 174256
rect 248860 174254 249748 174314
rect 214005 174251 214071 174254
rect 249742 174252 249748 174254
rect 249812 174252 249818 174316
rect 307661 174042 307727 174045
rect 307661 174040 310132 174042
rect 307661 173984 307666 174040
rect 307722 173984 310132 174040
rect 321326 174012 321386 174388
rect 307661 173982 310132 173984
rect 307661 173979 307727 173982
rect 249977 173770 250043 173773
rect 248860 173768 250043 173770
rect 248860 173712 249982 173768
rect 250038 173712 250043 173768
rect 248860 173710 250043 173712
rect 249977 173707 250043 173710
rect 213913 173634 213979 173637
rect 307661 173634 307727 173637
rect 213913 173632 217212 173634
rect 213913 173576 213918 173632
rect 213974 173576 217212 173632
rect 213913 173574 217212 173576
rect 307661 173632 310132 173634
rect 307661 173576 307666 173632
rect 307722 173576 310132 173632
rect 307661 173574 310132 173576
rect 213913 173571 213979 173574
rect 307661 173571 307727 173574
rect 252502 173362 252508 173364
rect 248860 173302 252508 173362
rect 252502 173300 252508 173302
rect 252572 173300 252578 173364
rect 306925 173226 306991 173229
rect 326654 173226 326660 173228
rect 306925 173224 310132 173226
rect 306925 173168 306930 173224
rect 306986 173168 310132 173224
rect 306925 173166 310132 173168
rect 321908 173166 326660 173226
rect 306925 173163 306991 173166
rect 326654 173164 326660 173166
rect 326724 173164 326730 173228
rect 214097 172954 214163 172957
rect 214097 172952 217212 172954
rect 214097 172896 214102 172952
rect 214158 172896 217212 172952
rect 214097 172894 217212 172896
rect 214097 172891 214163 172894
rect 249190 172818 249196 172820
rect 248860 172758 249196 172818
rect 249190 172756 249196 172758
rect 249260 172756 249266 172820
rect 307293 172682 307359 172685
rect 307293 172680 310132 172682
rect 307293 172624 307298 172680
rect 307354 172624 310132 172680
rect 307293 172622 310132 172624
rect 307293 172619 307359 172622
rect 249057 172546 249123 172549
rect 249057 172544 249258 172546
rect 249057 172488 249062 172544
rect 249118 172488 249258 172544
rect 249057 172486 249258 172488
rect 249057 172483 249123 172486
rect 249198 172410 249258 172486
rect 324313 172410 324379 172413
rect 248860 172350 249258 172410
rect 321908 172408 324379 172410
rect 321908 172352 324318 172408
rect 324374 172352 324379 172408
rect 321908 172350 324379 172352
rect 324313 172347 324379 172350
rect 213913 172274 213979 172277
rect 307569 172274 307635 172277
rect 213913 172272 217212 172274
rect 213913 172216 213918 172272
rect 213974 172216 217212 172272
rect 213913 172214 217212 172216
rect 307569 172272 310132 172274
rect 307569 172216 307574 172272
rect 307630 172216 310132 172272
rect 307569 172214 310132 172216
rect 213913 172211 213979 172214
rect 307569 172211 307635 172214
rect 249149 171866 249215 171869
rect 248860 171864 249215 171866
rect 248860 171808 249154 171864
rect 249210 171808 249215 171864
rect 248860 171806 249215 171808
rect 249149 171803 249215 171806
rect 307661 171866 307727 171869
rect 307661 171864 310132 171866
rect 307661 171808 307666 171864
rect 307722 171808 310132 171864
rect 307661 171806 310132 171808
rect 307661 171803 307727 171806
rect 325785 171730 325851 171733
rect 321908 171728 325851 171730
rect 321908 171672 325790 171728
rect 325846 171672 325851 171728
rect 321908 171670 325851 171672
rect 325785 171667 325851 171670
rect 168005 171594 168071 171597
rect 164694 171592 168071 171594
rect 164694 171536 168010 171592
rect 168066 171536 168071 171592
rect 164694 171534 168071 171536
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 168005 171531 168071 171534
rect 214005 171594 214071 171597
rect 214005 171592 217212 171594
rect 214005 171536 214010 171592
rect 214066 171536 217212 171592
rect 214005 171534 217212 171536
rect 214005 171531 214071 171534
rect 249333 171458 249399 171461
rect 248860 171456 249399 171458
rect 248860 171400 249338 171456
rect 249394 171400 249399 171456
rect 248860 171398 249399 171400
rect 249333 171395 249399 171398
rect 307477 171458 307543 171461
rect 307477 171456 310132 171458
rect 307477 171400 307482 171456
rect 307538 171400 310132 171456
rect 307477 171398 310132 171400
rect 307477 171395 307543 171398
rect 213913 171050 213979 171053
rect 307293 171050 307359 171053
rect 213913 171048 217212 171050
rect 213913 170992 213918 171048
rect 213974 170992 217212 171048
rect 213913 170990 217212 170992
rect 307293 171048 310132 171050
rect 307293 170992 307298 171048
rect 307354 170992 310132 171048
rect 307293 170990 310132 170992
rect 213913 170987 213979 170990
rect 307293 170987 307359 170990
rect 250069 170914 250135 170917
rect 327206 170914 327212 170916
rect 248860 170912 250135 170914
rect 248860 170856 250074 170912
rect 250130 170856 250135 170912
rect 248860 170854 250135 170856
rect 321908 170854 327212 170914
rect 250069 170851 250135 170854
rect 327206 170852 327212 170854
rect 327276 170852 327282 170916
rect 306557 170642 306623 170645
rect 306557 170640 310132 170642
rect 306557 170584 306562 170640
rect 306618 170584 310132 170640
rect 306557 170582 310132 170584
rect 306557 170579 306623 170582
rect 252461 170506 252527 170509
rect 248860 170504 252527 170506
rect 248860 170448 252466 170504
rect 252522 170448 252527 170504
rect 248860 170446 252527 170448
rect 252461 170443 252527 170446
rect 214925 170370 214991 170373
rect 214925 170368 217212 170370
rect 214925 170312 214930 170368
rect 214986 170312 217212 170368
rect 214925 170310 217212 170312
rect 214925 170307 214991 170310
rect 307661 170234 307727 170237
rect 307661 170232 310132 170234
rect 307661 170176 307666 170232
rect 307722 170176 310132 170232
rect 307661 170174 310132 170176
rect 307661 170171 307727 170174
rect 259678 170098 259684 170100
rect 248860 170038 259684 170098
rect 259678 170036 259684 170038
rect 259748 170036 259754 170100
rect 324313 170098 324379 170101
rect 321908 170096 324379 170098
rect 321908 170040 324318 170096
rect 324374 170040 324379 170096
rect 321908 170038 324379 170040
rect 324313 170035 324379 170038
rect 307661 169826 307727 169829
rect 307661 169824 310132 169826
rect 307661 169768 307666 169824
rect 307722 169768 310132 169824
rect 307661 169766 310132 169768
rect 307661 169763 307727 169766
rect 213913 169690 213979 169693
rect 213913 169688 217212 169690
rect 213913 169632 213918 169688
rect 213974 169632 217212 169688
rect 213913 169630 217212 169632
rect 213913 169627 213979 169630
rect 252737 169554 252803 169557
rect 248860 169552 252803 169554
rect 248860 169496 252742 169552
rect 252798 169496 252803 169552
rect 248860 169494 252803 169496
rect 252737 169491 252803 169494
rect 324313 169418 324379 169421
rect 321908 169416 324379 169418
rect 321908 169360 324318 169416
rect 324374 169360 324379 169416
rect 321908 169358 324379 169360
rect 324313 169355 324379 169358
rect 306557 169282 306623 169285
rect 306557 169280 310132 169282
rect 306557 169224 306562 169280
rect 306618 169224 310132 169280
rect 306557 169222 310132 169224
rect 306557 169219 306623 169222
rect 252461 169146 252527 169149
rect 248860 169144 252527 169146
rect 248860 169088 252466 169144
rect 252522 169088 252527 169144
rect 248860 169086 252527 169088
rect 252461 169083 252527 169086
rect 214005 169010 214071 169013
rect 214005 169008 217212 169010
rect 214005 168952 214010 169008
rect 214066 168952 217212 169008
rect 214005 168950 217212 168952
rect 214005 168947 214071 168950
rect 307661 168874 307727 168877
rect 307661 168872 310132 168874
rect 307661 168816 307666 168872
rect 307722 168816 310132 168872
rect 307661 168814 310132 168816
rect 307661 168811 307727 168814
rect 252369 168602 252435 168605
rect 324405 168602 324471 168605
rect 248860 168600 252435 168602
rect 248860 168544 252374 168600
rect 252430 168544 252435 168600
rect 248860 168542 252435 168544
rect 321908 168600 324471 168602
rect 321908 168544 324410 168600
rect 324466 168544 324471 168600
rect 321908 168542 324471 168544
rect 252369 168539 252435 168542
rect 324405 168539 324471 168542
rect 307293 168466 307359 168469
rect 307293 168464 310132 168466
rect 307293 168408 307298 168464
rect 307354 168408 310132 168464
rect 307293 168406 310132 168408
rect 307293 168403 307359 168406
rect 213913 168330 213979 168333
rect 213913 168328 217212 168330
rect 213913 168272 213918 168328
rect 213974 168272 217212 168328
rect 213913 168270 217212 168272
rect 213913 168267 213979 168270
rect 252461 168194 252527 168197
rect 248860 168192 252527 168194
rect 248860 168136 252466 168192
rect 252522 168136 252527 168192
rect 248860 168134 252527 168136
rect 252461 168131 252527 168134
rect 307477 168058 307543 168061
rect 307477 168056 310132 168058
rect 307477 168000 307482 168056
rect 307538 168000 310132 168056
rect 307477 167998 310132 168000
rect 307477 167995 307543 167998
rect 324313 167786 324379 167789
rect 321908 167784 324379 167786
rect 321908 167728 324318 167784
rect 324374 167728 324379 167784
rect 321908 167726 324379 167728
rect 324313 167723 324379 167726
rect 214005 167650 214071 167653
rect 252369 167650 252435 167653
rect 214005 167648 217212 167650
rect 214005 167592 214010 167648
rect 214066 167592 217212 167648
rect 214005 167590 217212 167592
rect 248860 167648 252435 167650
rect 248860 167592 252374 167648
rect 252430 167592 252435 167648
rect 248860 167590 252435 167592
rect 214005 167587 214071 167590
rect 252369 167587 252435 167590
rect 307569 167650 307635 167653
rect 307569 167648 310132 167650
rect 307569 167592 307574 167648
rect 307630 167592 310132 167648
rect 307569 167590 310132 167592
rect 307569 167587 307635 167590
rect 252001 167242 252067 167245
rect 248860 167240 252067 167242
rect 248860 167184 252006 167240
rect 252062 167184 252067 167240
rect 248860 167182 252067 167184
rect 252001 167179 252067 167182
rect 307661 167242 307727 167245
rect 307661 167240 310132 167242
rect 307661 167184 307666 167240
rect 307722 167184 310132 167240
rect 307661 167182 310132 167184
rect 307661 167179 307727 167182
rect 335854 167106 335860 167108
rect 321908 167046 335860 167106
rect 335854 167044 335860 167046
rect 335924 167044 335930 167108
rect 213913 166970 213979 166973
rect 213913 166968 217212 166970
rect 213913 166912 213918 166968
rect 213974 166912 217212 166968
rect 213913 166910 217212 166912
rect 213913 166907 213979 166910
rect 306557 166834 306623 166837
rect 306557 166832 310132 166834
rect 306557 166776 306562 166832
rect 306618 166776 310132 166832
rect 306557 166774 310132 166776
rect 306557 166771 306623 166774
rect 252461 166698 252527 166701
rect 248860 166696 252527 166698
rect 248860 166640 252466 166696
rect 252522 166640 252527 166696
rect 248860 166638 252527 166640
rect 252461 166635 252527 166638
rect 214097 166426 214163 166429
rect 306373 166426 306439 166429
rect 214097 166424 217212 166426
rect 214097 166368 214102 166424
rect 214158 166368 217212 166424
rect 214097 166366 217212 166368
rect 306373 166424 310132 166426
rect 306373 166368 306378 166424
rect 306434 166368 310132 166424
rect 306373 166366 310132 166368
rect 214097 166363 214163 166366
rect 306373 166363 306439 166366
rect 251909 166290 251975 166293
rect 327022 166290 327028 166292
rect 248860 166288 251975 166290
rect 248860 166232 251914 166288
rect 251970 166232 251975 166288
rect 248860 166230 251975 166232
rect 321908 166230 327028 166290
rect 251909 166227 251975 166230
rect 327022 166228 327028 166230
rect 327092 166228 327098 166292
rect 306465 165882 306531 165885
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 306465 165880 310132 165882
rect 306465 165824 306470 165880
rect 306526 165824 310132 165880
rect 306465 165822 310132 165824
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 306465 165819 306531 165822
rect 580165 165819 580231 165822
rect 214005 165746 214071 165749
rect 252369 165746 252435 165749
rect 214005 165744 217212 165746
rect 214005 165688 214010 165744
rect 214066 165688 217212 165744
rect 214005 165686 217212 165688
rect 248860 165744 252435 165746
rect 248860 165688 252374 165744
rect 252430 165688 252435 165744
rect 583520 165732 584960 165822
rect 248860 165686 252435 165688
rect 214005 165683 214071 165686
rect 252369 165683 252435 165686
rect 306465 165474 306531 165477
rect 324313 165474 324379 165477
rect 306465 165472 310132 165474
rect 306465 165416 306470 165472
rect 306526 165416 310132 165472
rect 306465 165414 310132 165416
rect 321908 165472 324379 165474
rect 321908 165416 324318 165472
rect 324374 165416 324379 165472
rect 321908 165414 324379 165416
rect 306465 165411 306531 165414
rect 324313 165411 324379 165414
rect 252461 165338 252527 165341
rect 248860 165336 252527 165338
rect 248860 165280 252466 165336
rect 252522 165280 252527 165336
rect 248860 165278 252527 165280
rect 252461 165275 252527 165278
rect 213913 165066 213979 165069
rect 307109 165066 307175 165069
rect 321277 165066 321343 165069
rect 213913 165064 217212 165066
rect 213913 165008 213918 165064
rect 213974 165008 217212 165064
rect 213913 165006 217212 165008
rect 307109 165064 310132 165066
rect 307109 165008 307114 165064
rect 307170 165008 310132 165064
rect 307109 165006 310132 165008
rect 321277 165064 321386 165066
rect 321277 165008 321282 165064
rect 321338 165008 321386 165064
rect 213913 165003 213979 165006
rect 307109 165003 307175 165006
rect 321277 165003 321386 165008
rect 251909 164794 251975 164797
rect 248860 164792 251975 164794
rect 248860 164736 251914 164792
rect 251970 164736 251975 164792
rect 321326 164764 321386 165003
rect 248860 164734 251975 164736
rect 251909 164731 251975 164734
rect 306373 164658 306439 164661
rect 306373 164656 310132 164658
rect 306373 164600 306378 164656
rect 306434 164600 310132 164656
rect 306373 164598 310132 164600
rect 306373 164595 306439 164598
rect 166206 164324 166212 164388
rect 166276 164386 166282 164388
rect 251449 164386 251515 164389
rect 166276 164326 217212 164386
rect 248860 164384 251515 164386
rect 248860 164328 251454 164384
rect 251510 164328 251515 164384
rect 248860 164326 251515 164328
rect 166276 164324 166282 164326
rect 251449 164323 251515 164326
rect 306373 164250 306439 164253
rect 306373 164248 310132 164250
rect 306373 164192 306378 164248
rect 306434 164192 310132 164248
rect 306373 164190 310132 164192
rect 306373 164187 306439 164190
rect 263726 163978 263732 163980
rect 248860 163918 263732 163978
rect 263726 163916 263732 163918
rect 263796 163916 263802 163980
rect 324313 163978 324379 163981
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 324313 163915 324379 163918
rect 306557 163842 306623 163845
rect 306557 163840 310132 163842
rect 306557 163784 306562 163840
rect 306618 163784 310132 163840
rect 306557 163782 310132 163784
rect 306557 163779 306623 163782
rect 213913 163706 213979 163709
rect 213913 163704 217212 163706
rect 213913 163648 213918 163704
rect 213974 163648 217212 163704
rect 213913 163646 217212 163648
rect 213913 163643 213979 163646
rect 251909 163434 251975 163437
rect 248860 163432 251975 163434
rect 248860 163376 251914 163432
rect 251970 163376 251975 163432
rect 248860 163374 251975 163376
rect 251909 163371 251975 163374
rect 306373 163434 306439 163437
rect 306373 163432 310132 163434
rect 306373 163376 306378 163432
rect 306434 163376 310132 163432
rect 306373 163374 310132 163376
rect 306373 163371 306439 163374
rect 324405 163162 324471 163165
rect 321908 163160 324471 163162
rect 321908 163104 324410 163160
rect 324466 163104 324471 163160
rect 321908 163102 324471 163104
rect 324405 163099 324471 163102
rect 214005 163026 214071 163029
rect 252185 163026 252251 163029
rect 214005 163024 217212 163026
rect 214005 162968 214010 163024
rect 214066 162968 217212 163024
rect 214005 162966 217212 162968
rect 248860 163024 252251 163026
rect 248860 162968 252190 163024
rect 252246 162968 252251 163024
rect 248860 162966 252251 162968
rect 214005 162963 214071 162966
rect 252185 162963 252251 162966
rect 306465 163026 306531 163029
rect 306465 163024 310132 163026
rect 306465 162968 306470 163024
rect 306526 162968 310132 163024
rect 306465 162966 310132 162968
rect 306465 162963 306531 162966
rect 252093 162482 252159 162485
rect 248860 162480 252159 162482
rect 248860 162424 252098 162480
rect 252154 162424 252159 162480
rect 248860 162422 252159 162424
rect 252093 162419 252159 162422
rect 306465 162482 306531 162485
rect 306465 162480 310132 162482
rect 306465 162424 306470 162480
rect 306526 162424 310132 162480
rect 306465 162422 310132 162424
rect 306465 162419 306531 162422
rect 217182 161938 217242 162316
rect 252461 162074 252527 162077
rect 248860 162072 252527 162074
rect 248860 162016 252466 162072
rect 252522 162016 252527 162072
rect 248860 162014 252527 162016
rect 252461 162011 252527 162014
rect 306557 162074 306623 162077
rect 306557 162072 310132 162074
rect 306557 162016 306562 162072
rect 306618 162016 310132 162072
rect 306557 162014 310132 162016
rect 306557 162011 306623 162014
rect 200070 161878 217242 161938
rect 166390 161468 166396 161532
rect 166460 161530 166466 161532
rect 200070 161530 200130 161878
rect 213913 161802 213979 161805
rect 321878 161802 321938 162452
rect 328678 161802 328684 161804
rect 213913 161800 217212 161802
rect 213913 161744 213918 161800
rect 213974 161744 217212 161800
rect 213913 161742 217212 161744
rect 321878 161742 328684 161802
rect 213913 161739 213979 161742
rect 328678 161740 328684 161742
rect 328748 161740 328754 161804
rect 306373 161666 306439 161669
rect 325877 161666 325943 161669
rect 306373 161664 310132 161666
rect 306373 161608 306378 161664
rect 306434 161608 310132 161664
rect 306373 161606 310132 161608
rect 321908 161664 325943 161666
rect 321908 161608 325882 161664
rect 325938 161608 325943 161664
rect 321908 161606 325943 161608
rect 306373 161603 306439 161606
rect 325877 161603 325943 161606
rect 252461 161530 252527 161533
rect 166460 161470 200130 161530
rect 248860 161528 252527 161530
rect 248860 161472 252466 161528
rect 252522 161472 252527 161528
rect 248860 161470 252527 161472
rect 166460 161468 166466 161470
rect 252461 161467 252527 161470
rect 306465 161258 306531 161261
rect 306465 161256 310132 161258
rect 306465 161200 306470 161256
rect 306526 161200 310132 161256
rect 306465 161198 310132 161200
rect 306465 161195 306531 161198
rect 213913 161122 213979 161125
rect 252461 161122 252527 161125
rect 213913 161120 217212 161122
rect 213913 161064 213918 161120
rect 213974 161064 217212 161120
rect 213913 161062 217212 161064
rect 248860 161120 252527 161122
rect 248860 161064 252466 161120
rect 252522 161064 252527 161120
rect 248860 161062 252527 161064
rect 213913 161059 213979 161062
rect 252461 161059 252527 161062
rect 306373 160850 306439 160853
rect 324313 160850 324379 160853
rect 306373 160848 310132 160850
rect 306373 160792 306378 160848
rect 306434 160792 310132 160848
rect 306373 160790 310132 160792
rect 321908 160848 324379 160850
rect 321908 160792 324318 160848
rect 324374 160792 324379 160848
rect 321908 160790 324379 160792
rect 306373 160787 306439 160790
rect 324313 160787 324379 160790
rect 259310 160652 259316 160716
rect 259380 160714 259386 160716
rect 269062 160714 269068 160716
rect 259380 160654 269068 160714
rect 259380 160652 259386 160654
rect 269062 160652 269068 160654
rect 269132 160652 269138 160716
rect 251357 160578 251423 160581
rect 248860 160576 251423 160578
rect 248860 160520 251362 160576
rect 251418 160520 251423 160576
rect 248860 160518 251423 160520
rect 251357 160515 251423 160518
rect 214005 160442 214071 160445
rect 306557 160442 306623 160445
rect 214005 160440 217212 160442
rect 214005 160384 214010 160440
rect 214066 160384 217212 160440
rect 214005 160382 217212 160384
rect 306557 160440 310132 160442
rect 306557 160384 306562 160440
rect 306618 160384 310132 160440
rect 306557 160382 310132 160384
rect 214005 160379 214071 160382
rect 306557 160379 306623 160382
rect 251909 160170 251975 160173
rect 324497 160170 324563 160173
rect 248860 160168 251975 160170
rect 248860 160112 251914 160168
rect 251970 160112 251975 160168
rect 248860 160110 251975 160112
rect 321908 160168 324563 160170
rect 321908 160112 324502 160168
rect 324558 160112 324563 160168
rect 321908 160110 324563 160112
rect 251909 160107 251975 160110
rect 324497 160107 324563 160110
rect 306557 160034 306623 160037
rect 306557 160032 310132 160034
rect 306557 159976 306562 160032
rect 306618 159976 310132 160032
rect 306557 159974 310132 159976
rect 306557 159971 306623 159974
rect 337878 159972 337884 160036
rect 337948 160034 337954 160036
rect 535494 160034 535500 160036
rect 337948 159974 535500 160034
rect 337948 159972 337954 159974
rect 535494 159972 535500 159974
rect 535564 159972 535570 160036
rect 213913 159762 213979 159765
rect 213913 159760 217212 159762
rect 213913 159704 213918 159760
rect 213974 159704 217212 159760
rect 213913 159702 217212 159704
rect 213913 159699 213979 159702
rect 251173 159626 251239 159629
rect 248860 159624 251239 159626
rect 248860 159568 251178 159624
rect 251234 159568 251239 159624
rect 248860 159566 251239 159568
rect 251173 159563 251239 159566
rect 306373 159626 306439 159629
rect 306373 159624 310132 159626
rect 306373 159568 306378 159624
rect 306434 159568 310132 159624
rect 306373 159566 310132 159568
rect 306373 159563 306439 159566
rect 324313 159354 324379 159357
rect 321908 159352 324379 159354
rect 321908 159296 324318 159352
rect 324374 159296 324379 159352
rect 321908 159294 324379 159296
rect 324313 159291 324379 159294
rect 251633 159218 251699 159221
rect 248860 159216 251699 159218
rect 248860 159160 251638 159216
rect 251694 159160 251699 159216
rect 248860 159158 251699 159160
rect 251633 159155 251699 159158
rect 214005 159082 214071 159085
rect 306465 159082 306531 159085
rect 214005 159080 217212 159082
rect 214005 159024 214010 159080
rect 214066 159024 217212 159080
rect 214005 159022 217212 159024
rect 306465 159080 310132 159082
rect 306465 159024 306470 159080
rect 306526 159024 310132 159080
rect 306465 159022 310132 159024
rect 214005 159019 214071 159022
rect 306465 159019 306531 159022
rect 256734 158810 256740 158812
rect 248860 158750 256740 158810
rect 256734 158748 256740 158750
rect 256804 158748 256810 158812
rect 337469 158810 337535 158813
rect 337878 158810 337884 158812
rect 337469 158808 337884 158810
rect 337469 158752 337474 158808
rect 337530 158752 337884 158808
rect 337469 158750 337884 158752
rect 337469 158747 337535 158750
rect 337878 158748 337884 158750
rect 337948 158748 337954 158812
rect 306557 158674 306623 158677
rect 306557 158672 310132 158674
rect 306557 158616 306562 158672
rect 306618 158616 310132 158672
rect 306557 158614 310132 158616
rect 306557 158611 306623 158614
rect 324313 158538 324379 158541
rect 321908 158536 324379 158538
rect 321908 158480 324318 158536
rect 324374 158480 324379 158536
rect 321908 158478 324379 158480
rect 324313 158475 324379 158478
rect 213453 157858 213519 157861
rect 217182 157858 217242 158372
rect 252461 158266 252527 158269
rect 248860 158264 252527 158266
rect 248860 158208 252466 158264
rect 252522 158208 252527 158264
rect 248860 158206 252527 158208
rect 252461 158203 252527 158206
rect 306373 158266 306439 158269
rect 306373 158264 310132 158266
rect 306373 158208 306378 158264
rect 306434 158208 310132 158264
rect 306373 158206 310132 158208
rect 306373 158203 306439 158206
rect 252369 157858 252435 157861
rect 213453 157856 217242 157858
rect 213453 157800 213458 157856
rect 213514 157800 217242 157856
rect 213453 157798 217242 157800
rect 248860 157856 252435 157858
rect 248860 157800 252374 157856
rect 252430 157800 252435 157856
rect 248860 157798 252435 157800
rect 213453 157795 213519 157798
rect 252369 157795 252435 157798
rect 306465 157858 306531 157861
rect 324405 157858 324471 157861
rect 306465 157856 310132 157858
rect 306465 157800 306470 157856
rect 306526 157800 310132 157856
rect 306465 157798 310132 157800
rect 321908 157856 324471 157858
rect 321908 157800 324410 157856
rect 324466 157800 324471 157856
rect 321908 157798 324471 157800
rect 306465 157795 306531 157798
rect 324405 157795 324471 157798
rect 200070 157662 217212 157722
rect 167678 157524 167684 157588
rect 167748 157586 167754 157588
rect 200070 157586 200130 157662
rect 167748 157526 200130 157586
rect 167748 157524 167754 157526
rect 167494 157388 167500 157452
rect 167564 157450 167570 157452
rect 213453 157450 213519 157453
rect 167564 157448 213519 157450
rect 167564 157392 213458 157448
rect 213514 157392 213519 157448
rect 167564 157390 213519 157392
rect 167564 157388 167570 157390
rect 213453 157387 213519 157390
rect 306925 157450 306991 157453
rect 306925 157448 310132 157450
rect 306925 157392 306930 157448
rect 306986 157392 310132 157448
rect 306925 157390 310132 157392
rect 306925 157387 306991 157390
rect 255446 157314 255452 157316
rect 248860 157254 255452 157314
rect 255446 157252 255452 157254
rect 255516 157252 255522 157316
rect 214097 157178 214163 157181
rect 214097 157176 217212 157178
rect 214097 157120 214102 157176
rect 214158 157120 217212 157176
rect 214097 157118 217212 157120
rect 214097 157115 214163 157118
rect 307477 157042 307543 157045
rect 324313 157042 324379 157045
rect 307477 157040 310132 157042
rect 307477 156984 307482 157040
rect 307538 156984 310132 157040
rect 307477 156982 310132 156984
rect 321908 157040 324379 157042
rect 321908 156984 324318 157040
rect 324374 156984 324379 157040
rect 321908 156982 324379 156984
rect 307477 156979 307543 156982
rect 324313 156979 324379 156982
rect 252461 156906 252527 156909
rect 248860 156904 252527 156906
rect 248860 156848 252466 156904
rect 252522 156848 252527 156904
rect 248860 156846 252527 156848
rect 252461 156843 252527 156846
rect 307569 156634 307635 156637
rect 307569 156632 310132 156634
rect 307569 156576 307574 156632
rect 307630 156576 310132 156632
rect 307569 156574 310132 156576
rect 307569 156571 307635 156574
rect 213913 156498 213979 156501
rect 213913 156496 217212 156498
rect 213913 156440 213918 156496
rect 213974 156440 217212 156496
rect 213913 156438 217212 156440
rect 213913 156435 213979 156438
rect 251541 156362 251607 156365
rect 324405 156362 324471 156365
rect 248860 156360 251607 156362
rect 248860 156304 251546 156360
rect 251602 156304 251607 156360
rect 248860 156302 251607 156304
rect 321908 156360 324471 156362
rect 321908 156304 324410 156360
rect 324466 156304 324471 156360
rect 321908 156302 324471 156304
rect 251541 156299 251607 156302
rect 324405 156299 324471 156302
rect 307661 156226 307727 156229
rect 307661 156224 310132 156226
rect 307661 156168 307666 156224
rect 307722 156168 310132 156224
rect 307661 156166 310132 156168
rect 307661 156163 307727 156166
rect 252461 155954 252527 155957
rect 248860 155952 252527 155954
rect 248860 155896 252466 155952
rect 252522 155896 252527 155952
rect 248860 155894 252527 155896
rect 252461 155891 252527 155894
rect 213913 155818 213979 155821
rect 213913 155816 217212 155818
rect 213913 155760 213918 155816
rect 213974 155760 217212 155816
rect 213913 155758 217212 155760
rect 213913 155755 213979 155758
rect 306741 155682 306807 155685
rect 306741 155680 310132 155682
rect 306741 155624 306746 155680
rect 306802 155624 310132 155680
rect 306741 155622 310132 155624
rect 306741 155619 306807 155622
rect 324681 155546 324747 155549
rect 321908 155544 324747 155546
rect 321908 155488 324686 155544
rect 324742 155488 324747 155544
rect 321908 155486 324747 155488
rect 324681 155483 324747 155486
rect 252461 155410 252527 155413
rect 248860 155408 252527 155410
rect 248860 155352 252466 155408
rect 252522 155352 252527 155408
rect 248860 155350 252527 155352
rect 252461 155347 252527 155350
rect 307477 155274 307543 155277
rect 307477 155272 310132 155274
rect 307477 155216 307482 155272
rect 307538 155216 310132 155272
rect 307477 155214 310132 155216
rect 307477 155211 307543 155214
rect 214557 155138 214623 155141
rect 214557 155136 217212 155138
rect 214557 155080 214562 155136
rect 214618 155080 217212 155136
rect 214557 155078 217212 155080
rect 214557 155075 214623 155078
rect 252369 155002 252435 155005
rect 248860 155000 252435 155002
rect 248860 154944 252374 155000
rect 252430 154944 252435 155000
rect 248860 154942 252435 154944
rect 252369 154939 252435 154942
rect 307385 154866 307451 154869
rect 307385 154864 310132 154866
rect 307385 154808 307390 154864
rect 307446 154808 310132 154864
rect 307385 154806 310132 154808
rect 307385 154803 307451 154806
rect 324313 154730 324379 154733
rect 321908 154728 324379 154730
rect 321908 154672 324318 154728
rect 324374 154672 324379 154728
rect 321908 154670 324379 154672
rect 324313 154667 324379 154670
rect 214005 154458 214071 154461
rect 249793 154458 249859 154461
rect 214005 154456 217212 154458
rect 214005 154400 214010 154456
rect 214066 154400 217212 154456
rect 214005 154398 217212 154400
rect 248860 154456 249859 154458
rect 248860 154400 249798 154456
rect 249854 154400 249859 154456
rect 248860 154398 249859 154400
rect 214005 154395 214071 154398
rect 249793 154395 249859 154398
rect 307569 154458 307635 154461
rect 307569 154456 310132 154458
rect 307569 154400 307574 154456
rect 307630 154400 310132 154456
rect 307569 154398 310132 154400
rect 307569 154395 307635 154398
rect 251725 154050 251791 154053
rect 248860 154048 251791 154050
rect 248860 153992 251730 154048
rect 251786 153992 251791 154048
rect 248860 153990 251791 153992
rect 251725 153987 251791 153990
rect 307661 154050 307727 154053
rect 324313 154050 324379 154053
rect 307661 154048 310132 154050
rect 307661 153992 307666 154048
rect 307722 153992 310132 154048
rect 307661 153990 310132 153992
rect 321908 154048 324379 154050
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 307661 153987 307727 153990
rect 324313 153987 324379 153990
rect 213913 153778 213979 153781
rect 213913 153776 217212 153778
rect 213913 153720 213918 153776
rect 213974 153720 217212 153776
rect 213913 153718 217212 153720
rect 213913 153715 213979 153718
rect 307477 153642 307543 153645
rect 307477 153640 310132 153642
rect 307477 153584 307482 153640
rect 307538 153584 310132 153640
rect 307477 153582 310132 153584
rect 307477 153579 307543 153582
rect 251173 153506 251239 153509
rect 248860 153504 251239 153506
rect 248860 153448 251178 153504
rect 251234 153448 251239 153504
rect 248860 153446 251239 153448
rect 251173 153443 251239 153446
rect 306649 153234 306715 153237
rect 323209 153234 323275 153237
rect 306649 153232 310132 153234
rect 306649 153176 306654 153232
rect 306710 153176 310132 153232
rect 306649 153174 310132 153176
rect 321908 153232 323275 153234
rect 321908 153176 323214 153232
rect 323270 153176 323275 153232
rect 321908 153174 323275 153176
rect 306649 153171 306715 153174
rect 323209 153171 323275 153174
rect 213913 153098 213979 153101
rect 252461 153098 252527 153101
rect 213913 153096 217212 153098
rect 213913 153040 213918 153096
rect 213974 153040 217212 153096
rect 213913 153038 217212 153040
rect 248860 153096 252527 153098
rect 248860 153040 252466 153096
rect 252522 153040 252527 153096
rect 248860 153038 252527 153040
rect 213913 153035 213979 153038
rect 252461 153035 252527 153038
rect 251766 152900 251772 152964
rect 251836 152962 251842 152964
rect 257613 152962 257679 152965
rect 251836 152960 257679 152962
rect 251836 152904 257618 152960
rect 257674 152904 257679 152960
rect 251836 152902 257679 152904
rect 251836 152900 251842 152902
rect 257613 152899 257679 152902
rect 260966 152690 260972 152692
rect 248860 152630 260972 152690
rect 260966 152628 260972 152630
rect 261036 152628 261042 152692
rect 306557 152690 306623 152693
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 306557 152688 310132 152690
rect 306557 152632 306562 152688
rect 306618 152632 310132 152688
rect 306557 152630 310132 152632
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 306557 152627 306623 152630
rect 580165 152627 580231 152630
rect 214005 152554 214071 152557
rect 214005 152552 217212 152554
rect 214005 152496 214010 152552
rect 214066 152496 217212 152552
rect 583520 152540 584960 152630
rect 214005 152494 217212 152496
rect 214005 152491 214071 152494
rect 324313 152418 324379 152421
rect 321908 152416 324379 152418
rect 321908 152360 324318 152416
rect 324374 152360 324379 152416
rect 321908 152358 324379 152360
rect 324313 152355 324379 152358
rect 305729 152282 305795 152285
rect 305729 152280 310132 152282
rect 305729 152224 305734 152280
rect 305790 152224 310132 152280
rect 305729 152222 310132 152224
rect 305729 152219 305795 152222
rect 252001 152146 252067 152149
rect 248860 152144 252067 152146
rect 248860 152088 252006 152144
rect 252062 152088 252067 152144
rect 248860 152086 252067 152088
rect 252001 152083 252067 152086
rect 213913 151874 213979 151877
rect 307661 151874 307727 151877
rect 213913 151872 217212 151874
rect 213913 151816 213918 151872
rect 213974 151816 217212 151872
rect 213913 151814 217212 151816
rect 307661 151872 310132 151874
rect 307661 151816 307666 151872
rect 307722 151816 310132 151872
rect 307661 151814 310132 151816
rect 213913 151811 213979 151814
rect 307661 151811 307727 151814
rect 252461 151738 252527 151741
rect 324313 151738 324379 151741
rect 248860 151736 252527 151738
rect 248860 151680 252466 151736
rect 252522 151680 252527 151736
rect 248860 151678 252527 151680
rect 321908 151736 324379 151738
rect 321908 151680 324318 151736
rect 324374 151680 324379 151736
rect 321908 151678 324379 151680
rect 252461 151675 252527 151678
rect 324313 151675 324379 151678
rect 307477 151466 307543 151469
rect 307477 151464 310132 151466
rect 307477 151408 307482 151464
rect 307538 151408 310132 151464
rect 307477 151406 310132 151408
rect 307477 151403 307543 151406
rect 214005 151194 214071 151197
rect 252645 151194 252711 151197
rect 214005 151192 217212 151194
rect 214005 151136 214010 151192
rect 214066 151136 217212 151192
rect 214005 151134 217212 151136
rect 248860 151192 252711 151194
rect 248860 151136 252650 151192
rect 252706 151136 252711 151192
rect 248860 151134 252711 151136
rect 214005 151131 214071 151134
rect 252645 151131 252711 151134
rect 307293 151058 307359 151061
rect 307293 151056 310132 151058
rect 307293 151000 307298 151056
rect 307354 151000 310132 151056
rect 307293 150998 310132 151000
rect 307293 150995 307359 150998
rect 329046 150996 329052 151060
rect 329116 151058 329122 151060
rect 343817 151058 343883 151061
rect 329116 151056 343883 151058
rect 329116 151000 343822 151056
rect 343878 151000 343883 151056
rect 329116 150998 343883 151000
rect 329116 150996 329122 150998
rect 343817 150995 343883 150998
rect 324313 150922 324379 150925
rect 321908 150920 324379 150922
rect 321908 150864 324318 150920
rect 324374 150864 324379 150920
rect 321908 150862 324379 150864
rect 324313 150859 324379 150862
rect 252369 150786 252435 150789
rect 248860 150784 252435 150786
rect 248860 150728 252374 150784
rect 252430 150728 252435 150784
rect 248860 150726 252435 150728
rect 252369 150723 252435 150726
rect 307661 150650 307727 150653
rect 307661 150648 310132 150650
rect 307661 150592 307666 150648
rect 307722 150592 310132 150648
rect 307661 150590 310132 150592
rect 307661 150587 307727 150590
rect 213913 150514 213979 150517
rect 213913 150512 217212 150514
rect 213913 150456 213918 150512
rect 213974 150456 217212 150512
rect 213913 150454 217212 150456
rect 213913 150451 213979 150454
rect 251909 150242 251975 150245
rect 248860 150240 251975 150242
rect 248860 150184 251914 150240
rect 251970 150184 251975 150240
rect 248860 150182 251975 150184
rect 251909 150179 251975 150182
rect 307477 150242 307543 150245
rect 307477 150240 310132 150242
rect 307477 150184 307482 150240
rect 307538 150184 310132 150240
rect 307477 150182 310132 150184
rect 307477 150179 307543 150182
rect 325601 150106 325667 150109
rect 321908 150104 325667 150106
rect 321908 150048 325606 150104
rect 325662 150048 325667 150104
rect 321908 150046 325667 150048
rect 325601 150043 325667 150046
rect 214649 149834 214715 149837
rect 251541 149834 251607 149837
rect 214649 149832 217212 149834
rect 214649 149776 214654 149832
rect 214710 149776 217212 149832
rect 214649 149774 217212 149776
rect 248860 149832 251607 149834
rect 248860 149776 251546 149832
rect 251602 149776 251607 149832
rect 248860 149774 251607 149776
rect 214649 149771 214715 149774
rect 251541 149771 251607 149774
rect 307661 149834 307727 149837
rect 307661 149832 310132 149834
rect 307661 149776 307666 149832
rect 307722 149776 310132 149832
rect 307661 149774 310132 149776
rect 307661 149771 307727 149774
rect 250621 149698 250687 149701
rect 259494 149698 259500 149700
rect 250621 149696 259500 149698
rect 250621 149640 250626 149696
rect 250682 149640 259500 149696
rect 250621 149638 259500 149640
rect 250621 149635 250687 149638
rect 259494 149636 259500 149638
rect 259564 149636 259570 149700
rect 264973 149698 265039 149701
rect 293902 149698 293908 149700
rect 264973 149696 293908 149698
rect 264973 149640 264978 149696
rect 265034 149640 293908 149696
rect 264973 149638 293908 149640
rect 264973 149635 265039 149638
rect 293902 149636 293908 149638
rect 293972 149636 293978 149700
rect 323025 149426 323091 149429
rect 321908 149424 323091 149426
rect 321908 149368 323030 149424
rect 323086 149368 323091 149424
rect 321908 149366 323091 149368
rect 323025 149363 323091 149366
rect 249885 149290 249951 149293
rect 248860 149288 249951 149290
rect 248860 149232 249890 149288
rect 249946 149232 249951 149288
rect 248860 149230 249951 149232
rect 249885 149227 249951 149230
rect 305637 149290 305703 149293
rect 305637 149288 310132 149290
rect 305637 149232 305642 149288
rect 305698 149232 310132 149288
rect 305637 149230 310132 149232
rect 305637 149227 305703 149230
rect 213913 149154 213979 149157
rect 213913 149152 217212 149154
rect 213913 149096 213918 149152
rect 213974 149096 217212 149152
rect 213913 149094 217212 149096
rect 213913 149091 213979 149094
rect 458766 149092 458772 149156
rect 458836 149154 458842 149156
rect 459553 149154 459619 149157
rect 458836 149152 459619 149154
rect 458836 149096 459558 149152
rect 459614 149096 459619 149152
rect 458836 149094 459619 149096
rect 458836 149092 458842 149094
rect 459553 149091 459619 149094
rect 252369 148882 252435 148885
rect 248860 148880 252435 148882
rect 248860 148824 252374 148880
rect 252430 148824 252435 148880
rect 248860 148822 252435 148824
rect 252369 148819 252435 148822
rect 307569 148882 307635 148885
rect 307569 148880 310132 148882
rect 307569 148824 307574 148880
rect 307630 148824 310132 148880
rect 307569 148822 310132 148824
rect 307569 148819 307635 148822
rect 324313 148610 324379 148613
rect 321908 148608 324379 148610
rect 321908 148552 324318 148608
rect 324374 148552 324379 148608
rect 321908 148550 324379 148552
rect 324313 148547 324379 148550
rect 213913 148474 213979 148477
rect 307661 148474 307727 148477
rect 213913 148472 217212 148474
rect 213913 148416 213918 148472
rect 213974 148416 217212 148472
rect 213913 148414 217212 148416
rect 307661 148472 310132 148474
rect 307661 148416 307666 148472
rect 307722 148416 310132 148472
rect 307661 148414 310132 148416
rect 213913 148411 213979 148414
rect 307661 148411 307727 148414
rect 252461 148338 252527 148341
rect 248860 148336 252527 148338
rect 248860 148280 252466 148336
rect 252522 148280 252527 148336
rect 248860 148278 252527 148280
rect 252461 148275 252527 148278
rect 307477 148066 307543 148069
rect 307477 148064 310132 148066
rect 307477 148008 307482 148064
rect 307538 148008 310132 148064
rect 307477 148006 310132 148008
rect 307477 148003 307543 148006
rect 214557 147930 214623 147933
rect 251265 147930 251331 147933
rect 214557 147928 217212 147930
rect 214557 147872 214562 147928
rect 214618 147872 217212 147928
rect 214557 147870 217212 147872
rect 248860 147928 251331 147930
rect 248860 147872 251270 147928
rect 251326 147872 251331 147928
rect 248860 147870 251331 147872
rect 214557 147867 214623 147870
rect 251265 147867 251331 147870
rect 324405 147794 324471 147797
rect 321908 147792 324471 147794
rect 321908 147736 324410 147792
rect 324466 147736 324471 147792
rect 321908 147734 324471 147736
rect 324405 147731 324471 147734
rect 396574 147732 396580 147796
rect 396644 147794 396650 147796
rect 439497 147794 439563 147797
rect 439957 147794 440023 147797
rect 396644 147792 440023 147794
rect 396644 147736 439502 147792
rect 439558 147736 439962 147792
rect 440018 147736 440023 147792
rect 396644 147734 440023 147736
rect 396644 147732 396650 147734
rect 439497 147731 439563 147734
rect 439957 147731 440023 147734
rect 451406 147732 451412 147796
rect 451476 147794 451482 147796
rect 451549 147794 451615 147797
rect 451476 147792 451615 147794
rect 451476 147736 451554 147792
rect 451610 147736 451615 147792
rect 451476 147734 451615 147736
rect 451476 147732 451482 147734
rect 451549 147731 451615 147734
rect 307569 147658 307635 147661
rect 307569 147656 310132 147658
rect 307569 147600 307574 147656
rect 307630 147600 310132 147656
rect 307569 147598 310132 147600
rect 307569 147595 307635 147598
rect 252461 147522 252527 147525
rect 248860 147520 252527 147522
rect 248860 147464 252466 147520
rect 252522 147464 252527 147520
rect 248860 147462 252527 147464
rect 252461 147459 252527 147462
rect 213913 147250 213979 147253
rect 307477 147250 307543 147253
rect 213913 147248 217212 147250
rect 213913 147192 213918 147248
rect 213974 147192 217212 147248
rect 213913 147190 217212 147192
rect 307477 147248 310132 147250
rect 307477 147192 307482 147248
rect 307538 147192 310132 147248
rect 307477 147190 310132 147192
rect 213913 147187 213979 147190
rect 307477 147187 307543 147190
rect 324313 147114 324379 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 324313 147051 324379 147054
rect 251173 146978 251239 146981
rect 248860 146976 251239 146978
rect 248860 146920 251178 146976
rect 251234 146920 251239 146976
rect 248860 146918 251239 146920
rect 251173 146915 251239 146918
rect 422201 146978 422267 146981
rect 450118 146978 450124 146980
rect 422201 146976 450124 146978
rect 422201 146920 422206 146976
rect 422262 146920 450124 146976
rect 422201 146918 450124 146920
rect 422201 146915 422267 146918
rect 450118 146916 450124 146918
rect 450188 146916 450194 146980
rect 307661 146842 307727 146845
rect 307661 146840 310132 146842
rect 307661 146784 307666 146840
rect 307722 146784 310132 146840
rect 307661 146782 310132 146784
rect 307661 146779 307727 146782
rect 214649 146570 214715 146573
rect 252369 146570 252435 146573
rect 214649 146568 217212 146570
rect 214649 146512 214654 146568
rect 214710 146512 217212 146568
rect 214649 146510 217212 146512
rect 248860 146568 252435 146570
rect 248860 146512 252374 146568
rect 252430 146512 252435 146568
rect 248860 146510 252435 146512
rect 214649 146507 214715 146510
rect 252369 146507 252435 146510
rect 308489 146434 308555 146437
rect 308489 146432 310132 146434
rect 308489 146376 308494 146432
rect 308550 146376 310132 146432
rect 308489 146374 310132 146376
rect 308489 146371 308555 146374
rect 324313 146298 324379 146301
rect 321908 146296 324379 146298
rect 321908 146240 324318 146296
rect 324374 146240 324379 146296
rect 321908 146238 324379 146240
rect 324313 146235 324379 146238
rect 251909 146026 251975 146029
rect 248860 146024 251975 146026
rect 248860 145968 251914 146024
rect 251970 145968 251975 146024
rect 248860 145966 251975 145968
rect 251909 145963 251975 145966
rect 214005 145890 214071 145893
rect 307477 145890 307543 145893
rect 214005 145888 217212 145890
rect 214005 145832 214010 145888
rect 214066 145832 217212 145888
rect 214005 145830 217212 145832
rect 307477 145888 310132 145890
rect 307477 145832 307482 145888
rect 307538 145832 310132 145888
rect 307477 145830 310132 145832
rect 214005 145827 214071 145830
rect 307477 145827 307543 145830
rect 252461 145618 252527 145621
rect 248860 145616 252527 145618
rect 248860 145560 252466 145616
rect 252522 145560 252527 145616
rect 248860 145558 252527 145560
rect 252461 145555 252527 145558
rect 397453 145618 397519 145621
rect 449249 145618 449315 145621
rect 397453 145616 400108 145618
rect 397453 145560 397458 145616
rect 397514 145560 400108 145616
rect 397453 145558 400108 145560
rect 449206 145616 449315 145618
rect 449206 145560 449254 145616
rect 449310 145560 449315 145616
rect 397453 145555 397519 145558
rect 449206 145555 449315 145560
rect 307661 145482 307727 145485
rect 324405 145482 324471 145485
rect 307661 145480 310132 145482
rect 307661 145424 307666 145480
rect 307722 145424 310132 145480
rect 307661 145422 310132 145424
rect 321908 145480 324471 145482
rect 321908 145424 324410 145480
rect 324466 145424 324471 145480
rect 321908 145422 324471 145424
rect 307661 145419 307727 145422
rect 324405 145419 324471 145422
rect 213913 145210 213979 145213
rect 213913 145208 217212 145210
rect 213913 145152 213918 145208
rect 213974 145152 217212 145208
rect 213913 145150 217212 145152
rect 213913 145147 213979 145150
rect 252093 145074 252159 145077
rect 248860 145072 252159 145074
rect 248860 145016 252098 145072
rect 252154 145016 252159 145072
rect 248860 145014 252159 145016
rect 252093 145011 252159 145014
rect 306557 145074 306623 145077
rect 306557 145072 310132 145074
rect 306557 145016 306562 145072
rect 306618 145016 310132 145072
rect 449206 145044 449266 145555
rect 306557 145014 310132 145016
rect 306557 145011 306623 145014
rect 324313 144802 324379 144805
rect 321908 144800 324379 144802
rect 321908 144744 324318 144800
rect 324374 144744 324379 144800
rect 321908 144742 324379 144744
rect 324313 144739 324379 144742
rect 251541 144666 251607 144669
rect 248860 144664 251607 144666
rect 248860 144608 251546 144664
rect 251602 144608 251607 144664
rect 248860 144606 251607 144608
rect 251541 144603 251607 144606
rect 307201 144666 307267 144669
rect 307201 144664 310132 144666
rect 307201 144608 307206 144664
rect 307262 144608 310132 144664
rect 307201 144606 310132 144608
rect 307201 144603 307267 144606
rect 213913 144530 213979 144533
rect 213913 144528 217212 144530
rect 213913 144472 213918 144528
rect 213974 144472 217212 144528
rect 213913 144470 217212 144472
rect 213913 144467 213979 144470
rect 452561 144394 452627 144397
rect 449788 144392 452627 144394
rect 449788 144336 452566 144392
rect 452622 144336 452627 144392
rect 449788 144334 452627 144336
rect 452561 144331 452627 144334
rect 307385 144258 307451 144261
rect 397453 144258 397519 144261
rect 307385 144256 310132 144258
rect 307385 144200 307390 144256
rect 307446 144200 310132 144256
rect 307385 144198 310132 144200
rect 397453 144256 400108 144258
rect 397453 144200 397458 144256
rect 397514 144200 400108 144256
rect 397453 144198 400108 144200
rect 307385 144195 307451 144198
rect 397453 144195 397519 144198
rect 252461 144122 252527 144125
rect 248860 144120 252527 144122
rect 248860 144064 252466 144120
rect 252522 144064 252527 144120
rect 248860 144062 252527 144064
rect 252461 144059 252527 144062
rect 252645 144122 252711 144125
rect 292614 144122 292620 144124
rect 252645 144120 292620 144122
rect 252645 144064 252650 144120
rect 252706 144064 292620 144120
rect 252645 144062 292620 144064
rect 252645 144059 252711 144062
rect 292614 144060 292620 144062
rect 292684 144060 292690 144124
rect 324405 143986 324471 143989
rect 321908 143984 324471 143986
rect 321908 143928 324410 143984
rect 324466 143928 324471 143984
rect 321908 143926 324471 143928
rect 324405 143923 324471 143926
rect 307477 143850 307543 143853
rect 200070 143790 217212 143850
rect 307477 143848 310132 143850
rect 307477 143792 307482 143848
rect 307538 143792 310132 143848
rect 307477 143790 310132 143792
rect 166206 143652 166212 143716
rect 166276 143714 166282 143716
rect 200070 143714 200130 143790
rect 307477 143787 307543 143790
rect 252185 143714 252251 143717
rect 166276 143654 200130 143714
rect 248860 143712 252251 143714
rect 248860 143656 252190 143712
rect 252246 143656 252251 143712
rect 248860 143654 252251 143656
rect 166276 143652 166282 143654
rect 252185 143651 252251 143654
rect 397545 143714 397611 143717
rect 397545 143712 400108 143714
rect 397545 143656 397550 143712
rect 397606 143656 400108 143712
rect 397545 143654 400108 143656
rect 397545 143651 397611 143654
rect 307293 143442 307359 143445
rect 449341 143444 449407 143445
rect 307293 143440 310132 143442
rect 307293 143384 307298 143440
rect 307354 143384 310132 143440
rect 307293 143382 310132 143384
rect 449341 143440 449388 143444
rect 449452 143442 449458 143444
rect 449341 143384 449346 143440
rect 307293 143379 307359 143382
rect 449341 143380 449388 143384
rect 449452 143382 449498 143442
rect 449452 143380 449458 143382
rect 449341 143379 449407 143380
rect 213913 143306 213979 143309
rect 449525 143306 449591 143309
rect 213913 143304 217212 143306
rect 213913 143248 213918 143304
rect 213974 143248 217212 143304
rect 213913 143246 217212 143248
rect 449525 143304 449634 143306
rect 449525 143248 449530 143304
rect 449586 143248 449634 143304
rect 213913 143243 213979 143246
rect 449525 143243 449634 143248
rect 251725 143170 251791 143173
rect 324313 143170 324379 143173
rect 248860 143168 251791 143170
rect 248860 143112 251730 143168
rect 251786 143112 251791 143168
rect 248860 143110 251791 143112
rect 321908 143168 324379 143170
rect 321908 143112 324318 143168
rect 324374 143112 324379 143168
rect 321908 143110 324379 143112
rect 251725 143107 251791 143110
rect 324313 143107 324379 143110
rect 307661 143034 307727 143037
rect 449574 143034 449634 143243
rect 307661 143032 310132 143034
rect 307661 142976 307666 143032
rect 307722 142976 310132 143032
rect 449574 143004 449788 143034
rect 307661 142974 310132 142976
rect 449604 142974 449818 143004
rect 307661 142971 307727 142974
rect 321553 142898 321619 142901
rect 321510 142896 321619 142898
rect 321510 142840 321558 142896
rect 321614 142840 321619 142896
rect 449758 142898 449818 142974
rect 452469 142898 452535 142901
rect 449758 142896 452535 142898
rect 449758 142868 452474 142896
rect 321510 142835 321619 142840
rect 449788 142840 452474 142868
rect 452530 142840 452535 142896
rect 449788 142838 452535 142840
rect 452469 142835 452535 142838
rect 252461 142762 252527 142765
rect 248860 142760 252527 142762
rect 248860 142704 252466 142760
rect 252522 142704 252527 142760
rect 248860 142702 252527 142704
rect 252461 142699 252527 142702
rect 213913 142626 213979 142629
rect 251081 142626 251147 142629
rect 265014 142626 265020 142628
rect 213913 142624 217212 142626
rect 213913 142568 213918 142624
rect 213974 142568 217212 142624
rect 213913 142566 217212 142568
rect 251081 142624 265020 142626
rect 251081 142568 251086 142624
rect 251142 142568 265020 142624
rect 251081 142566 265020 142568
rect 213913 142563 213979 142566
rect 251081 142563 251147 142566
rect 265014 142564 265020 142566
rect 265084 142564 265090 142628
rect 307477 142490 307543 142493
rect 307477 142488 310132 142490
rect 307477 142432 307482 142488
rect 307538 142432 310132 142488
rect 321510 142460 321570 142835
rect 307477 142430 310132 142432
rect 307477 142427 307543 142430
rect 451457 142354 451523 142357
rect 449788 142352 451523 142354
rect 449788 142296 451462 142352
rect 451518 142296 451523 142352
rect 449788 142294 451523 142296
rect 451457 142291 451523 142294
rect 263542 142218 263548 142220
rect 248860 142158 263548 142218
rect 263542 142156 263548 142158
rect 263612 142156 263618 142220
rect 397545 142218 397611 142221
rect 397545 142216 400108 142218
rect 397545 142160 397550 142216
rect 397606 142160 400108 142216
rect 397545 142158 400108 142160
rect 397545 142155 397611 142158
rect 307661 142082 307727 142085
rect 307661 142080 310132 142082
rect 307661 142024 307666 142080
rect 307722 142024 310132 142080
rect 307661 142022 310132 142024
rect 307661 142019 307727 142022
rect 214005 141946 214071 141949
rect 214005 141944 217212 141946
rect 214005 141888 214010 141944
rect 214066 141888 217212 141944
rect 214005 141886 217212 141888
rect 214005 141883 214071 141886
rect 262254 141810 262260 141812
rect 248860 141750 262260 141810
rect 262254 141748 262260 141750
rect 262324 141748 262330 141812
rect 307334 141612 307340 141676
rect 307404 141674 307410 141676
rect 324313 141674 324379 141677
rect 307404 141614 310132 141674
rect 321908 141672 324379 141674
rect 321908 141616 324318 141672
rect 324374 141616 324379 141672
rect 321908 141614 324379 141616
rect 307404 141612 307410 141614
rect 324313 141611 324379 141614
rect 397453 141674 397519 141677
rect 397453 141672 400108 141674
rect 397453 141616 397458 141672
rect 397514 141616 400108 141672
rect 397453 141614 400108 141616
rect 397453 141611 397519 141614
rect 449433 141538 449499 141541
rect 449390 141536 449499 141538
rect 449390 141480 449438 141536
rect 449494 141480 449499 141536
rect 449390 141475 449499 141480
rect 251725 141402 251791 141405
rect 248860 141400 251791 141402
rect 248860 141344 251730 141400
rect 251786 141344 251791 141400
rect 248860 141342 251791 141344
rect 251725 141339 251791 141342
rect 213913 141266 213979 141269
rect 307569 141266 307635 141269
rect 213913 141264 217212 141266
rect 213913 141208 213918 141264
rect 213974 141208 217212 141264
rect 213913 141206 217212 141208
rect 307569 141264 310132 141266
rect 307569 141208 307574 141264
rect 307630 141208 310132 141264
rect 307569 141206 310132 141208
rect 213913 141203 213979 141206
rect 307569 141203 307635 141206
rect 449390 140964 449450 141475
rect 251214 140858 251220 140860
rect 248860 140798 251220 140858
rect 251214 140796 251220 140798
rect 251284 140796 251290 140860
rect 307661 140858 307727 140861
rect 324405 140858 324471 140861
rect 307661 140856 310132 140858
rect 307661 140800 307666 140856
rect 307722 140800 310132 140856
rect 307661 140798 310132 140800
rect 321908 140856 324471 140858
rect 321908 140800 324410 140856
rect 324466 140800 324471 140856
rect 321908 140798 324471 140800
rect 307661 140795 307727 140798
rect 324405 140795 324471 140798
rect 213177 140586 213243 140589
rect 213177 140584 217212 140586
rect 213177 140528 213182 140584
rect 213238 140528 217212 140584
rect 213177 140526 217212 140528
rect 213177 140523 213243 140526
rect 255262 140450 255268 140452
rect 248860 140390 255268 140450
rect 255262 140388 255268 140390
rect 255332 140388 255338 140452
rect 307569 140450 307635 140453
rect 307569 140448 310132 140450
rect 307569 140392 307574 140448
rect 307630 140392 310132 140448
rect 307569 140390 310132 140392
rect 307569 140387 307635 140390
rect 397361 140314 397427 140317
rect 451917 140314 451983 140317
rect 397361 140312 400108 140314
rect 397361 140256 397366 140312
rect 397422 140256 400108 140312
rect 397361 140254 400108 140256
rect 449788 140312 451983 140314
rect 449788 140256 451922 140312
rect 451978 140256 451983 140312
rect 449788 140254 451983 140256
rect 397361 140251 397427 140254
rect 451917 140251 451983 140254
rect 324313 140178 324379 140181
rect 321908 140176 324379 140178
rect 321908 140120 324318 140176
rect 324374 140120 324379 140176
rect 321908 140118 324379 140120
rect 324313 140115 324379 140118
rect 306557 140042 306623 140045
rect 400121 140042 400187 140045
rect 306557 140040 310132 140042
rect 306557 139984 306562 140040
rect 306618 139984 310132 140040
rect 306557 139982 310132 139984
rect 400078 140040 400187 140042
rect 400078 139984 400126 140040
rect 400182 139984 400187 140040
rect 306557 139979 306623 139982
rect 400078 139979 400187 139984
rect 213913 139906 213979 139909
rect 256918 139906 256924 139908
rect 213913 139904 217212 139906
rect 213913 139848 213918 139904
rect 213974 139848 217212 139904
rect 213913 139846 217212 139848
rect 248860 139846 256924 139906
rect 213913 139843 213979 139846
rect 256918 139844 256924 139846
rect 256988 139844 256994 139908
rect 307661 139634 307727 139637
rect 307661 139632 310132 139634
rect 307661 139576 307666 139632
rect 307722 139576 310132 139632
rect 400078 139604 400138 139979
rect 307661 139574 310132 139576
rect 307661 139571 307727 139574
rect 251725 139498 251791 139501
rect 248860 139496 251791 139498
rect 248860 139440 251730 139496
rect 251786 139440 251791 139496
rect 248860 139438 251791 139440
rect 251725 139435 251791 139438
rect 580349 139362 580415 139365
rect 583520 139362 584960 139452
rect 580349 139360 584960 139362
rect 217182 138818 217242 139196
rect 307477 139090 307543 139093
rect 307477 139088 310132 139090
rect 307477 139032 307482 139088
rect 307538 139032 310132 139088
rect 307477 139030 310132 139032
rect 307477 139027 307543 139030
rect 252461 138954 252527 138957
rect 248860 138952 252527 138954
rect 248860 138896 252466 138952
rect 252522 138896 252527 138952
rect 248860 138894 252527 138896
rect 252461 138891 252527 138894
rect 200070 138758 217242 138818
rect 167678 138076 167684 138140
rect 167748 138138 167754 138140
rect 200070 138138 200130 138758
rect 213913 138682 213979 138685
rect 307661 138682 307727 138685
rect 321878 138682 321938 139332
rect 580349 139304 580354 139360
rect 580410 139304 584960 139360
rect 580349 139302 584960 139304
rect 580349 139299 580415 139302
rect 583520 139212 584960 139302
rect 397453 138954 397519 138957
rect 451273 138954 451339 138957
rect 397453 138952 400108 138954
rect 397453 138896 397458 138952
rect 397514 138896 400108 138952
rect 397453 138894 400108 138896
rect 449788 138952 451339 138954
rect 449788 138896 451278 138952
rect 451334 138896 451339 138952
rect 449788 138894 451339 138896
rect 397453 138891 397519 138894
rect 451273 138891 451339 138894
rect 328494 138682 328500 138684
rect 213913 138680 217212 138682
rect 213913 138624 213918 138680
rect 213974 138624 217212 138680
rect 213913 138622 217212 138624
rect 307661 138680 310132 138682
rect 307661 138624 307666 138680
rect 307722 138624 310132 138680
rect 307661 138622 310132 138624
rect 321878 138622 328500 138682
rect 213913 138619 213979 138622
rect 307661 138619 307727 138622
rect 328494 138620 328500 138622
rect 328564 138620 328570 138684
rect 251725 138546 251791 138549
rect 324313 138546 324379 138549
rect 248860 138544 251791 138546
rect 248860 138488 251730 138544
rect 251786 138488 251791 138544
rect 248860 138486 251791 138488
rect 321908 138544 324379 138546
rect 321908 138488 324318 138544
rect 324374 138488 324379 138544
rect 321908 138486 324379 138488
rect 251725 138483 251791 138486
rect 324313 138483 324379 138486
rect 307569 138274 307635 138277
rect 452101 138274 452167 138277
rect 307569 138272 310132 138274
rect 307569 138216 307574 138272
rect 307630 138216 310132 138272
rect 307569 138214 310132 138216
rect 449788 138272 452167 138274
rect 449788 138216 452106 138272
rect 452162 138216 452167 138272
rect 449788 138214 452167 138216
rect 307569 138211 307635 138214
rect 452101 138211 452167 138214
rect 167748 138078 200130 138138
rect 167748 138076 167754 138078
rect 214097 138002 214163 138005
rect 251357 138002 251423 138005
rect 449985 138002 450051 138005
rect 214097 138000 217212 138002
rect 214097 137944 214102 138000
rect 214158 137944 217212 138000
rect 214097 137942 217212 137944
rect 248860 138000 251423 138002
rect 248860 137944 251362 138000
rect 251418 137944 251423 138000
rect 248860 137942 251423 137944
rect 214097 137939 214163 137942
rect 251357 137939 251423 137942
rect 449758 138000 450051 138002
rect 449758 137944 449990 138000
rect 450046 137944 450051 138000
rect 449758 137942 450051 137944
rect 306741 137866 306807 137869
rect 324313 137866 324379 137869
rect 306741 137864 310132 137866
rect 306741 137808 306746 137864
rect 306802 137808 310132 137864
rect 306741 137806 310132 137808
rect 321908 137864 324379 137866
rect 321908 137808 324318 137864
rect 324374 137808 324379 137864
rect 321908 137806 324379 137808
rect 306741 137803 306807 137806
rect 324313 137803 324379 137806
rect 252461 137594 252527 137597
rect 248860 137592 252527 137594
rect 248860 137536 252466 137592
rect 252522 137536 252527 137592
rect 248860 137534 252527 137536
rect 252461 137531 252527 137534
rect 397453 137594 397519 137597
rect 397453 137592 400108 137594
rect 397453 137536 397458 137592
rect 397514 137536 400108 137592
rect 449758 137564 449818 137942
rect 449985 137939 450051 137942
rect 397453 137534 400108 137536
rect 397453 137531 397519 137534
rect 307661 137458 307727 137461
rect 307661 137456 310132 137458
rect 307661 137400 307666 137456
rect 307722 137400 310132 137456
rect 307661 137398 310132 137400
rect 307661 137395 307727 137398
rect 213913 137322 213979 137325
rect 213913 137320 217212 137322
rect 213913 137264 213918 137320
rect 213974 137264 217212 137320
rect 213913 137262 217212 137264
rect 213913 137259 213979 137262
rect 250621 137050 250687 137053
rect 248860 137048 250687 137050
rect 248860 136992 250626 137048
rect 250682 136992 250687 137048
rect 248860 136990 250687 136992
rect 250621 136987 250687 136990
rect 307150 136988 307156 137052
rect 307220 137050 307226 137052
rect 323301 137050 323367 137053
rect 307220 136990 310132 137050
rect 321908 137048 323367 137050
rect 321908 136992 323306 137048
rect 323362 136992 323367 137048
rect 321908 136990 323367 136992
rect 307220 136988 307226 136990
rect 323301 136987 323367 136990
rect 397545 136914 397611 136917
rect 397545 136912 400108 136914
rect 397545 136856 397550 136912
rect 397606 136856 400108 136912
rect 397545 136854 400108 136856
rect 397545 136851 397611 136854
rect 214005 136642 214071 136645
rect 254526 136642 254532 136644
rect 214005 136640 217212 136642
rect 214005 136584 214010 136640
rect 214066 136584 217212 136640
rect 214005 136582 217212 136584
rect 248860 136582 254532 136642
rect 214005 136579 214071 136582
rect 254526 136580 254532 136582
rect 254596 136580 254602 136644
rect 306741 136642 306807 136645
rect 306741 136640 310132 136642
rect 306741 136584 306746 136640
rect 306802 136584 310132 136640
rect 306741 136582 310132 136584
rect 306741 136579 306807 136582
rect 341374 136580 341380 136644
rect 341444 136642 341450 136644
rect 390185 136642 390251 136645
rect 450537 136642 450603 136645
rect 341444 136640 390251 136642
rect 341444 136584 390190 136640
rect 390246 136584 390251 136640
rect 341444 136582 390251 136584
rect 341444 136580 341450 136582
rect 390185 136579 390251 136582
rect 449758 136640 450603 136642
rect 449758 136584 450542 136640
rect 450598 136584 450603 136640
rect 449758 136582 450603 136584
rect 323393 136370 323459 136373
rect 321908 136368 323459 136370
rect 321908 136312 323398 136368
rect 323454 136312 323459 136368
rect 321908 136310 323459 136312
rect 323393 136307 323459 136310
rect 252461 136234 252527 136237
rect 248860 136232 252527 136234
rect 248860 136176 252466 136232
rect 252522 136176 252527 136232
rect 248860 136174 252527 136176
rect 252461 136171 252527 136174
rect 306557 136234 306623 136237
rect 306557 136232 310132 136234
rect 306557 136176 306562 136232
rect 306618 136176 310132 136232
rect 449758 136204 449818 136582
rect 450537 136579 450603 136582
rect 306557 136174 310132 136176
rect 306557 136171 306623 136174
rect 214097 135962 214163 135965
rect 214097 135960 217212 135962
rect 214097 135904 214102 135960
rect 214158 135904 217212 135960
rect 214097 135902 217212 135904
rect 214097 135899 214163 135902
rect 251725 135690 251791 135693
rect 248860 135688 251791 135690
rect 248860 135632 251730 135688
rect 251786 135632 251791 135688
rect 248860 135630 251791 135632
rect 251725 135627 251791 135630
rect 306925 135690 306991 135693
rect 306925 135688 310132 135690
rect 306925 135632 306930 135688
rect 306986 135632 310132 135688
rect 306925 135630 310132 135632
rect 306925 135627 306991 135630
rect 324313 135554 324379 135557
rect 450077 135554 450143 135557
rect 321908 135552 324379 135554
rect 321908 135496 324318 135552
rect 324374 135496 324379 135552
rect 321908 135494 324379 135496
rect 449788 135552 450143 135554
rect 449788 135496 450082 135552
rect 450138 135496 450143 135552
rect 449788 135494 450143 135496
rect 324313 135491 324379 135494
rect 450077 135491 450143 135494
rect 397453 135418 397519 135421
rect 397453 135416 400108 135418
rect 397453 135360 397458 135416
rect 397514 135360 400108 135416
rect 397453 135358 400108 135360
rect 397453 135355 397519 135358
rect 213913 135282 213979 135285
rect 252369 135282 252435 135285
rect 213913 135280 217212 135282
rect 213913 135224 213918 135280
rect 213974 135224 217212 135280
rect 213913 135222 217212 135224
rect 248860 135280 252435 135282
rect 248860 135224 252374 135280
rect 252430 135224 252435 135280
rect 248860 135222 252435 135224
rect 213913 135219 213979 135222
rect 252369 135219 252435 135222
rect 307661 135282 307727 135285
rect 307661 135280 310132 135282
rect 307661 135224 307666 135280
rect 307722 135224 310132 135280
rect 307661 135222 310132 135224
rect 307661 135219 307727 135222
rect 307477 134874 307543 134877
rect 307477 134872 310132 134874
rect 307477 134816 307482 134872
rect 307538 134816 310132 134872
rect 307477 134814 310132 134816
rect 307477 134811 307543 134814
rect 251449 134738 251515 134741
rect 324313 134738 324379 134741
rect 248860 134736 251515 134738
rect 248860 134680 251454 134736
rect 251510 134680 251515 134736
rect 248860 134678 251515 134680
rect 321908 134736 324379 134738
rect 321908 134680 324318 134736
rect 324374 134680 324379 134736
rect 321908 134678 324379 134680
rect 251449 134675 251515 134678
rect 324313 134675 324379 134678
rect 397453 134738 397519 134741
rect 397453 134736 400108 134738
rect 397453 134680 397458 134736
rect 397514 134680 400108 134736
rect 397453 134678 400108 134680
rect 397453 134675 397519 134678
rect 214005 134602 214071 134605
rect 214005 134600 217212 134602
rect 214005 134544 214010 134600
rect 214066 134544 217212 134600
rect 214005 134542 217212 134544
rect 214005 134539 214071 134542
rect 270033 134466 270099 134469
rect 307334 134466 307340 134468
rect 270033 134464 307340 134466
rect 270033 134408 270038 134464
rect 270094 134408 307340 134464
rect 270033 134406 307340 134408
rect 270033 134403 270099 134406
rect 307334 134404 307340 134406
rect 307404 134404 307410 134468
rect 307569 134466 307635 134469
rect 307569 134464 310132 134466
rect 307569 134408 307574 134464
rect 307630 134408 310132 134464
rect 307569 134406 310132 134408
rect 307569 134403 307635 134406
rect 252461 134330 252527 134333
rect 248860 134328 252527 134330
rect 248860 134272 252466 134328
rect 252522 134272 252527 134328
rect 248860 134270 252527 134272
rect 252461 134267 252527 134270
rect 451917 134194 451983 134197
rect 449788 134192 451983 134194
rect 449788 134136 451922 134192
rect 451978 134136 451983 134192
rect 449788 134134 451983 134136
rect 451917 134131 451983 134134
rect 307661 134058 307727 134061
rect 324405 134058 324471 134061
rect 307661 134056 310132 134058
rect 307661 134000 307666 134056
rect 307722 134000 310132 134056
rect 307661 133998 310132 134000
rect 321908 134056 324471 134058
rect 321908 134000 324410 134056
rect 324466 134000 324471 134056
rect 321908 133998 324471 134000
rect 307661 133995 307727 133998
rect 324405 133995 324471 133998
rect 213913 133922 213979 133925
rect 213913 133920 217212 133922
rect 213913 133864 213918 133920
rect 213974 133864 217212 133920
rect 213913 133862 217212 133864
rect 213913 133859 213979 133862
rect 251357 133786 251423 133789
rect 248860 133784 251423 133786
rect 248860 133728 251362 133784
rect 251418 133728 251423 133784
rect 248860 133726 251423 133728
rect 251357 133723 251423 133726
rect 307477 133650 307543 133653
rect 307477 133648 310132 133650
rect 307477 133592 307482 133648
rect 307538 133592 310132 133648
rect 307477 133590 310132 133592
rect 307477 133587 307543 133590
rect 451038 133514 451044 133516
rect 449788 133454 451044 133514
rect 451038 133452 451044 133454
rect 451108 133514 451114 133516
rect 452193 133514 452259 133517
rect 451108 133512 452259 133514
rect 451108 133456 452198 133512
rect 452254 133456 452259 133512
rect 451108 133454 452259 133456
rect 451108 133452 451114 133454
rect 452193 133451 452259 133454
rect 214005 133378 214071 133381
rect 252369 133378 252435 133381
rect 214005 133376 217212 133378
rect 214005 133320 214010 133376
rect 214066 133320 217212 133376
rect 214005 133318 217212 133320
rect 248860 133376 252435 133378
rect 248860 133320 252374 133376
rect 252430 133320 252435 133376
rect 248860 133318 252435 133320
rect 214005 133315 214071 133318
rect 252369 133315 252435 133318
rect 397453 133378 397519 133381
rect 397453 133376 400108 133378
rect 397453 133320 397458 133376
rect 397514 133320 400108 133376
rect 397453 133318 400108 133320
rect 397453 133315 397519 133318
rect 307569 133242 307635 133245
rect 324313 133242 324379 133245
rect 307569 133240 310132 133242
rect 307569 133184 307574 133240
rect 307630 133184 310132 133240
rect 307569 133182 310132 133184
rect 321908 133240 324379 133242
rect 321908 133184 324318 133240
rect 324374 133184 324379 133240
rect 321908 133182 324379 133184
rect 307569 133179 307635 133182
rect 324313 133179 324379 133182
rect 252461 132834 252527 132837
rect 248860 132832 252527 132834
rect 248860 132776 252466 132832
rect 252522 132776 252527 132832
rect 248860 132774 252527 132776
rect 252461 132771 252527 132774
rect 213913 132698 213979 132701
rect 307661 132698 307727 132701
rect 397545 132698 397611 132701
rect 213913 132696 217212 132698
rect 213913 132640 213918 132696
rect 213974 132640 217212 132696
rect 213913 132638 217212 132640
rect 307661 132696 310132 132698
rect 307661 132640 307666 132696
rect 307722 132640 310132 132696
rect 307661 132638 310132 132640
rect 397545 132696 400108 132698
rect 397545 132640 397550 132696
rect 397606 132640 400108 132696
rect 397545 132638 400108 132640
rect 213913 132635 213979 132638
rect 307661 132635 307727 132638
rect 397545 132635 397611 132638
rect 252461 132426 252527 132429
rect 248860 132424 252527 132426
rect 248860 132368 252466 132424
rect 252522 132368 252527 132424
rect 248860 132366 252527 132368
rect 252461 132363 252527 132366
rect 307477 132290 307543 132293
rect 307477 132288 310132 132290
rect 307477 132232 307482 132288
rect 307538 132232 310132 132288
rect 307477 132230 310132 132232
rect 307477 132227 307543 132230
rect 166390 131412 166396 131476
rect 166460 131474 166466 131476
rect 217182 131474 217242 131988
rect 251541 131882 251607 131885
rect 248860 131880 251607 131882
rect 248860 131824 251546 131880
rect 251602 131824 251607 131880
rect 248860 131822 251607 131824
rect 251541 131819 251607 131822
rect 307569 131882 307635 131885
rect 321878 131882 321938 132396
rect 398741 132154 398807 132157
rect 451406 132154 451412 132156
rect 398741 132152 400108 132154
rect 398741 132096 398746 132152
rect 398802 132096 400108 132152
rect 398741 132094 400108 132096
rect 449788 132094 451412 132154
rect 398741 132091 398807 132094
rect 451406 132092 451412 132094
rect 451476 132092 451482 132156
rect 323485 131882 323551 131885
rect 307569 131880 310132 131882
rect 307569 131824 307574 131880
rect 307630 131824 310132 131880
rect 307569 131822 310132 131824
rect 321878 131880 323551 131882
rect 321878 131824 323490 131880
rect 323546 131824 323551 131880
rect 321878 131822 323551 131824
rect 307569 131819 307635 131822
rect 323485 131819 323551 131822
rect 252093 131474 252159 131477
rect 166460 131414 217242 131474
rect 248860 131472 252159 131474
rect 248860 131416 252098 131472
rect 252154 131416 252159 131472
rect 248860 131414 252159 131416
rect 166460 131412 166466 131414
rect 252093 131411 252159 131414
rect 307661 131474 307727 131477
rect 307661 131472 310132 131474
rect 307661 131416 307666 131472
rect 307722 131416 310132 131472
rect 307661 131414 310132 131416
rect 307661 131411 307727 131414
rect 213269 131338 213335 131341
rect 321878 131338 321938 131716
rect 331438 131338 331444 131340
rect 213269 131336 217212 131338
rect 213269 131280 213274 131336
rect 213330 131280 217212 131336
rect 213269 131278 217212 131280
rect 321878 131278 331444 131338
rect 213269 131275 213335 131278
rect 331438 131276 331444 131278
rect 331508 131276 331514 131340
rect 323485 131202 323551 131205
rect 342294 131202 342300 131204
rect 323485 131200 342300 131202
rect 323485 131144 323490 131200
rect 323546 131144 342300 131200
rect 323485 131142 342300 131144
rect 323485 131139 323551 131142
rect 342294 131140 342300 131142
rect 342364 131140 342370 131204
rect 449758 131202 449818 131308
rect 449985 131202 450051 131205
rect 449758 131200 450051 131202
rect 449758 131144 449990 131200
rect 450046 131144 450051 131200
rect 449758 131142 450051 131144
rect 449985 131139 450051 131142
rect 307109 131066 307175 131069
rect 307109 131064 310132 131066
rect 307109 131008 307114 131064
rect 307170 131008 310132 131064
rect 307109 131006 310132 131008
rect 307109 131003 307175 131006
rect 252461 130930 252527 130933
rect 324313 130930 324379 130933
rect 248860 130928 252527 130930
rect 248860 130872 252466 130928
rect 252522 130872 252527 130928
rect 248860 130870 252527 130872
rect 321908 130928 324379 130930
rect 321908 130872 324318 130928
rect 324374 130872 324379 130928
rect 321908 130870 324379 130872
rect 252461 130867 252527 130870
rect 324313 130867 324379 130870
rect 452561 130794 452627 130797
rect 449788 130792 452627 130794
rect 449788 130764 452566 130792
rect 449758 130736 452566 130764
rect 452622 130736 452627 130792
rect 449758 130734 452627 130736
rect 213913 130658 213979 130661
rect 307569 130658 307635 130661
rect 397545 130658 397611 130661
rect 213913 130656 217212 130658
rect 213913 130600 213918 130656
rect 213974 130600 217212 130656
rect 213913 130598 217212 130600
rect 307569 130656 310132 130658
rect 307569 130600 307574 130656
rect 307630 130600 310132 130656
rect 307569 130598 310132 130600
rect 397545 130656 400108 130658
rect 397545 130600 397550 130656
rect 397606 130600 400108 130656
rect 397545 130598 400108 130600
rect 213913 130595 213979 130598
rect 307569 130595 307635 130598
rect 397545 130595 397611 130598
rect 252461 130522 252527 130525
rect 248860 130520 252527 130522
rect 248860 130464 252466 130520
rect 252522 130464 252527 130520
rect 248860 130462 252527 130464
rect 252461 130459 252527 130462
rect 449390 130522 449450 130628
rect 449758 130522 449818 130734
rect 452561 130731 452627 130734
rect 449390 130462 449818 130522
rect 307477 130250 307543 130253
rect 307477 130248 310132 130250
rect 307477 130192 307482 130248
rect 307538 130192 310132 130248
rect 307477 130190 310132 130192
rect 307477 130187 307543 130190
rect 449390 130117 449450 130462
rect 252369 130114 252435 130117
rect 324405 130114 324471 130117
rect 248860 130112 252435 130114
rect 248860 130056 252374 130112
rect 252430 130056 252435 130112
rect 248860 130054 252435 130056
rect 321908 130112 324471 130114
rect 321908 130056 324410 130112
rect 324466 130056 324471 130112
rect 321908 130054 324471 130056
rect 449390 130112 449499 130117
rect 449390 130056 449438 130112
rect 449494 130056 449499 130112
rect 449390 130054 449499 130056
rect 252369 130051 252435 130054
rect 324405 130051 324471 130054
rect 449433 130051 449499 130054
rect 397453 129978 397519 129981
rect 398189 129978 398255 129981
rect 200070 129918 217212 129978
rect 397453 129976 400108 129978
rect 397453 129920 397458 129976
rect 397514 129920 398194 129976
rect 398250 129920 400108 129976
rect 397453 129918 400108 129920
rect 167494 129780 167500 129844
rect 167564 129842 167570 129844
rect 200070 129842 200130 129918
rect 397453 129915 397519 129918
rect 398189 129915 398255 129918
rect 167564 129782 200130 129842
rect 307661 129842 307727 129845
rect 307661 129840 310132 129842
rect 307661 129784 307666 129840
rect 307722 129784 310132 129840
rect 307661 129782 310132 129784
rect 167564 129780 167570 129782
rect 307661 129779 307727 129782
rect 252461 129570 252527 129573
rect 248860 129568 252527 129570
rect 248860 129512 252466 129568
rect 252522 129512 252527 129568
rect 248860 129510 252527 129512
rect 252461 129507 252527 129510
rect 324313 129434 324379 129437
rect 452561 129434 452627 129437
rect 321908 129432 324379 129434
rect 321908 129376 324318 129432
rect 324374 129376 324379 129432
rect 321908 129374 324379 129376
rect 449788 129432 452627 129434
rect 449788 129376 452566 129432
rect 452622 129376 452627 129432
rect 449788 129374 452627 129376
rect 324313 129371 324379 129374
rect 452561 129371 452627 129374
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 306557 129298 306623 129301
rect 306557 129296 310132 129298
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 66161 129235 66227 129238
rect 217182 128890 217242 129268
rect 306557 129240 306562 129296
rect 306618 129240 310132 129296
rect 306557 129238 310132 129240
rect 306557 129235 306623 129238
rect 251449 129162 251515 129165
rect 449893 129162 449959 129165
rect 248860 129160 251515 129162
rect 248860 129104 251454 129160
rect 251510 129104 251515 129160
rect 248860 129102 251515 129104
rect 251449 129099 251515 129102
rect 449758 129160 449959 129162
rect 449758 129104 449898 129160
rect 449954 129104 449959 129160
rect 449758 129102 449959 129104
rect 200070 128830 217242 128890
rect 307109 128890 307175 128893
rect 307109 128888 310132 128890
rect 307109 128832 307114 128888
rect 307170 128832 310132 128888
rect 307109 128830 310132 128832
rect 169150 128420 169156 128484
rect 169220 128482 169226 128484
rect 200070 128482 200130 128830
rect 307109 128827 307175 128830
rect 213913 128754 213979 128757
rect 397453 128754 397519 128757
rect 213913 128752 217212 128754
rect 213913 128696 213918 128752
rect 213974 128696 217212 128752
rect 213913 128694 217212 128696
rect 397453 128752 400108 128754
rect 397453 128696 397458 128752
rect 397514 128696 400108 128752
rect 449758 128724 449818 129102
rect 449893 129099 449959 129102
rect 397453 128694 400108 128696
rect 213913 128691 213979 128694
rect 397453 128691 397519 128694
rect 252369 128618 252435 128621
rect 324405 128618 324471 128621
rect 248860 128616 252435 128618
rect 248860 128560 252374 128616
rect 252430 128560 252435 128616
rect 248860 128558 252435 128560
rect 321908 128616 324471 128618
rect 321908 128560 324410 128616
rect 324466 128560 324471 128616
rect 321908 128558 324471 128560
rect 252369 128555 252435 128558
rect 324405 128555 324471 128558
rect 169220 128422 200130 128482
rect 169220 128420 169226 128422
rect 301630 128420 301636 128484
rect 301700 128482 301706 128484
rect 301700 128422 310132 128482
rect 301700 128420 301706 128422
rect 252461 128210 252527 128213
rect 248860 128208 252527 128210
rect 248860 128152 252466 128208
rect 252522 128152 252527 128208
rect 248860 128150 252527 128152
rect 252461 128147 252527 128150
rect 65517 128074 65583 128077
rect 68142 128074 68816 128080
rect 65517 128072 68816 128074
rect 65517 128016 65522 128072
rect 65578 128020 68816 128072
rect 65578 128016 68202 128020
rect 65517 128014 68202 128016
rect 65517 128011 65583 128014
rect 214833 128074 214899 128077
rect 307661 128074 307727 128077
rect 214833 128072 217212 128074
rect 214833 128016 214838 128072
rect 214894 128016 217212 128072
rect 214833 128014 217212 128016
rect 307661 128072 310132 128074
rect 307661 128016 307666 128072
rect 307722 128016 310132 128072
rect 307661 128014 310132 128016
rect 214833 128011 214899 128014
rect 307661 128011 307727 128014
rect 397453 127938 397519 127941
rect 398649 127938 398715 127941
rect 397453 127936 400108 127938
rect 397453 127880 397458 127936
rect 397514 127880 398654 127936
rect 398710 127880 400108 127936
rect 397453 127878 400108 127880
rect 397453 127875 397519 127878
rect 398649 127875 398715 127878
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 251633 127666 251699 127669
rect 248860 127664 251699 127666
rect 248860 127608 251638 127664
rect 251694 127608 251699 127664
rect 248860 127606 251699 127608
rect 251633 127603 251699 127606
rect 307109 127666 307175 127669
rect 307109 127664 310132 127666
rect 307109 127608 307114 127664
rect 307170 127608 310132 127664
rect 307109 127606 310132 127608
rect 307109 127603 307175 127606
rect 213913 127394 213979 127397
rect 452101 127394 452167 127397
rect 213913 127392 217212 127394
rect 213913 127336 213918 127392
rect 213974 127336 217212 127392
rect 213913 127334 217212 127336
rect 449788 127392 452167 127394
rect 449788 127336 452106 127392
rect 452162 127336 452167 127392
rect 449788 127334 452167 127336
rect 213913 127331 213979 127334
rect 452101 127331 452167 127334
rect 251909 127258 251975 127261
rect 248860 127256 251975 127258
rect 248860 127200 251914 127256
rect 251970 127200 251975 127256
rect 248860 127198 251975 127200
rect 251909 127195 251975 127198
rect 306741 127258 306807 127261
rect 306741 127256 310132 127258
rect 306741 127200 306746 127256
rect 306802 127200 310132 127256
rect 306741 127198 310132 127200
rect 306741 127195 306807 127198
rect 324405 127122 324471 127125
rect 321908 127120 324471 127122
rect 321908 127064 324410 127120
rect 324466 127064 324471 127120
rect 321908 127062 324471 127064
rect 324405 127059 324471 127062
rect 307661 126850 307727 126853
rect 307661 126848 310132 126850
rect 307661 126792 307666 126848
rect 307722 126792 310132 126848
rect 307661 126790 310132 126792
rect 307661 126787 307727 126790
rect 214005 126714 214071 126717
rect 252461 126714 252527 126717
rect 214005 126712 217212 126714
rect 214005 126656 214010 126712
rect 214066 126656 217212 126712
rect 214005 126654 217212 126656
rect 248860 126712 252527 126714
rect 248860 126656 252466 126712
rect 252522 126656 252527 126712
rect 248860 126654 252527 126656
rect 214005 126651 214071 126654
rect 252461 126651 252527 126654
rect 397453 126714 397519 126717
rect 452561 126714 452627 126717
rect 397453 126712 400108 126714
rect 397453 126656 397458 126712
rect 397514 126656 400108 126712
rect 397453 126654 400108 126656
rect 449788 126712 452627 126714
rect 449788 126656 452566 126712
rect 452622 126656 452627 126712
rect 449788 126654 452627 126656
rect 397453 126651 397519 126654
rect 452561 126651 452627 126654
rect 301446 126380 301452 126444
rect 301516 126442 301522 126444
rect 301516 126382 310132 126442
rect 301516 126380 301522 126382
rect 67633 126306 67699 126309
rect 68142 126306 68816 126312
rect 67633 126304 68816 126306
rect 67633 126248 67638 126304
rect 67694 126252 68816 126304
rect 251766 126306 251772 126308
rect 67694 126248 68202 126252
rect 67633 126246 68202 126248
rect 67633 126243 67699 126246
rect 248860 126246 251772 126306
rect 251766 126244 251772 126246
rect 251836 126244 251842 126308
rect 325601 126306 325667 126309
rect 321908 126304 325667 126306
rect 321908 126248 325606 126304
rect 325662 126248 325667 126304
rect 321908 126246 325667 126248
rect 325601 126243 325667 126246
rect 213913 126034 213979 126037
rect 397545 126034 397611 126037
rect 580257 126034 580323 126037
rect 583520 126034 584960 126124
rect 213913 126032 217212 126034
rect 213913 125976 213918 126032
rect 213974 125976 217212 126032
rect 213913 125974 217212 125976
rect 397545 126032 400108 126034
rect 397545 125976 397550 126032
rect 397606 125976 400108 126032
rect 397545 125974 400108 125976
rect 580257 126032 584960 126034
rect 580257 125976 580262 126032
rect 580318 125976 584960 126032
rect 580257 125974 584960 125976
rect 213913 125971 213979 125974
rect 397545 125971 397611 125974
rect 580257 125971 580323 125974
rect 306741 125898 306807 125901
rect 306741 125896 310132 125898
rect 306741 125840 306746 125896
rect 306802 125840 310132 125896
rect 583520 125884 584960 125974
rect 306741 125838 310132 125840
rect 306741 125835 306807 125838
rect 252093 125762 252159 125765
rect 248860 125760 252159 125762
rect 248860 125704 252098 125760
rect 252154 125704 252159 125760
rect 248860 125702 252159 125704
rect 252093 125699 252159 125702
rect 306741 125490 306807 125493
rect 322974 125490 322980 125492
rect 306741 125488 310132 125490
rect 306741 125432 306746 125488
rect 306802 125432 310132 125488
rect 306741 125430 310132 125432
rect 321908 125430 322980 125490
rect 306741 125427 306807 125430
rect 322974 125428 322980 125430
rect 323044 125428 323050 125492
rect 214005 125354 214071 125357
rect 251909 125354 251975 125357
rect 214005 125352 217212 125354
rect 214005 125296 214010 125352
rect 214066 125296 217212 125352
rect 214005 125294 217212 125296
rect 248860 125352 251975 125354
rect 248860 125296 251914 125352
rect 251970 125296 251975 125352
rect 248860 125294 251975 125296
rect 214005 125291 214071 125294
rect 251909 125291 251975 125294
rect 397453 125354 397519 125357
rect 451549 125354 451615 125357
rect 452561 125354 452627 125357
rect 397453 125352 400108 125354
rect 397453 125296 397458 125352
rect 397514 125296 400108 125352
rect 397453 125294 400108 125296
rect 449788 125352 452627 125354
rect 449788 125296 451554 125352
rect 451610 125296 452566 125352
rect 452622 125296 452627 125352
rect 449788 125294 452627 125296
rect 397453 125291 397519 125294
rect 451549 125291 451615 125294
rect 452561 125291 452627 125294
rect 67541 125218 67607 125221
rect 68142 125218 68816 125224
rect 67541 125216 68816 125218
rect 67541 125160 67546 125216
rect 67602 125164 68816 125216
rect 67602 125160 68202 125164
rect 67541 125158 68202 125160
rect 67541 125155 67607 125158
rect -960 123572 480 123812
rect 307661 125082 307727 125085
rect 307661 125080 310132 125082
rect 307661 125024 307666 125080
rect 307722 125024 310132 125080
rect 307661 125022 310132 125024
rect 307661 125019 307727 125022
rect 252461 124810 252527 124813
rect 324313 124810 324379 124813
rect 248860 124808 252527 124810
rect 248860 124752 252466 124808
rect 252522 124752 252527 124808
rect 248860 124750 252527 124752
rect 321908 124808 324379 124810
rect 321908 124752 324318 124808
rect 324374 124752 324379 124808
rect 321908 124750 324379 124752
rect 252461 124747 252527 124750
rect 324313 124747 324379 124750
rect 213913 124674 213979 124677
rect 307017 124674 307083 124677
rect 451273 124674 451339 124677
rect 213913 124672 217212 124674
rect 213913 124616 213918 124672
rect 213974 124616 217212 124672
rect 213913 124614 217212 124616
rect 307017 124672 310132 124674
rect 307017 124616 307022 124672
rect 307078 124616 310132 124672
rect 307017 124614 310132 124616
rect 449788 124672 451339 124674
rect 449788 124616 451278 124672
rect 451334 124616 451339 124672
rect 449788 124614 451339 124616
rect 213913 124611 213979 124614
rect 307017 124611 307083 124614
rect 451273 124611 451339 124614
rect 251357 124402 251423 124405
rect 248860 124400 251423 124402
rect 248860 124344 251362 124400
rect 251418 124344 251423 124400
rect 248860 124342 251423 124344
rect 251357 124339 251423 124342
rect 307109 124266 307175 124269
rect 307109 124264 310132 124266
rect 307109 124208 307114 124264
rect 307170 124208 310132 124264
rect 307109 124206 310132 124208
rect 307109 124203 307175 124206
rect 214005 124130 214071 124133
rect 214005 124128 217212 124130
rect 214005 124072 214010 124128
rect 214066 124072 217212 124128
rect 214005 124070 217212 124072
rect 214005 124067 214071 124070
rect 252461 123994 252527 123997
rect 451641 123994 451707 123997
rect 248860 123992 252527 123994
rect 248860 123936 252466 123992
rect 252522 123936 252527 123992
rect 449788 123992 451707 123994
rect 248860 123934 252527 123936
rect 252461 123931 252527 123934
rect 306557 123858 306623 123861
rect 306557 123856 310132 123858
rect 306557 123800 306562 123856
rect 306618 123800 310132 123856
rect 306557 123798 310132 123800
rect 306557 123795 306623 123798
rect 67449 123586 67515 123589
rect 68142 123586 68816 123592
rect 67449 123584 68816 123586
rect 67449 123528 67454 123584
rect 67510 123532 68816 123584
rect 67510 123528 68202 123532
rect 67449 123526 68202 123528
rect 67449 123523 67515 123526
rect 213913 123450 213979 123453
rect 252369 123450 252435 123453
rect 213913 123448 217212 123450
rect 213913 123392 213918 123448
rect 213974 123392 217212 123448
rect 213913 123390 217212 123392
rect 248860 123448 252435 123450
rect 248860 123392 252374 123448
rect 252430 123392 252435 123448
rect 248860 123390 252435 123392
rect 213913 123387 213979 123390
rect 252369 123387 252435 123390
rect 307109 123450 307175 123453
rect 321878 123450 321938 123964
rect 449788 123936 451646 123992
rect 451702 123936 451707 123992
rect 449788 123934 451707 123936
rect 451641 123931 451707 123934
rect 397453 123858 397519 123861
rect 397453 123856 400108 123858
rect 397453 123800 397458 123856
rect 397514 123800 400108 123856
rect 397453 123798 400108 123800
rect 397453 123795 397519 123798
rect 323485 123450 323551 123453
rect 307109 123448 310132 123450
rect 307109 123392 307114 123448
rect 307170 123392 310132 123448
rect 307109 123390 310132 123392
rect 321878 123448 323551 123450
rect 321878 123392 323490 123448
rect 323546 123392 323551 123448
rect 321878 123390 323551 123392
rect 307109 123387 307175 123390
rect 323485 123387 323551 123390
rect 398189 123178 398255 123181
rect 321908 123118 325710 123178
rect 251173 123042 251239 123045
rect 248860 123040 251239 123042
rect 248860 122984 251178 123040
rect 251234 122984 251239 123040
rect 248860 122982 251239 122984
rect 251173 122979 251239 122982
rect 307661 123042 307727 123045
rect 325650 123042 325710 123118
rect 398189 123176 400108 123178
rect 398189 123120 398194 123176
rect 398250 123120 400108 123176
rect 398189 123118 400108 123120
rect 398189 123115 398255 123118
rect 329046 123042 329052 123044
rect 307661 123040 310132 123042
rect 307661 122984 307666 123040
rect 307722 122984 310132 123040
rect 307661 122982 310132 122984
rect 325650 122982 329052 123042
rect 307661 122979 307727 122982
rect 329046 122980 329052 122982
rect 329116 122980 329122 123044
rect 323485 122906 323551 122909
rect 335670 122906 335676 122908
rect 323485 122904 335676 122906
rect 323485 122848 323490 122904
rect 323546 122848 335676 122904
rect 323485 122846 335676 122848
rect 323485 122843 323551 122846
rect 335670 122844 335676 122846
rect 335740 122844 335746 122908
rect 214005 122770 214071 122773
rect 214005 122768 217212 122770
rect 214005 122712 214010 122768
rect 214066 122712 217212 122768
rect 214005 122710 217212 122712
rect 214005 122707 214071 122710
rect 66069 122634 66135 122637
rect 68142 122634 68816 122640
rect 66069 122632 68816 122634
rect 66069 122576 66074 122632
rect 66130 122580 68816 122632
rect 452561 122634 452627 122637
rect 66130 122576 68202 122580
rect 66069 122574 68202 122576
rect 66069 122571 66135 122574
rect 449788 122632 452627 122634
rect 449788 122576 452566 122632
rect 452622 122576 452627 122632
rect 449788 122574 452627 122576
rect 452561 122571 452627 122574
rect 252461 122498 252527 122501
rect 248860 122496 252527 122498
rect 248860 122440 252466 122496
rect 252522 122440 252527 122496
rect 248860 122438 252527 122440
rect 252461 122435 252527 122438
rect 307477 122498 307543 122501
rect 324313 122498 324379 122501
rect 307477 122496 310132 122498
rect 307477 122440 307482 122496
rect 307538 122440 310132 122496
rect 307477 122438 310132 122440
rect 321908 122496 324379 122498
rect 321908 122440 324318 122496
rect 324374 122440 324379 122496
rect 321908 122438 324379 122440
rect 307477 122435 307543 122438
rect 324313 122435 324379 122438
rect 321645 122226 321711 122229
rect 321645 122224 321754 122226
rect 321645 122168 321650 122224
rect 321706 122168 321754 122224
rect 321645 122163 321754 122168
rect 213913 122090 213979 122093
rect 251357 122090 251423 122093
rect 213913 122088 217212 122090
rect 213913 122032 213918 122088
rect 213974 122032 217212 122088
rect 213913 122030 217212 122032
rect 248860 122088 251423 122090
rect 248860 122032 251362 122088
rect 251418 122032 251423 122088
rect 248860 122030 251423 122032
rect 213913 122027 213979 122030
rect 251357 122027 251423 122030
rect 307569 122090 307635 122093
rect 307569 122088 310132 122090
rect 307569 122032 307574 122088
rect 307630 122032 310132 122088
rect 307569 122030 310132 122032
rect 307569 122027 307635 122030
rect 307661 121682 307727 121685
rect 307661 121680 310132 121682
rect 307661 121624 307666 121680
rect 307722 121624 310132 121680
rect 321694 121652 321754 122163
rect 397453 121954 397519 121957
rect 397453 121952 400108 121954
rect 397453 121896 397458 121952
rect 397514 121896 400108 121952
rect 397453 121894 400108 121896
rect 397453 121891 397519 121894
rect 307661 121622 310132 121624
rect 307661 121619 307727 121622
rect 252001 121546 252067 121549
rect 248860 121544 252067 121546
rect 248860 121488 252006 121544
rect 252062 121488 252067 121544
rect 248860 121486 252067 121488
rect 449758 121546 449818 121788
rect 451038 121546 451044 121548
rect 449758 121486 451044 121546
rect 252001 121483 252067 121486
rect 451038 121484 451044 121486
rect 451108 121484 451114 121548
rect 214005 121410 214071 121413
rect 214005 121408 217212 121410
rect 214005 121352 214010 121408
rect 214066 121352 217212 121408
rect 214005 121350 217212 121352
rect 214005 121347 214071 121350
rect 306741 121274 306807 121277
rect 397453 121274 397519 121277
rect 306741 121272 310132 121274
rect 306741 121216 306746 121272
rect 306802 121216 310132 121272
rect 306741 121214 310132 121216
rect 397453 121272 400108 121274
rect 397453 121216 397458 121272
rect 397514 121216 400108 121272
rect 397453 121214 400108 121216
rect 306741 121211 306807 121214
rect 397453 121211 397519 121214
rect 252461 121138 252527 121141
rect 248860 121136 252527 121138
rect 248860 121080 252466 121136
rect 252522 121080 252527 121136
rect 248860 121078 252527 121080
rect 252461 121075 252527 121078
rect 67357 120866 67423 120869
rect 68142 120866 68816 120872
rect 67357 120864 68816 120866
rect 67357 120808 67362 120864
rect 67418 120812 68816 120864
rect 67418 120808 68202 120812
rect 67357 120806 68202 120808
rect 67357 120803 67423 120806
rect 307569 120866 307635 120869
rect 324313 120866 324379 120869
rect 307569 120864 310132 120866
rect 307569 120808 307574 120864
rect 307630 120808 310132 120864
rect 307569 120806 310132 120808
rect 321908 120864 324379 120866
rect 321908 120808 324318 120864
rect 324374 120808 324379 120864
rect 321908 120806 324379 120808
rect 307569 120803 307635 120806
rect 324313 120803 324379 120806
rect 213913 120730 213979 120733
rect 213913 120728 217212 120730
rect 213913 120672 213918 120728
rect 213974 120672 217212 120728
rect 213913 120670 217212 120672
rect 213913 120667 213979 120670
rect 251817 120594 251883 120597
rect 248860 120592 251883 120594
rect 248860 120536 251822 120592
rect 251878 120536 251883 120592
rect 248860 120534 251883 120536
rect 251817 120531 251883 120534
rect 307661 120458 307727 120461
rect 450077 120458 450143 120461
rect 307661 120456 310132 120458
rect 307661 120400 307666 120456
rect 307722 120400 310132 120456
rect 307661 120398 310132 120400
rect 449788 120456 450143 120458
rect 449788 120400 450082 120456
rect 450138 120400 450143 120456
rect 449788 120398 450143 120400
rect 307661 120395 307727 120398
rect 450077 120395 450143 120398
rect 252277 120186 252343 120189
rect 324405 120186 324471 120189
rect 248860 120184 252343 120186
rect 248860 120128 252282 120184
rect 252338 120128 252343 120184
rect 248860 120126 252343 120128
rect 321908 120184 324471 120186
rect 321908 120128 324410 120184
rect 324466 120128 324471 120184
rect 321908 120126 324471 120128
rect 252277 120123 252343 120126
rect 324405 120123 324471 120126
rect 214005 120050 214071 120053
rect 307569 120050 307635 120053
rect 214005 120048 217212 120050
rect 214005 119992 214010 120048
rect 214066 119992 217212 120048
rect 214005 119990 217212 119992
rect 307569 120048 310132 120050
rect 307569 119992 307574 120048
rect 307630 119992 310132 120048
rect 307569 119990 310132 119992
rect 214005 119987 214071 119990
rect 307569 119987 307635 119990
rect 397453 119914 397519 119917
rect 397453 119912 400108 119914
rect 397453 119856 397458 119912
rect 397514 119856 400108 119912
rect 397453 119854 400108 119856
rect 397453 119851 397519 119854
rect 251357 119642 251423 119645
rect 248860 119640 251423 119642
rect 248860 119584 251362 119640
rect 251418 119584 251423 119640
rect 248860 119582 251423 119584
rect 251357 119579 251423 119582
rect 307477 119642 307543 119645
rect 307477 119640 310132 119642
rect 307477 119584 307482 119640
rect 307538 119584 310132 119640
rect 307477 119582 310132 119584
rect 307477 119579 307543 119582
rect 213913 119506 213979 119509
rect 213913 119504 217212 119506
rect 213913 119448 213918 119504
rect 213974 119448 217212 119504
rect 213913 119446 217212 119448
rect 213913 119443 213979 119446
rect 324313 119370 324379 119373
rect 321908 119368 324379 119370
rect 321908 119312 324318 119368
rect 324374 119312 324379 119368
rect 321908 119310 324379 119312
rect 324313 119307 324379 119310
rect 252461 119234 252527 119237
rect 248860 119232 252527 119234
rect 248860 119176 252466 119232
rect 252522 119176 252527 119232
rect 248860 119174 252527 119176
rect 252461 119171 252527 119174
rect 307661 119098 307727 119101
rect 396717 119098 396783 119101
rect 307661 119096 310132 119098
rect 307661 119040 307666 119096
rect 307722 119040 310132 119096
rect 307661 119038 310132 119040
rect 396717 119096 400108 119098
rect 396717 119040 396722 119096
rect 396778 119040 400108 119096
rect 396717 119038 400108 119040
rect 307661 119035 307727 119038
rect 396717 119035 396783 119038
rect 214097 118826 214163 118829
rect 252277 118826 252343 118829
rect 214097 118824 217212 118826
rect 214097 118768 214102 118824
rect 214158 118768 217212 118824
rect 214097 118766 217212 118768
rect 248860 118824 252343 118826
rect 248860 118768 252282 118824
rect 252338 118768 252343 118824
rect 248860 118766 252343 118768
rect 449758 118826 449818 119748
rect 458766 118826 458772 118828
rect 449758 118766 458772 118826
rect 214097 118763 214163 118766
rect 252277 118763 252343 118766
rect 458766 118764 458772 118766
rect 458836 118764 458842 118828
rect 307569 118690 307635 118693
rect 307569 118688 310132 118690
rect 307569 118632 307574 118688
rect 307630 118632 310132 118688
rect 307569 118630 310132 118632
rect 307569 118627 307635 118630
rect 324957 118554 325023 118557
rect 321908 118552 325023 118554
rect 321908 118496 324962 118552
rect 325018 118496 325023 118552
rect 321908 118494 325023 118496
rect 324957 118491 325023 118494
rect 252461 118282 252527 118285
rect 248860 118280 252527 118282
rect 248860 118224 252466 118280
rect 252522 118224 252527 118280
rect 248860 118222 252527 118224
rect 252461 118219 252527 118222
rect 306557 118282 306623 118285
rect 306557 118280 310132 118282
rect 306557 118224 306562 118280
rect 306618 118224 310132 118280
rect 306557 118222 310132 118224
rect 306557 118219 306623 118222
rect 214005 118146 214071 118149
rect 449758 118146 449818 118388
rect 454166 118146 454172 118148
rect 214005 118144 217212 118146
rect 214005 118088 214010 118144
rect 214066 118088 217212 118144
rect 214005 118086 217212 118088
rect 449758 118086 454172 118146
rect 214005 118083 214071 118086
rect 454166 118084 454172 118086
rect 454236 118084 454242 118148
rect 251817 117874 251883 117877
rect 248860 117872 251883 117874
rect 248860 117816 251822 117872
rect 251878 117816 251883 117872
rect 248860 117814 251883 117816
rect 251817 117811 251883 117814
rect 307661 117874 307727 117877
rect 324313 117874 324379 117877
rect 307661 117872 310132 117874
rect 307661 117816 307666 117872
rect 307722 117816 310132 117872
rect 307661 117814 310132 117816
rect 321908 117872 324379 117874
rect 321908 117816 324318 117872
rect 324374 117816 324379 117872
rect 321908 117814 324379 117816
rect 307661 117811 307727 117814
rect 324313 117811 324379 117814
rect 398281 117874 398347 117877
rect 452469 117874 452535 117877
rect 398281 117872 400108 117874
rect 398281 117816 398286 117872
rect 398342 117816 400108 117872
rect 398281 117814 400108 117816
rect 449788 117872 452535 117874
rect 449788 117816 452474 117872
rect 452530 117816 452535 117872
rect 449788 117814 452535 117816
rect 398281 117811 398347 117814
rect 452469 117811 452535 117814
rect 213913 117466 213979 117469
rect 307661 117466 307727 117469
rect 213913 117464 217212 117466
rect 213913 117408 213918 117464
rect 213974 117408 217212 117464
rect 213913 117406 217212 117408
rect 307661 117464 310132 117466
rect 307661 117408 307666 117464
rect 307722 117408 310132 117464
rect 307661 117406 310132 117408
rect 213913 117403 213979 117406
rect 307661 117403 307727 117406
rect 251725 117330 251791 117333
rect 248860 117328 251791 117330
rect 248860 117272 251730 117328
rect 251786 117272 251791 117328
rect 248860 117270 251791 117272
rect 251725 117267 251791 117270
rect 346342 117268 346348 117332
rect 346412 117330 346418 117332
rect 347221 117330 347287 117333
rect 346412 117328 347287 117330
rect 346412 117272 347226 117328
rect 347282 117272 347287 117328
rect 346412 117270 347287 117272
rect 346412 117268 346418 117270
rect 347221 117267 347287 117270
rect 397453 117194 397519 117197
rect 397453 117192 400108 117194
rect 397453 117136 397458 117192
rect 397514 117136 400108 117192
rect 397453 117134 400108 117136
rect 397453 117131 397519 117134
rect 306741 117058 306807 117061
rect 323158 117058 323164 117060
rect 306741 117056 310132 117058
rect 306741 117000 306746 117056
rect 306802 117000 310132 117056
rect 306741 116998 310132 117000
rect 321908 116998 323164 117058
rect 306741 116995 306807 116998
rect 323158 116996 323164 116998
rect 323228 116996 323234 117060
rect 449341 117058 449407 117061
rect 449341 117056 449450 117058
rect 449341 117000 449346 117056
rect 449402 117000 449450 117056
rect 449341 116995 449450 117000
rect 251357 116922 251423 116925
rect 248860 116920 251423 116922
rect 248860 116864 251362 116920
rect 251418 116864 251423 116920
rect 248860 116862 251423 116864
rect 251357 116859 251423 116862
rect 214005 116786 214071 116789
rect 214005 116784 217212 116786
rect 214005 116728 214010 116784
rect 214066 116728 217212 116784
rect 214005 116726 217212 116728
rect 214005 116723 214071 116726
rect 307477 116650 307543 116653
rect 307477 116648 310132 116650
rect 307477 116592 307482 116648
rect 307538 116592 310132 116648
rect 307477 116590 310132 116592
rect 307477 116587 307543 116590
rect 398925 116514 398991 116517
rect 398925 116512 400108 116514
rect 398925 116456 398930 116512
rect 398986 116456 400108 116512
rect 449390 116484 449450 116995
rect 398925 116454 400108 116456
rect 398925 116451 398991 116454
rect 252369 116378 252435 116381
rect 324313 116378 324379 116381
rect 248860 116376 252435 116378
rect 248860 116320 252374 116376
rect 252430 116320 252435 116376
rect 248860 116318 252435 116320
rect 321908 116376 324379 116378
rect 321908 116320 324318 116376
rect 324374 116320 324379 116376
rect 321908 116318 324379 116320
rect 252369 116315 252435 116318
rect 324313 116315 324379 116318
rect 307293 116242 307359 116245
rect 307293 116240 310132 116242
rect 307293 116184 307298 116240
rect 307354 116184 310132 116240
rect 307293 116182 310132 116184
rect 307293 116179 307359 116182
rect 213913 116106 213979 116109
rect 213913 116104 217212 116106
rect 213913 116048 213918 116104
rect 213974 116048 217212 116104
rect 213913 116046 217212 116048
rect 213913 116043 213979 116046
rect 252461 115970 252527 115973
rect 248860 115968 252527 115970
rect 248860 115912 252466 115968
rect 252522 115912 252527 115968
rect 248860 115910 252527 115912
rect 252461 115907 252527 115910
rect 451549 115834 451615 115837
rect 449788 115832 451615 115834
rect 449788 115776 451554 115832
rect 451610 115776 451615 115832
rect 449788 115774 451615 115776
rect 451549 115771 451615 115774
rect 307109 115698 307175 115701
rect 307109 115696 310132 115698
rect 307109 115640 307114 115696
rect 307170 115640 310132 115696
rect 307109 115638 310132 115640
rect 307109 115635 307175 115638
rect 324313 115562 324379 115565
rect 321908 115560 324379 115562
rect 321908 115504 324318 115560
rect 324374 115504 324379 115560
rect 321908 115502 324379 115504
rect 324313 115499 324379 115502
rect 214005 115426 214071 115429
rect 252277 115426 252343 115429
rect 214005 115424 217212 115426
rect 214005 115368 214010 115424
rect 214066 115368 217212 115424
rect 214005 115366 217212 115368
rect 248860 115424 252343 115426
rect 248860 115368 252282 115424
rect 252338 115368 252343 115424
rect 248860 115366 252343 115368
rect 214005 115363 214071 115366
rect 252277 115363 252343 115366
rect 307569 115290 307635 115293
rect 307569 115288 310132 115290
rect 307569 115232 307574 115288
rect 307630 115232 310132 115288
rect 307569 115230 310132 115232
rect 307569 115227 307635 115230
rect 397453 115154 397519 115157
rect 397453 115152 400108 115154
rect 397453 115096 397458 115152
rect 397514 115096 400108 115152
rect 397453 115094 400108 115096
rect 397453 115091 397519 115094
rect 251909 115018 251975 115021
rect 451365 115018 451431 115021
rect 248860 115016 251975 115018
rect 248860 114960 251914 115016
rect 251970 114960 251975 115016
rect 248860 114958 251975 114960
rect 449788 115016 451431 115018
rect 449788 114960 451370 115016
rect 451426 114960 451431 115016
rect 449788 114958 451431 114960
rect 251909 114955 251975 114958
rect 451365 114955 451431 114958
rect 213913 114882 213979 114885
rect 307661 114882 307727 114885
rect 213913 114880 217212 114882
rect 213913 114824 213918 114880
rect 213974 114824 217212 114880
rect 213913 114822 217212 114824
rect 307661 114880 310132 114882
rect 307661 114824 307666 114880
rect 307722 114824 310132 114880
rect 307661 114822 310132 114824
rect 213913 114819 213979 114822
rect 307661 114819 307727 114822
rect 321908 114686 325710 114746
rect 325650 114610 325710 114686
rect 329782 114610 329788 114612
rect 325650 114550 329788 114610
rect 329782 114548 329788 114550
rect 329852 114548 329858 114612
rect 251725 114474 251791 114477
rect 248860 114472 251791 114474
rect 248860 114416 251730 114472
rect 251786 114416 251791 114472
rect 248860 114414 251791 114416
rect 251725 114411 251791 114414
rect 306925 114474 306991 114477
rect 397453 114474 397519 114477
rect 306925 114472 310132 114474
rect 306925 114416 306930 114472
rect 306986 114416 310132 114472
rect 306925 114414 310132 114416
rect 397453 114472 400108 114474
rect 397453 114416 397458 114472
rect 397514 114416 400108 114472
rect 397453 114414 400108 114416
rect 306925 114411 306991 114414
rect 397453 114411 397519 114414
rect 214005 114202 214071 114205
rect 214005 114200 217212 114202
rect 214005 114144 214010 114200
rect 214066 114144 217212 114200
rect 214005 114142 217212 114144
rect 214005 114139 214071 114142
rect 251633 114066 251699 114069
rect 248860 114064 251699 114066
rect 248860 114008 251638 114064
rect 251694 114008 251699 114064
rect 248860 114006 251699 114008
rect 251633 114003 251699 114006
rect 306557 114066 306623 114069
rect 324313 114066 324379 114069
rect 306557 114064 310132 114066
rect 306557 114008 306562 114064
rect 306618 114008 310132 114064
rect 306557 114006 310132 114008
rect 321908 114064 324379 114066
rect 321908 114008 324318 114064
rect 324374 114008 324379 114064
rect 321908 114006 324379 114008
rect 306557 114003 306623 114006
rect 324313 114003 324379 114006
rect 271781 113930 271847 113933
rect 291694 113930 291700 113932
rect 271781 113928 291700 113930
rect 271781 113872 271786 113928
rect 271842 113872 291700 113928
rect 271781 113870 291700 113872
rect 271781 113867 271847 113870
rect 291694 113868 291700 113870
rect 291764 113868 291770 113932
rect 252502 113732 252508 113796
rect 252572 113794 252578 113796
rect 278129 113794 278195 113797
rect 452469 113794 452535 113797
rect 252572 113792 278195 113794
rect 252572 113736 278134 113792
rect 278190 113736 278195 113792
rect 252572 113734 278195 113736
rect 449788 113792 452535 113794
rect 449788 113736 452474 113792
rect 452530 113736 452535 113792
rect 449788 113734 452535 113736
rect 252572 113732 252578 113734
rect 278129 113731 278195 113734
rect 452469 113731 452535 113734
rect 305678 113596 305684 113660
rect 305748 113658 305754 113660
rect 305748 113598 310132 113658
rect 305748 113596 305754 113598
rect 213913 113522 213979 113525
rect 251357 113522 251423 113525
rect 213913 113520 217212 113522
rect 213913 113464 213918 113520
rect 213974 113464 217212 113520
rect 213913 113462 217212 113464
rect 248860 113520 251423 113522
rect 248860 113464 251362 113520
rect 251418 113464 251423 113520
rect 248860 113462 251423 113464
rect 213913 113459 213979 113462
rect 251357 113459 251423 113462
rect 307661 113250 307727 113253
rect 324405 113250 324471 113253
rect 307661 113248 310132 113250
rect 307661 113192 307666 113248
rect 307722 113192 310132 113248
rect 307661 113190 310132 113192
rect 321908 113248 324471 113250
rect 321908 113192 324410 113248
rect 324466 113192 324471 113248
rect 321908 113190 324471 113192
rect 307661 113187 307727 113190
rect 324405 113187 324471 113190
rect 252461 113114 252527 113117
rect 248860 113112 252527 113114
rect 248860 113056 252466 113112
rect 252522 113056 252527 113112
rect 248860 113054 252527 113056
rect 252461 113051 252527 113054
rect 397453 113114 397519 113117
rect 397453 113112 400108 113114
rect 397453 113056 397458 113112
rect 397514 113056 400108 113112
rect 397453 113054 400108 113056
rect 397453 113051 397519 113054
rect 214005 112842 214071 112845
rect 214005 112840 217212 112842
rect 214005 112784 214010 112840
rect 214066 112784 217212 112840
rect 214005 112782 217212 112784
rect 214005 112779 214071 112782
rect 252461 112706 252527 112709
rect 248860 112704 252527 112706
rect 248860 112648 252466 112704
rect 252522 112648 252527 112704
rect 248860 112646 252527 112648
rect 252461 112643 252527 112646
rect 299974 112644 299980 112708
rect 300044 112706 300050 112708
rect 300044 112646 310132 112706
rect 300044 112644 300050 112646
rect 326337 112434 326403 112437
rect 396574 112434 396580 112436
rect 326337 112432 396580 112434
rect 307477 112298 307543 112301
rect 307477 112296 310132 112298
rect 307477 112240 307482 112296
rect 307538 112240 310132 112296
rect 307477 112238 310132 112240
rect 307477 112235 307543 112238
rect 213913 112162 213979 112165
rect 251633 112162 251699 112165
rect 213913 112160 217212 112162
rect 213913 112104 213918 112160
rect 213974 112104 217212 112160
rect 213913 112102 217212 112104
rect 248860 112160 251699 112162
rect 248860 112104 251638 112160
rect 251694 112104 251699 112160
rect 248860 112102 251699 112104
rect 213913 112099 213979 112102
rect 251633 112099 251699 112102
rect 307661 111890 307727 111893
rect 321878 111890 321938 112404
rect 326337 112376 326342 112432
rect 326398 112376 396580 112432
rect 326337 112374 396580 112376
rect 326337 112371 326403 112374
rect 396574 112372 396580 112374
rect 396644 112372 396650 112436
rect 449758 112434 449818 112948
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect 449934 112434 449940 112436
rect 449758 112374 449940 112434
rect 449934 112372 449940 112374
rect 450004 112372 450010 112436
rect 331254 111890 331260 111892
rect 307661 111888 310132 111890
rect 307661 111832 307666 111888
rect 307722 111832 310132 111888
rect 307661 111830 310132 111832
rect 321878 111830 331260 111890
rect 307661 111827 307727 111830
rect 331254 111828 331260 111830
rect 331324 111828 331330 111892
rect 399569 111890 399635 111893
rect 400078 111890 400138 112268
rect 399569 111888 400138 111890
rect 399569 111832 399574 111888
rect 399630 111832 400138 111888
rect 399569 111830 400138 111832
rect 399569 111827 399635 111830
rect 168281 111754 168347 111757
rect 252093 111754 252159 111757
rect 452561 111754 452627 111757
rect 164694 111752 168347 111754
rect 164694 111696 168286 111752
rect 168342 111696 168347 111752
rect 164694 111694 168347 111696
rect 248860 111752 252159 111754
rect 248860 111696 252098 111752
rect 252154 111696 252159 111752
rect 449788 111752 452627 111754
rect 248860 111694 252159 111696
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 168281 111691 168347 111694
rect 252093 111691 252159 111694
rect 213913 111482 213979 111485
rect 307477 111482 307543 111485
rect 213913 111480 217212 111482
rect 213913 111424 213918 111480
rect 213974 111424 217212 111480
rect 213913 111422 217212 111424
rect 307477 111480 310132 111482
rect 307477 111424 307482 111480
rect 307538 111424 310132 111480
rect 307477 111422 310132 111424
rect 213913 111419 213979 111422
rect 307477 111419 307543 111422
rect 252001 111210 252067 111213
rect 248860 111208 252067 111210
rect 248860 111152 252006 111208
rect 252062 111152 252067 111208
rect 248860 111150 252067 111152
rect 252001 111147 252067 111150
rect 307569 111074 307635 111077
rect 321878 111074 321938 111724
rect 449788 111696 452566 111752
rect 452622 111696 452627 111752
rect 449788 111694 452627 111696
rect 452561 111691 452627 111694
rect 334014 111074 334020 111076
rect 307569 111072 310132 111074
rect 307569 111016 307574 111072
rect 307630 111016 310132 111072
rect 307569 111014 310132 111016
rect 321878 111014 334020 111074
rect 307569 111011 307635 111014
rect 334014 111012 334020 111014
rect 334084 111012 334090 111076
rect 397453 111074 397519 111077
rect 452469 111074 452535 111077
rect 397453 111072 400108 111074
rect 397453 111016 397458 111072
rect 397514 111016 400108 111072
rect 397453 111014 400108 111016
rect 449788 111072 452535 111074
rect 449788 111016 452474 111072
rect 452530 111016 452535 111072
rect 449788 111014 452535 111016
rect 397453 111011 397519 111014
rect 452469 111011 452535 111014
rect 324957 110938 325023 110941
rect 321908 110936 325023 110938
rect 321908 110880 324962 110936
rect 325018 110880 325023 110936
rect 321908 110878 325023 110880
rect 324957 110875 325023 110878
rect 214741 110802 214807 110805
rect 252502 110802 252508 110804
rect 214741 110800 217212 110802
rect 214741 110744 214746 110800
rect 214802 110744 217212 110800
rect 214741 110742 217212 110744
rect 248860 110742 252508 110802
rect 214741 110739 214807 110742
rect 252502 110740 252508 110742
rect 252572 110740 252578 110804
rect 307661 110666 307727 110669
rect 307661 110664 310132 110666
rect 307661 110608 307666 110664
rect 307722 110608 310132 110664
rect 307661 110606 310132 110608
rect 307661 110603 307727 110606
rect 397453 110394 397519 110397
rect 397453 110392 400108 110394
rect 397453 110336 397458 110392
rect 397514 110336 400108 110392
rect 397453 110334 400108 110336
rect 397453 110331 397519 110334
rect 214005 110258 214071 110261
rect 251909 110258 251975 110261
rect 214005 110256 217212 110258
rect 214005 110200 214010 110256
rect 214066 110200 217212 110256
rect 214005 110198 217212 110200
rect 248860 110256 251975 110258
rect 248860 110200 251914 110256
rect 251970 110200 251975 110256
rect 248860 110198 251975 110200
rect 214005 110195 214071 110198
rect 251909 110195 251975 110198
rect 307477 110258 307543 110261
rect 307477 110256 310132 110258
rect 307477 110200 307482 110256
rect 307538 110200 310132 110256
rect 307477 110198 310132 110200
rect 307477 110195 307543 110198
rect 167821 110122 167887 110125
rect 324313 110122 324379 110125
rect 164694 110120 167887 110122
rect 164694 110064 167826 110120
rect 167882 110064 167887 110120
rect 164694 110062 167887 110064
rect 321908 110120 324379 110122
rect 321908 110064 324318 110120
rect 324374 110064 324379 110120
rect 321908 110062 324379 110064
rect 167821 110059 167887 110062
rect 324313 110059 324379 110062
rect 252461 109850 252527 109853
rect 248860 109848 252527 109850
rect 248860 109792 252466 109848
rect 252522 109792 252527 109848
rect 248860 109790 252527 109792
rect 252461 109787 252527 109790
rect 307569 109850 307635 109853
rect 307569 109848 310132 109850
rect 307569 109792 307574 109848
rect 307630 109792 310132 109848
rect 307569 109790 310132 109792
rect 307569 109787 307635 109790
rect 452101 109714 452167 109717
rect 449788 109712 452167 109714
rect 449788 109656 452106 109712
rect 452162 109656 452167 109712
rect 449788 109654 452167 109656
rect 452101 109651 452167 109654
rect 213913 109578 213979 109581
rect 397729 109578 397795 109581
rect 213913 109576 217212 109578
rect 213913 109520 213918 109576
rect 213974 109520 217212 109576
rect 213913 109518 217212 109520
rect 397729 109576 400108 109578
rect 397729 109520 397734 109576
rect 397790 109520 400108 109576
rect 397729 109518 400108 109520
rect 213913 109515 213979 109518
rect 397729 109515 397795 109518
rect 252093 109306 252159 109309
rect 248860 109304 252159 109306
rect 248860 109248 252098 109304
rect 252154 109248 252159 109304
rect 248860 109246 252159 109248
rect 252093 109243 252159 109246
rect 307661 109306 307727 109309
rect 307661 109304 310132 109306
rect 307661 109248 307666 109304
rect 307722 109248 310132 109304
rect 307661 109246 310132 109248
rect 307661 109243 307727 109246
rect 321510 109173 321570 109412
rect 251081 109170 251147 109173
rect 251214 109170 251220 109172
rect 251081 109168 251220 109170
rect 251081 109112 251086 109168
rect 251142 109112 251220 109168
rect 251081 109110 251220 109112
rect 251081 109107 251147 109110
rect 251214 109108 251220 109110
rect 251284 109108 251290 109172
rect 321510 109168 321619 109173
rect 321510 109112 321558 109168
rect 321614 109112 321619 109168
rect 321510 109110 321619 109112
rect 321553 109107 321619 109110
rect 451549 109034 451615 109037
rect 452837 109034 452903 109037
rect 449788 109032 452903 109034
rect 449788 108976 451554 109032
rect 451610 108976 452842 109032
rect 452898 108976 452903 109032
rect 449788 108974 452903 108976
rect 451549 108971 451615 108974
rect 452837 108971 452903 108974
rect 214005 108898 214071 108901
rect 252461 108898 252527 108901
rect 214005 108896 217212 108898
rect 214005 108840 214010 108896
rect 214066 108840 217212 108896
rect 214005 108838 217212 108840
rect 248860 108896 252527 108898
rect 248860 108840 252466 108896
rect 252522 108840 252527 108896
rect 248860 108838 252527 108840
rect 214005 108835 214071 108838
rect 252461 108835 252527 108838
rect 307477 108898 307543 108901
rect 307477 108896 310132 108898
rect 307477 108840 307482 108896
rect 307538 108840 310132 108896
rect 307477 108838 310132 108840
rect 307477 108835 307543 108838
rect 168097 108762 168163 108765
rect 164694 108760 168163 108762
rect 164694 108704 168102 108760
rect 168158 108704 168163 108760
rect 164694 108702 168163 108704
rect 168097 108699 168163 108702
rect 324262 108626 324268 108628
rect 321908 108566 324268 108626
rect 324262 108564 324268 108566
rect 324332 108626 324338 108628
rect 324405 108626 324471 108629
rect 324332 108624 324471 108626
rect 324332 108568 324410 108624
rect 324466 108568 324471 108624
rect 324332 108566 324471 108568
rect 324332 108564 324338 108566
rect 324405 108563 324471 108566
rect 307661 108490 307727 108493
rect 307661 108488 310132 108490
rect 307661 108432 307666 108488
rect 307722 108432 310132 108488
rect 307661 108430 310132 108432
rect 307661 108427 307727 108430
rect 252369 108354 252435 108357
rect 322054 108354 322060 108356
rect 248860 108352 252435 108354
rect 248860 108296 252374 108352
rect 252430 108296 252435 108352
rect 248860 108294 252435 108296
rect 252369 108291 252435 108294
rect 321878 108294 322060 108354
rect 213913 108218 213979 108221
rect 213913 108216 217212 108218
rect 213913 108160 213918 108216
rect 213974 108160 217212 108216
rect 213913 108158 217212 108160
rect 213913 108155 213979 108158
rect 307569 108082 307635 108085
rect 307569 108080 310132 108082
rect 307569 108024 307574 108080
rect 307630 108024 310132 108080
rect 307569 108022 310132 108024
rect 307569 108019 307635 108022
rect 252277 107946 252343 107949
rect 248860 107944 252343 107946
rect 248860 107888 252282 107944
rect 252338 107888 252343 107944
rect 248860 107886 252343 107888
rect 252277 107883 252343 107886
rect 321878 107780 321938 108294
rect 322054 108292 322060 108294
rect 322124 108354 322130 108356
rect 324313 108354 324379 108357
rect 322124 108352 324379 108354
rect 322124 108296 324318 108352
rect 324374 108296 324379 108352
rect 322124 108294 324379 108296
rect 322124 108292 322130 108294
rect 324313 108291 324379 108294
rect 397453 108218 397519 108221
rect 451733 108218 451799 108221
rect 397453 108216 400108 108218
rect 397453 108160 397458 108216
rect 397514 108160 400108 108216
rect 397453 108158 400108 108160
rect 449788 108216 451799 108218
rect 449788 108160 451738 108216
rect 451794 108160 451799 108216
rect 449788 108158 451799 108160
rect 397453 108155 397519 108158
rect 451733 108155 451799 108158
rect 305637 107674 305703 107677
rect 307477 107674 307543 107677
rect 305637 107672 307543 107674
rect 305637 107616 305642 107672
rect 305698 107616 307482 107672
rect 307538 107616 307543 107672
rect 305637 107614 307543 107616
rect 305637 107611 305703 107614
rect 307477 107611 307543 107614
rect 307661 107674 307727 107677
rect 307661 107672 310132 107674
rect 307661 107616 307666 107672
rect 307722 107616 310132 107672
rect 307661 107614 310132 107616
rect 307661 107611 307727 107614
rect 214005 107538 214071 107541
rect 252185 107538 252251 107541
rect 214005 107536 217212 107538
rect 214005 107480 214010 107536
rect 214066 107480 217212 107536
rect 214005 107478 217212 107480
rect 248860 107536 252251 107538
rect 248860 107480 252190 107536
rect 252246 107480 252251 107536
rect 248860 107478 252251 107480
rect 214005 107475 214071 107478
rect 252185 107475 252251 107478
rect 307477 107266 307543 107269
rect 307477 107264 310132 107266
rect 307477 107208 307482 107264
rect 307538 107208 310132 107264
rect 307477 107206 310132 107208
rect 307477 107203 307543 107206
rect 325049 107130 325115 107133
rect 321908 107128 325115 107130
rect 321908 107072 325054 107128
rect 325110 107072 325115 107128
rect 321908 107070 325115 107072
rect 325049 107067 325115 107070
rect 251817 106994 251883 106997
rect 248860 106992 251883 106994
rect 248860 106936 251822 106992
rect 251878 106936 251883 106992
rect 248860 106934 251883 106936
rect 251817 106931 251883 106934
rect 213913 106858 213979 106861
rect 307569 106858 307635 106861
rect 400078 106858 400138 107508
rect 452561 106994 452627 106997
rect 449788 106992 452627 106994
rect 449788 106936 452566 106992
rect 452622 106936 452627 106992
rect 449788 106934 452627 106936
rect 452561 106931 452627 106934
rect 213913 106856 217212 106858
rect 213913 106800 213918 106856
rect 213974 106800 217212 106856
rect 213913 106798 217212 106800
rect 307569 106856 310132 106858
rect 307569 106800 307574 106856
rect 307630 106800 310132 106856
rect 307569 106798 310132 106800
rect 393270 106798 400138 106858
rect 213913 106795 213979 106798
rect 307569 106795 307635 106798
rect 252093 106586 252159 106589
rect 248860 106584 252159 106586
rect 248860 106528 252098 106584
rect 252154 106528 252159 106584
rect 248860 106526 252159 106528
rect 252093 106523 252159 106526
rect 307661 106450 307727 106453
rect 307661 106448 310132 106450
rect 307661 106392 307666 106448
rect 307722 106392 310132 106448
rect 307661 106390 310132 106392
rect 307661 106387 307727 106390
rect 382774 106388 382780 106452
rect 382844 106450 382850 106452
rect 393270 106450 393330 106798
rect 382844 106390 393330 106450
rect 382844 106388 382850 106390
rect 305729 106314 305795 106317
rect 307477 106314 307543 106317
rect 322933 106314 322999 106317
rect 323301 106314 323367 106317
rect 305729 106312 307543 106314
rect 305729 106256 305734 106312
rect 305790 106256 307482 106312
rect 307538 106256 307543 106312
rect 305729 106254 307543 106256
rect 321908 106312 323367 106314
rect 321908 106256 322938 106312
rect 322994 106256 323306 106312
rect 323362 106256 323367 106312
rect 321908 106254 323367 106256
rect 305729 106251 305795 106254
rect 307477 106251 307543 106254
rect 322933 106251 322999 106254
rect 323301 106251 323367 106254
rect 397637 106314 397703 106317
rect 451273 106314 451339 106317
rect 397637 106312 400108 106314
rect 397637 106256 397642 106312
rect 397698 106256 400108 106312
rect 397637 106254 400108 106256
rect 449788 106312 451339 106314
rect 449788 106256 451278 106312
rect 451334 106256 451339 106312
rect 449788 106254 451339 106256
rect 397637 106251 397703 106254
rect 451273 106251 451339 106254
rect 213913 106178 213979 106181
rect 213913 106176 217212 106178
rect 213913 106120 213918 106176
rect 213974 106120 217212 106176
rect 213913 106118 217212 106120
rect 213913 106115 213979 106118
rect 251909 106042 251975 106045
rect 248860 106040 251975 106042
rect 248860 105984 251914 106040
rect 251970 105984 251975 106040
rect 248860 105982 251975 105984
rect 251909 105979 251975 105982
rect 307569 105906 307635 105909
rect 307569 105904 310132 105906
rect 307569 105848 307574 105904
rect 307630 105848 310132 105904
rect 307569 105846 310132 105848
rect 307569 105843 307635 105846
rect 214005 105634 214071 105637
rect 252461 105634 252527 105637
rect 214005 105632 217212 105634
rect 214005 105576 214010 105632
rect 214066 105576 217212 105632
rect 214005 105574 217212 105576
rect 248860 105632 252527 105634
rect 248860 105576 252466 105632
rect 252522 105576 252527 105632
rect 248860 105574 252527 105576
rect 214005 105571 214071 105574
rect 252461 105571 252527 105574
rect 397453 105634 397519 105637
rect 397453 105632 400108 105634
rect 397453 105576 397458 105632
rect 397514 105576 400108 105632
rect 397453 105574 400108 105576
rect 397453 105571 397519 105574
rect 305913 105498 305979 105501
rect 324313 105498 324379 105501
rect 305913 105496 310132 105498
rect 305913 105440 305918 105496
rect 305974 105440 310132 105496
rect 305913 105438 310132 105440
rect 321908 105496 324379 105498
rect 321908 105440 324318 105496
rect 324374 105440 324379 105496
rect 321908 105438 324379 105440
rect 305913 105435 305979 105438
rect 324313 105435 324379 105438
rect 251357 105090 251423 105093
rect 248860 105088 251423 105090
rect 248860 105032 251362 105088
rect 251418 105032 251423 105088
rect 248860 105030 251423 105032
rect 251357 105027 251423 105030
rect 307661 105090 307727 105093
rect 307661 105088 310132 105090
rect 307661 105032 307666 105088
rect 307722 105032 310132 105088
rect 307661 105030 310132 105032
rect 307661 105027 307727 105030
rect 213913 104954 213979 104957
rect 452561 104954 452627 104957
rect 213913 104952 217212 104954
rect 213913 104896 213918 104952
rect 213974 104896 217212 104952
rect 213913 104894 217212 104896
rect 449788 104952 452627 104954
rect 449788 104896 452566 104952
rect 452622 104896 452627 104952
rect 449788 104894 452627 104896
rect 213913 104891 213979 104894
rect 452561 104891 452627 104894
rect 324497 104818 324563 104821
rect 321908 104816 324563 104818
rect 321908 104760 324502 104816
rect 324558 104760 324563 104816
rect 321908 104758 324563 104760
rect 324497 104755 324563 104758
rect 251909 104682 251975 104685
rect 248860 104680 251975 104682
rect 248860 104624 251914 104680
rect 251970 104624 251975 104680
rect 248860 104622 251975 104624
rect 251909 104619 251975 104622
rect 307477 104682 307543 104685
rect 307477 104680 310132 104682
rect 307477 104624 307482 104680
rect 307538 104624 310132 104680
rect 307477 104622 310132 104624
rect 307477 104619 307543 104622
rect 214005 104274 214071 104277
rect 307661 104274 307727 104277
rect 214005 104272 217212 104274
rect 214005 104216 214010 104272
rect 214066 104216 217212 104272
rect 214005 104214 217212 104216
rect 307661 104272 310132 104274
rect 307661 104216 307666 104272
rect 307722 104216 310132 104272
rect 307661 104214 310132 104216
rect 214005 104211 214071 104214
rect 307661 104211 307727 104214
rect 252461 104138 252527 104141
rect 248860 104136 252527 104138
rect 248860 104080 252466 104136
rect 252522 104080 252527 104136
rect 248860 104078 252527 104080
rect 252461 104075 252527 104078
rect 398005 104138 398071 104141
rect 450169 104138 450235 104141
rect 398005 104136 400108 104138
rect 398005 104080 398010 104136
rect 398066 104080 400108 104136
rect 398005 104078 400108 104080
rect 449788 104136 450235 104138
rect 449788 104080 450174 104136
rect 450230 104080 450235 104136
rect 449788 104078 450235 104080
rect 398005 104075 398071 104078
rect 450169 104075 450235 104078
rect 324313 104002 324379 104005
rect 321908 104000 324379 104002
rect 321908 103944 324318 104000
rect 324374 103944 324379 104000
rect 321908 103942 324379 103944
rect 324313 103939 324379 103942
rect 307569 103866 307635 103869
rect 307569 103864 310132 103866
rect 307569 103808 307574 103864
rect 307630 103808 310132 103864
rect 307569 103806 310132 103808
rect 307569 103803 307635 103806
rect 251725 103730 251791 103733
rect 248860 103728 251791 103730
rect 248860 103672 251730 103728
rect 251786 103672 251791 103728
rect 248860 103670 251791 103672
rect 251725 103667 251791 103670
rect 213913 103594 213979 103597
rect 397545 103594 397611 103597
rect 213913 103592 217212 103594
rect 213913 103536 213918 103592
rect 213974 103536 217212 103592
rect 213913 103534 217212 103536
rect 397545 103592 400108 103594
rect 397545 103536 397550 103592
rect 397606 103536 400108 103592
rect 397545 103534 400108 103536
rect 213913 103531 213979 103534
rect 397545 103531 397611 103534
rect 307569 103458 307635 103461
rect 307569 103456 310132 103458
rect 307569 103400 307574 103456
rect 307630 103400 310132 103456
rect 307569 103398 310132 103400
rect 307569 103395 307635 103398
rect 252001 103186 252067 103189
rect 248860 103184 252067 103186
rect 248860 103128 252006 103184
rect 252062 103128 252067 103184
rect 248860 103126 252067 103128
rect 252001 103123 252067 103126
rect 307477 103050 307543 103053
rect 307477 103048 310132 103050
rect 307477 102992 307482 103048
rect 307538 102992 310132 103048
rect 307477 102990 310132 102992
rect 307477 102987 307543 102990
rect 214005 102914 214071 102917
rect 214005 102912 217212 102914
rect 214005 102856 214010 102912
rect 214066 102856 217212 102912
rect 214005 102854 217212 102856
rect 214005 102851 214071 102854
rect 321694 102781 321754 103156
rect 397545 102914 397611 102917
rect 452561 102914 452627 102917
rect 397545 102912 400108 102914
rect 397545 102856 397550 102912
rect 397606 102856 400108 102912
rect 397545 102854 400108 102856
rect 449788 102912 452627 102914
rect 449788 102856 452566 102912
rect 452622 102856 452627 102912
rect 449788 102854 452627 102856
rect 397545 102851 397611 102854
rect 452561 102851 452627 102854
rect 252369 102778 252435 102781
rect 248860 102776 252435 102778
rect 248860 102720 252374 102776
rect 252430 102720 252435 102776
rect 248860 102718 252435 102720
rect 252369 102715 252435 102718
rect 321645 102776 321754 102781
rect 321645 102720 321650 102776
rect 321706 102720 321754 102776
rect 321645 102718 321754 102720
rect 321645 102715 321711 102718
rect 373206 102716 373212 102780
rect 373276 102778 373282 102780
rect 374637 102778 374703 102781
rect 373276 102776 374703 102778
rect 373276 102720 374642 102776
rect 374698 102720 374703 102776
rect 373276 102718 374703 102720
rect 373276 102716 373282 102718
rect 374637 102715 374703 102718
rect 307661 102506 307727 102509
rect 324313 102506 324379 102509
rect 307661 102504 310132 102506
rect 307661 102448 307666 102504
rect 307722 102448 310132 102504
rect 307661 102446 310132 102448
rect 321908 102504 324379 102506
rect 321908 102448 324318 102504
rect 324374 102448 324379 102504
rect 321908 102446 324379 102448
rect 307661 102443 307727 102446
rect 324313 102443 324379 102446
rect 66069 102370 66135 102373
rect 68142 102370 68816 102376
rect 66069 102368 68816 102370
rect 66069 102312 66074 102368
rect 66130 102316 68816 102368
rect 66130 102312 68202 102316
rect 66069 102310 68202 102312
rect 66069 102307 66135 102310
rect 213913 102234 213979 102237
rect 252461 102234 252527 102237
rect 213913 102232 217212 102234
rect 213913 102176 213918 102232
rect 213974 102176 217212 102232
rect 213913 102174 217212 102176
rect 248860 102232 252527 102234
rect 248860 102176 252466 102232
rect 252522 102176 252527 102232
rect 248860 102174 252527 102176
rect 213913 102171 213979 102174
rect 252461 102171 252527 102174
rect 307477 102098 307543 102101
rect 307477 102096 310132 102098
rect 307477 102040 307482 102096
rect 307538 102040 310132 102096
rect 307477 102038 310132 102040
rect 307477 102035 307543 102038
rect 449758 101962 449818 102068
rect 449893 101962 449959 101965
rect 449758 101960 449959 101962
rect 449758 101904 449898 101960
rect 449954 101904 449959 101960
rect 449758 101902 449959 101904
rect 449893 101899 449959 101902
rect 252277 101826 252343 101829
rect 248860 101824 252343 101826
rect 248860 101768 252282 101824
rect 252338 101768 252343 101824
rect 248860 101766 252343 101768
rect 252277 101763 252343 101766
rect 306741 101690 306807 101693
rect 306741 101688 310132 101690
rect 306741 101632 306746 101688
rect 306802 101632 310132 101688
rect 306741 101630 310132 101632
rect 306741 101627 306807 101630
rect 215017 101554 215083 101557
rect 215017 101552 217212 101554
rect 215017 101496 215022 101552
rect 215078 101496 217212 101552
rect 215017 101494 217212 101496
rect 215017 101491 215083 101494
rect 252461 101418 252527 101421
rect 248860 101416 252527 101418
rect 248860 101360 252466 101416
rect 252522 101360 252527 101416
rect 248860 101358 252527 101360
rect 252461 101355 252527 101358
rect 307569 101282 307635 101285
rect 307569 101280 310132 101282
rect 307569 101224 307574 101280
rect 307630 101224 310132 101280
rect 307569 101222 310132 101224
rect 307569 101219 307635 101222
rect 321694 101149 321754 101660
rect 397545 101554 397611 101557
rect 397545 101552 400108 101554
rect 397545 101496 397550 101552
rect 397606 101496 400108 101552
rect 397545 101494 400108 101496
rect 397545 101491 397611 101494
rect 305821 101146 305887 101149
rect 307477 101146 307543 101149
rect 305821 101144 307543 101146
rect 305821 101088 305826 101144
rect 305882 101088 307482 101144
rect 307538 101088 307543 101144
rect 305821 101086 307543 101088
rect 321694 101144 321803 101149
rect 321694 101088 321742 101144
rect 321798 101088 321803 101144
rect 321694 101086 321803 101088
rect 305821 101083 305887 101086
rect 307477 101083 307543 101086
rect 321737 101083 321803 101086
rect 213913 101010 213979 101013
rect 449390 101012 449450 101388
rect 213913 101008 217212 101010
rect 213913 100952 213918 101008
rect 213974 100952 217212 101008
rect 213913 100950 217212 100952
rect 213913 100947 213979 100950
rect 449382 100948 449388 101012
rect 449452 100948 449458 101012
rect 252001 100874 252067 100877
rect 248860 100872 252067 100874
rect 248860 100816 252006 100872
rect 252062 100816 252067 100872
rect 248860 100814 252067 100816
rect 252001 100811 252067 100814
rect 307661 100874 307727 100877
rect 324405 100874 324471 100877
rect 307661 100872 310132 100874
rect 307661 100816 307666 100872
rect 307722 100816 310132 100872
rect 307661 100814 310132 100816
rect 321908 100872 324471 100874
rect 321908 100816 324410 100872
rect 324466 100816 324471 100872
rect 321908 100814 324471 100816
rect 307661 100811 307727 100814
rect 324405 100811 324471 100814
rect 397637 100874 397703 100877
rect 397637 100872 400108 100874
rect 397637 100816 397642 100872
rect 397698 100816 400108 100872
rect 397637 100814 400108 100816
rect 397637 100811 397703 100814
rect 67265 100738 67331 100741
rect 68142 100738 68816 100744
rect 67265 100736 68816 100738
rect 67265 100680 67270 100736
rect 67326 100684 68816 100736
rect 538254 100738 538260 100740
rect 67326 100680 68202 100684
rect 67265 100678 68202 100680
rect 67265 100675 67331 100678
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 460890 100678 538260 100738
rect 252461 100466 252527 100469
rect 248860 100464 252527 100466
rect 248860 100408 252466 100464
rect 252522 100408 252527 100464
rect 248860 100406 252527 100408
rect 252461 100403 252527 100406
rect 307569 100466 307635 100469
rect 307569 100464 310132 100466
rect 307569 100408 307574 100464
rect 307630 100408 310132 100464
rect 307569 100406 310132 100408
rect 307569 100403 307635 100406
rect 214005 100330 214071 100333
rect 214005 100328 217212 100330
rect 214005 100272 214010 100328
rect 214066 100272 217212 100328
rect 214005 100270 217212 100272
rect 214005 100267 214071 100270
rect 309225 100194 309291 100197
rect 324313 100194 324379 100197
rect 452561 100194 452627 100197
rect 296670 100192 309291 100194
rect 296670 100136 309230 100192
rect 309286 100136 309291 100192
rect 296670 100134 309291 100136
rect 321908 100192 324379 100194
rect 321908 100136 324318 100192
rect 324374 100136 324379 100192
rect 321908 100134 324379 100136
rect 449788 100192 452627 100194
rect 449788 100136 452566 100192
rect 452622 100136 452627 100192
rect 449788 100134 452627 100136
rect 288198 99996 288204 100060
rect 288268 100058 288274 100060
rect 296670 100058 296730 100134
rect 309225 100131 309291 100134
rect 324313 100131 324379 100134
rect 452561 100131 452627 100134
rect 288268 99998 296730 100058
rect 308262 99998 310132 100058
rect 288268 99996 288274 99998
rect 251725 99922 251791 99925
rect 248860 99920 251791 99922
rect 248860 99864 251730 99920
rect 251786 99864 251791 99920
rect 248860 99862 251791 99864
rect 251725 99859 251791 99862
rect 304206 99724 304212 99788
rect 304276 99786 304282 99788
rect 308262 99786 308322 99998
rect 460890 99922 460950 100678
rect 538254 100676 538260 100678
rect 538324 100676 538330 100740
rect 449390 99862 460950 99922
rect 449390 99788 449450 99862
rect 304276 99726 308322 99786
rect 304276 99724 304282 99726
rect 449382 99724 449388 99788
rect 449452 99724 449458 99788
rect 213913 99650 213979 99653
rect 307661 99650 307727 99653
rect 213913 99648 217212 99650
rect 213913 99592 213918 99648
rect 213974 99592 217212 99648
rect 213913 99590 217212 99592
rect 307661 99648 310132 99650
rect 307661 99592 307666 99648
rect 307722 99592 310132 99648
rect 307661 99590 310132 99592
rect 213913 99587 213979 99590
rect 307661 99587 307727 99590
rect 252369 99514 252435 99517
rect 248860 99512 252435 99514
rect 248860 99456 252374 99512
rect 252430 99456 252435 99512
rect 248860 99454 252435 99456
rect 252369 99451 252435 99454
rect 397545 99514 397611 99517
rect 397545 99512 400108 99514
rect 397545 99456 397550 99512
rect 397606 99456 400108 99512
rect 449390 99484 449450 99724
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 397545 99454 400108 99456
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 397545 99451 397611 99454
rect 580165 99451 580231 99454
rect 324405 99378 324471 99381
rect 321908 99376 324471 99378
rect 321908 99320 324410 99376
rect 324466 99320 324471 99376
rect 583520 99364 584960 99454
rect 321908 99318 324471 99320
rect 324405 99315 324471 99318
rect 307569 99106 307635 99109
rect 307569 99104 310132 99106
rect 307569 99048 307574 99104
rect 307630 99048 310132 99104
rect 307569 99046 310132 99048
rect 307569 99043 307635 99046
rect 214005 98970 214071 98973
rect 251173 98970 251239 98973
rect 214005 98968 217212 98970
rect 214005 98912 214010 98968
rect 214066 98912 217212 98968
rect 214005 98910 217212 98912
rect 248860 98968 251239 98970
rect 248860 98912 251178 98968
rect 251234 98912 251239 98968
rect 248860 98910 251239 98912
rect 214005 98907 214071 98910
rect 251173 98907 251239 98910
rect 399109 98834 399175 98837
rect 399109 98832 400108 98834
rect 399109 98776 399114 98832
rect 399170 98776 400108 98832
rect 399109 98774 400108 98776
rect 399109 98771 399175 98774
rect 307201 98698 307267 98701
rect 307201 98696 310132 98698
rect 307201 98640 307206 98696
rect 307262 98640 310132 98696
rect 307201 98638 310132 98640
rect 307201 98635 307267 98638
rect 251817 98562 251883 98565
rect 248860 98560 251883 98562
rect 248860 98504 251822 98560
rect 251878 98504 251883 98560
rect 248860 98502 251883 98504
rect 251817 98499 251883 98502
rect 213913 98290 213979 98293
rect 307661 98290 307727 98293
rect 213913 98288 217212 98290
rect 213913 98232 213918 98288
rect 213974 98232 217212 98288
rect 213913 98230 217212 98232
rect 307661 98288 310132 98290
rect 307661 98232 307666 98288
rect 307722 98232 310132 98288
rect 307661 98230 310132 98232
rect 213913 98227 213979 98230
rect 307661 98227 307727 98230
rect 321878 98154 321938 98532
rect 332542 98154 332548 98156
rect 321878 98094 332548 98154
rect 332542 98092 332548 98094
rect 332612 98092 332618 98156
rect 452285 98154 452351 98157
rect 449788 98152 452351 98154
rect 449788 98096 452290 98152
rect 452346 98096 452351 98152
rect 449788 98094 452351 98096
rect 452285 98091 452351 98094
rect 251541 98018 251607 98021
rect 248860 98016 251607 98018
rect 248860 97960 251546 98016
rect 251602 97960 251607 98016
rect 248860 97958 251607 97960
rect 251541 97955 251607 97958
rect 306966 97820 306972 97884
rect 307036 97882 307042 97884
rect 307036 97822 310132 97882
rect 307036 97820 307042 97822
rect 213913 97610 213979 97613
rect 252185 97610 252251 97613
rect 213913 97608 217212 97610
rect 213913 97552 213918 97608
rect 213974 97552 217212 97608
rect 213913 97550 217212 97552
rect 248860 97608 252251 97610
rect 248860 97552 252190 97608
rect 252246 97552 252251 97608
rect 248860 97550 252251 97552
rect 213913 97547 213979 97550
rect 252185 97547 252251 97550
rect 307661 97474 307727 97477
rect 307661 97472 310132 97474
rect 307661 97416 307666 97472
rect 307722 97416 310132 97472
rect 307661 97414 310132 97416
rect 307661 97411 307727 97414
rect 321510 97341 321570 97852
rect 452561 97474 452627 97477
rect 449788 97472 452627 97474
rect 449788 97416 452566 97472
rect 452622 97416 452627 97472
rect 449788 97414 452627 97416
rect 452561 97411 452627 97414
rect 321461 97336 321570 97341
rect 321461 97280 321466 97336
rect 321522 97280 321570 97336
rect 321461 97278 321570 97280
rect 397545 97338 397611 97341
rect 397545 97336 400108 97338
rect 397545 97280 397550 97336
rect 397606 97280 400108 97336
rect 397545 97278 400108 97280
rect 321461 97275 321527 97278
rect 397545 97275 397611 97278
rect 251173 97066 251239 97069
rect 251909 97066 251975 97069
rect 248860 97064 251975 97066
rect 248860 97008 251178 97064
rect 251234 97008 251914 97064
rect 251970 97008 251975 97064
rect 248860 97006 251975 97008
rect 251173 97003 251239 97006
rect 251909 97003 251975 97006
rect 307569 97066 307635 97069
rect 324313 97066 324379 97069
rect 307569 97064 310132 97066
rect 307569 97008 307574 97064
rect 307630 97008 310132 97064
rect 307569 97006 310132 97008
rect 321908 97064 324379 97066
rect 321908 97008 324318 97064
rect 324374 97008 324379 97064
rect 321908 97006 324379 97008
rect 307569 97003 307635 97006
rect 324313 97003 324379 97006
rect 214557 96930 214623 96933
rect 214557 96928 217212 96930
rect 214557 96872 214562 96928
rect 214618 96872 217212 96928
rect 214557 96870 217212 96872
rect 214557 96867 214623 96870
rect 249793 96658 249859 96661
rect 252093 96658 252159 96661
rect 248860 96656 252159 96658
rect 248860 96600 249798 96656
rect 249854 96600 252098 96656
rect 252154 96600 252159 96656
rect 248860 96598 252159 96600
rect 249793 96595 249859 96598
rect 252093 96595 252159 96598
rect 307661 96658 307727 96661
rect 396901 96658 396967 96661
rect 307661 96656 310132 96658
rect 307661 96600 307666 96656
rect 307722 96600 310132 96656
rect 307661 96598 310132 96600
rect 396901 96656 400108 96658
rect 396901 96600 396906 96656
rect 396962 96600 400108 96656
rect 396901 96598 400108 96600
rect 307661 96595 307727 96598
rect 396901 96595 396967 96598
rect 213913 96386 213979 96389
rect 213913 96384 217212 96386
rect 213913 96328 213918 96384
rect 213974 96328 217212 96384
rect 213913 96326 217212 96328
rect 213913 96323 213979 96326
rect 251265 96250 251331 96253
rect 248860 96248 251331 96250
rect 248860 96192 251270 96248
rect 251326 96192 251331 96248
rect 248860 96190 251331 96192
rect 251265 96187 251331 96190
rect 307661 96250 307727 96253
rect 307661 96248 310132 96250
rect 307661 96192 307666 96248
rect 307722 96192 310132 96248
rect 307661 96190 310132 96192
rect 307661 96187 307727 96190
rect 321326 95706 321386 96356
rect 450118 96114 450124 96116
rect 449788 96054 450124 96114
rect 450118 96052 450124 96054
rect 450188 96052 450194 96116
rect 333094 95706 333100 95708
rect 315990 95646 333100 95706
rect 261334 95372 261340 95436
rect 261404 95434 261410 95436
rect 315990 95434 316050 95646
rect 333094 95644 333100 95646
rect 333164 95644 333170 95708
rect 261404 95374 316050 95434
rect 261404 95372 261410 95374
rect 442993 95298 443059 95301
rect 443821 95298 443887 95301
rect 534390 95298 534396 95300
rect 442993 95296 534396 95298
rect 442993 95240 442998 95296
rect 443054 95240 443826 95296
rect 443882 95240 534396 95296
rect 442993 95238 534396 95240
rect 442993 95235 443059 95238
rect 443821 95235 443887 95238
rect 534390 95236 534396 95238
rect 534460 95236 534466 95300
rect 175917 95162 175983 95165
rect 324262 95162 324268 95164
rect 175917 95160 324268 95162
rect 175917 95104 175922 95160
rect 175978 95104 324268 95160
rect 175917 95102 324268 95104
rect 175917 95099 175983 95102
rect 324262 95100 324268 95102
rect 324332 95100 324338 95164
rect 151721 94892 151787 94893
rect 106472 94828 106478 94892
rect 106542 94890 106548 94892
rect 106774 94890 106780 94892
rect 106542 94830 106780 94890
rect 106542 94828 106548 94830
rect 106774 94828 106780 94830
rect 106844 94828 106850 94892
rect 151721 94890 151766 94892
rect 151674 94888 151766 94890
rect 151674 94832 151726 94888
rect 151674 94830 151766 94832
rect 151721 94828 151766 94830
rect 151830 94828 151836 94892
rect 151721 94827 151787 94828
rect 94957 94756 95023 94757
rect 113173 94756 113239 94757
rect 94912 94692 94918 94756
rect 94982 94754 95023 94756
rect 94982 94752 95074 94754
rect 95018 94696 95074 94752
rect 94982 94694 95074 94696
rect 94982 94692 95023 94694
rect 113136 94692 113142 94756
rect 113206 94754 113239 94756
rect 115841 94756 115907 94757
rect 126513 94756 126579 94757
rect 115841 94754 115862 94756
rect 113206 94752 113298 94754
rect 113234 94696 113298 94752
rect 113206 94694 113298 94696
rect 115770 94752 115862 94754
rect 115770 94696 115846 94752
rect 115770 94694 115862 94696
rect 113206 94692 113239 94694
rect 94957 94691 95023 94692
rect 113173 94691 113239 94692
rect 115841 94692 115862 94694
rect 115926 94692 115932 94756
rect 126464 94692 126470 94756
rect 126534 94754 126579 94756
rect 126534 94752 126626 94754
rect 126574 94696 126626 94752
rect 126534 94694 126626 94696
rect 126534 94692 126579 94694
rect 115841 94691 115907 94692
rect 126513 94691 126579 94692
rect 128118 93876 128124 93940
rect 128188 93938 128194 93940
rect 166206 93938 166212 93940
rect 128188 93878 166212 93938
rect 128188 93876 128194 93878
rect 166206 93876 166212 93878
rect 166276 93876 166282 93940
rect 171726 93740 171732 93804
rect 171796 93802 171802 93804
rect 324497 93802 324563 93805
rect 171796 93800 324563 93802
rect 171796 93744 324502 93800
rect 324558 93744 324563 93800
rect 171796 93742 324563 93744
rect 171796 93740 171802 93742
rect 324497 93739 324563 93742
rect 430389 93802 430455 93805
rect 453297 93802 453363 93805
rect 430389 93800 453363 93802
rect 430389 93744 430394 93800
rect 430450 93744 453302 93800
rect 453358 93744 453363 93800
rect 430389 93742 453363 93744
rect 430389 93739 430455 93742
rect 453297 93739 453363 93742
rect 130745 93668 130811 93669
rect 130694 93666 130700 93668
rect 130654 93606 130700 93666
rect 130764 93664 130811 93668
rect 130806 93608 130811 93664
rect 130694 93604 130700 93606
rect 130764 93604 130811 93608
rect 173566 93604 173572 93668
rect 173636 93666 173642 93668
rect 324405 93666 324471 93669
rect 173636 93664 324471 93666
rect 173636 93608 324410 93664
rect 324466 93608 324471 93664
rect 173636 93606 324471 93608
rect 173636 93604 173642 93606
rect 130745 93603 130811 93604
rect 324405 93603 324471 93606
rect 97257 93532 97323 93533
rect 113817 93532 113883 93533
rect 97206 93530 97212 93532
rect 97166 93470 97212 93530
rect 97276 93528 97323 93532
rect 113766 93530 113772 93532
rect 97318 93472 97323 93528
rect 97206 93468 97212 93470
rect 97276 93468 97323 93472
rect 113726 93470 113772 93530
rect 113836 93528 113883 93532
rect 113878 93472 113883 93528
rect 113766 93468 113772 93470
rect 113836 93468 113883 93472
rect 97257 93467 97323 93468
rect 113817 93467 113883 93468
rect 110137 93260 110203 93261
rect 110086 93258 110092 93260
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 110137 93195 110203 93196
rect 87137 92444 87203 92445
rect 98177 92444 98243 92445
rect 87086 92442 87092 92444
rect 87046 92382 87092 92442
rect 87156 92440 87203 92444
rect 98126 92442 98132 92444
rect 87198 92384 87203 92440
rect 87086 92380 87092 92382
rect 87156 92380 87203 92384
rect 98086 92382 98132 92442
rect 98196 92440 98243 92444
rect 98238 92384 98243 92440
rect 98126 92380 98132 92382
rect 98196 92380 98243 92384
rect 98494 92380 98500 92444
rect 98564 92442 98570 92444
rect 98637 92442 98703 92445
rect 98564 92440 98703 92442
rect 98564 92384 98642 92440
rect 98698 92384 98703 92440
rect 98564 92382 98703 92384
rect 98564 92380 98570 92382
rect 87137 92379 87203 92380
rect 98177 92379 98243 92380
rect 98637 92379 98703 92382
rect 106774 92380 106780 92444
rect 106844 92442 106850 92444
rect 107377 92442 107443 92445
rect 116761 92444 116827 92445
rect 116710 92442 116716 92444
rect 106844 92440 107443 92442
rect 106844 92384 107382 92440
rect 107438 92384 107443 92440
rect 106844 92382 107443 92384
rect 116670 92382 116716 92442
rect 116780 92440 116827 92444
rect 116822 92384 116827 92440
rect 106844 92380 106850 92382
rect 107377 92379 107443 92382
rect 116710 92380 116716 92382
rect 116780 92380 116827 92384
rect 120206 92380 120212 92444
rect 120276 92442 120282 92444
rect 120349 92442 120415 92445
rect 120276 92440 120415 92442
rect 120276 92384 120354 92440
rect 120410 92384 120415 92440
rect 120276 92382 120415 92384
rect 120276 92380 120282 92382
rect 116761 92379 116827 92380
rect 120349 92379 120415 92382
rect 124029 92444 124095 92445
rect 125777 92444 125843 92445
rect 129457 92444 129523 92445
rect 133137 92444 133203 92445
rect 135713 92444 135779 92445
rect 151537 92444 151603 92445
rect 152089 92444 152155 92445
rect 124029 92440 124076 92444
rect 124140 92442 124146 92444
rect 125726 92442 125732 92444
rect 124029 92384 124034 92440
rect 124029 92380 124076 92384
rect 124140 92382 124186 92442
rect 125686 92382 125732 92442
rect 125796 92440 125843 92444
rect 129406 92442 129412 92444
rect 125838 92384 125843 92440
rect 124140 92380 124146 92382
rect 125726 92380 125732 92382
rect 125796 92380 125843 92384
rect 129366 92382 129412 92442
rect 129476 92440 129523 92444
rect 133086 92442 133092 92444
rect 129518 92384 129523 92440
rect 129406 92380 129412 92382
rect 129476 92380 129523 92384
rect 133046 92382 133092 92442
rect 133156 92440 133203 92444
rect 135662 92442 135668 92444
rect 133198 92384 133203 92440
rect 133086 92380 133092 92382
rect 133156 92380 133203 92384
rect 135622 92382 135668 92442
rect 135732 92440 135779 92444
rect 151486 92442 151492 92444
rect 135774 92384 135779 92440
rect 135662 92380 135668 92382
rect 135732 92380 135779 92384
rect 151446 92382 151492 92442
rect 151556 92440 151603 92444
rect 152038 92442 152044 92444
rect 151598 92384 151603 92440
rect 151486 92380 151492 92382
rect 151556 92380 151603 92384
rect 151998 92382 152044 92442
rect 152108 92440 152155 92444
rect 152150 92384 152155 92440
rect 152038 92380 152044 92382
rect 152108 92380 152155 92384
rect 170254 92380 170260 92444
rect 170324 92442 170330 92444
rect 324313 92442 324379 92445
rect 170324 92440 324379 92442
rect 170324 92384 324318 92440
rect 324374 92384 324379 92440
rect 170324 92382 324379 92384
rect 170324 92380 170330 92382
rect 124029 92379 124095 92380
rect 125777 92379 125843 92380
rect 129457 92379 129523 92380
rect 133137 92379 133203 92380
rect 135713 92379 135779 92380
rect 151537 92379 151603 92380
rect 152089 92379 152155 92380
rect 324313 92379 324379 92382
rect 114134 92244 114140 92308
rect 114204 92306 114210 92308
rect 207749 92306 207815 92309
rect 114204 92304 207815 92306
rect 114204 92248 207754 92304
rect 207810 92248 207815 92304
rect 114204 92246 207815 92248
rect 114204 92244 114210 92246
rect 207749 92243 207815 92246
rect 119654 92108 119660 92172
rect 119724 92170 119730 92172
rect 167678 92170 167684 92172
rect 119724 92110 167684 92170
rect 119724 92108 119730 92110
rect 167678 92108 167684 92110
rect 167748 92108 167754 92172
rect 99598 91700 99604 91764
rect 99668 91762 99674 91764
rect 99741 91762 99807 91765
rect 117129 91764 117195 91765
rect 117078 91762 117084 91764
rect 99668 91760 99807 91762
rect 99668 91704 99746 91760
rect 99802 91704 99807 91760
rect 99668 91702 99807 91704
rect 117038 91702 117084 91762
rect 117148 91760 117195 91764
rect 117190 91704 117195 91760
rect 99668 91700 99674 91702
rect 99741 91699 99807 91702
rect 117078 91700 117084 91702
rect 117148 91700 117195 91704
rect 305494 91700 305500 91764
rect 305564 91762 305570 91764
rect 316033 91762 316099 91765
rect 305564 91760 316099 91762
rect 305564 91704 316038 91760
rect 316094 91704 316099 91760
rect 305564 91702 316099 91704
rect 305564 91700 305570 91702
rect 117129 91699 117195 91700
rect 316033 91699 316099 91702
rect 109166 91564 109172 91628
rect 109236 91626 109242 91628
rect 110321 91626 110387 91629
rect 109236 91624 110387 91626
rect 109236 91568 110326 91624
rect 110382 91568 110387 91624
rect 109236 91566 110387 91568
rect 109236 91564 109242 91566
rect 110321 91563 110387 91566
rect 131982 91564 131988 91628
rect 132052 91626 132058 91628
rect 132217 91626 132283 91629
rect 151353 91628 151419 91629
rect 151302 91626 151308 91628
rect 132052 91624 132283 91626
rect 132052 91568 132222 91624
rect 132278 91568 132283 91624
rect 132052 91566 132283 91568
rect 151262 91566 151308 91626
rect 151372 91624 151419 91628
rect 151414 91568 151419 91624
rect 132052 91564 132058 91566
rect 132217 91563 132283 91566
rect 151302 91564 151308 91566
rect 151372 91564 151419 91568
rect 151353 91563 151419 91564
rect 122833 91492 122899 91493
rect 122782 91428 122788 91492
rect 122852 91490 122899 91492
rect 122852 91488 122944 91490
rect 122894 91432 122944 91488
rect 122852 91430 122944 91432
rect 122852 91428 122899 91430
rect 122833 91427 122899 91428
rect 101806 91292 101812 91356
rect 101876 91354 101882 91356
rect 101949 91354 102015 91357
rect 101876 91352 102015 91354
rect 101876 91296 101954 91352
rect 102010 91296 102015 91352
rect 101876 91294 102015 91296
rect 101876 91292 101882 91294
rect 101949 91291 102015 91294
rect 104198 91292 104204 91356
rect 104268 91354 104274 91356
rect 104801 91354 104867 91357
rect 104268 91352 104867 91354
rect 104268 91296 104806 91352
rect 104862 91296 104867 91352
rect 104268 91294 104867 91296
rect 104268 91292 104274 91294
rect 104801 91291 104867 91294
rect 107694 91292 107700 91356
rect 107764 91354 107770 91356
rect 108941 91354 109007 91357
rect 107764 91352 109007 91354
rect 107764 91296 108946 91352
rect 109002 91296 109007 91352
rect 107764 91294 109007 91296
rect 107764 91292 107770 91294
rect 108941 91291 109007 91294
rect 112294 91292 112300 91356
rect 112364 91354 112370 91356
rect 112437 91354 112503 91357
rect 112364 91352 112503 91354
rect 112364 91296 112442 91352
rect 112498 91296 112503 91352
rect 112364 91294 112503 91296
rect 112364 91292 112370 91294
rect 112437 91291 112503 91294
rect 124438 91292 124444 91356
rect 124508 91354 124514 91356
rect 125409 91354 125475 91357
rect 124508 91352 125475 91354
rect 124508 91296 125414 91352
rect 125470 91296 125475 91352
rect 124508 91294 125475 91296
rect 124508 91292 124514 91294
rect 125409 91291 125475 91294
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75361 91218 75427 91221
rect 74828 91216 75427 91218
rect 74828 91160 75366 91216
rect 75422 91160 75427 91216
rect 74828 91158 75427 91160
rect 74828 91156 74834 91158
rect 75361 91155 75427 91158
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85481 91218 85547 91221
rect 84396 91216 85547 91218
rect 84396 91160 85486 91216
rect 85542 91160 85547 91216
rect 84396 91158 85547 91160
rect 84396 91156 84402 91158
rect 85481 91155 85547 91158
rect 85614 91156 85620 91220
rect 85684 91218 85690 91220
rect 86401 91218 86467 91221
rect 85684 91216 86467 91218
rect 85684 91160 86406 91216
rect 86462 91160 86467 91216
rect 85684 91158 86467 91160
rect 85684 91156 85690 91158
rect 86401 91155 86467 91158
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 86788 91156 86794 91158
rect 86861 91155 86927 91158
rect 88926 91156 88932 91220
rect 88996 91218 89002 91220
rect 89621 91218 89687 91221
rect 88996 91216 89687 91218
rect 88996 91160 89626 91216
rect 89682 91160 89687 91216
rect 88996 91158 89687 91160
rect 88996 91156 89002 91158
rect 89621 91155 89687 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 90633 91218 90699 91221
rect 90284 91216 90699 91218
rect 90284 91160 90638 91216
rect 90694 91160 90699 91216
rect 90284 91158 90699 91160
rect 90284 91156 90290 91158
rect 90633 91155 90699 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92381 91218 92447 91221
rect 91388 91216 92447 91218
rect 91388 91160 92386 91216
rect 92442 91160 92447 91216
rect 91388 91158 92447 91160
rect 91388 91156 91394 91158
rect 92381 91155 92447 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 93894 91156 93900 91220
rect 93964 91218 93970 91220
rect 95141 91218 95207 91221
rect 93964 91216 95207 91218
rect 93964 91160 95146 91216
rect 95202 91160 95207 91216
rect 93964 91158 95207 91160
rect 93964 91156 93970 91158
rect 95141 91155 95207 91158
rect 96102 91156 96108 91220
rect 96172 91218 96178 91220
rect 96521 91218 96587 91221
rect 96172 91216 96587 91218
rect 96172 91160 96526 91216
rect 96582 91160 96587 91216
rect 96172 91158 96587 91160
rect 96172 91156 96178 91158
rect 96521 91155 96587 91158
rect 97022 91156 97028 91220
rect 97092 91218 97098 91220
rect 97901 91218 97967 91221
rect 99281 91220 99347 91221
rect 99230 91218 99236 91220
rect 97092 91216 97967 91218
rect 97092 91160 97906 91216
rect 97962 91160 97967 91216
rect 97092 91158 97967 91160
rect 99190 91158 99236 91218
rect 99300 91216 99347 91220
rect 99342 91160 99347 91216
rect 97092 91156 97098 91158
rect 97901 91155 97967 91158
rect 99230 91156 99236 91158
rect 99300 91156 99347 91160
rect 100518 91156 100524 91220
rect 100588 91218 100594 91220
rect 100661 91218 100727 91221
rect 101673 91220 101739 91221
rect 102041 91220 102107 91221
rect 102961 91220 103027 91221
rect 103329 91220 103395 91221
rect 101622 91218 101628 91220
rect 100588 91216 100727 91218
rect 100588 91160 100666 91216
rect 100722 91160 100727 91216
rect 100588 91158 100727 91160
rect 101582 91158 101628 91218
rect 101692 91216 101739 91220
rect 101990 91218 101996 91220
rect 101734 91160 101739 91216
rect 100588 91156 100594 91158
rect 99281 91155 99347 91156
rect 100661 91155 100727 91158
rect 101622 91156 101628 91158
rect 101692 91156 101739 91160
rect 101950 91158 101996 91218
rect 102060 91216 102107 91220
rect 102910 91218 102916 91220
rect 102102 91160 102107 91216
rect 101990 91156 101996 91158
rect 102060 91156 102107 91160
rect 102870 91158 102916 91218
rect 102980 91216 103027 91220
rect 103278 91218 103284 91220
rect 103022 91160 103027 91216
rect 102910 91156 102916 91158
rect 102980 91156 103027 91160
rect 103238 91158 103284 91218
rect 103348 91216 103395 91220
rect 103390 91160 103395 91216
rect 103278 91156 103284 91158
rect 103348 91156 103395 91160
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104709 91218 104775 91221
rect 104636 91216 104775 91218
rect 104636 91160 104714 91216
rect 104770 91160 104775 91216
rect 104636 91158 104775 91160
rect 104636 91156 104642 91158
rect 101673 91155 101739 91156
rect 102041 91155 102107 91156
rect 102961 91155 103027 91156
rect 103329 91155 103395 91156
rect 104709 91155 104775 91158
rect 105118 91156 105124 91220
rect 105188 91218 105194 91220
rect 105721 91218 105787 91221
rect 105188 91216 105787 91218
rect 105188 91160 105726 91216
rect 105782 91160 105787 91216
rect 105188 91158 105787 91160
rect 105188 91156 105194 91158
rect 105721 91155 105787 91158
rect 106038 91156 106044 91220
rect 106108 91156 106114 91220
rect 106406 91156 106412 91220
rect 106476 91218 106482 91220
rect 107469 91218 107535 91221
rect 106476 91216 107535 91218
rect 106476 91160 107474 91216
rect 107530 91160 107535 91216
rect 106476 91158 107535 91160
rect 106476 91156 106482 91158
rect 106046 91082 106106 91156
rect 107469 91155 107535 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108849 91218 108915 91221
rect 108132 91216 108915 91218
rect 108132 91160 108854 91216
rect 108910 91160 108915 91216
rect 108132 91158 108915 91160
rect 108132 91156 108138 91158
rect 108849 91155 108915 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 109769 91218 109835 91221
rect 109604 91216 109835 91218
rect 109604 91160 109774 91216
rect 109830 91160 109835 91216
rect 109604 91158 109835 91160
rect 109604 91156 109610 91158
rect 109769 91155 109835 91158
rect 110638 91156 110644 91220
rect 110708 91218 110714 91220
rect 111057 91218 111123 91221
rect 110708 91216 111123 91218
rect 110708 91160 111062 91216
rect 111118 91160 111123 91216
rect 110708 91158 111123 91160
rect 110708 91156 110714 91158
rect 111057 91155 111123 91158
rect 111190 91156 111196 91220
rect 111260 91218 111266 91220
rect 111701 91218 111767 91221
rect 111260 91216 111767 91218
rect 111260 91160 111706 91216
rect 111762 91160 111767 91216
rect 111260 91158 111767 91160
rect 111260 91156 111266 91158
rect 111701 91155 111767 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 113081 91218 113147 91221
rect 111996 91216 113147 91218
rect 111996 91160 113086 91216
rect 113142 91160 113147 91216
rect 111996 91158 113147 91160
rect 111996 91156 112002 91158
rect 113081 91155 113147 91158
rect 115054 91156 115060 91220
rect 115124 91218 115130 91220
rect 115289 91218 115355 91221
rect 115124 91216 115355 91218
rect 115124 91160 115294 91216
rect 115350 91160 115355 91216
rect 115124 91158 115355 91160
rect 115124 91156 115130 91158
rect 115289 91155 115355 91158
rect 115422 91156 115428 91220
rect 115492 91218 115498 91220
rect 115841 91218 115907 91221
rect 118049 91220 118115 91221
rect 117998 91218 118004 91220
rect 115492 91216 115907 91218
rect 115492 91160 115846 91216
rect 115902 91160 115907 91216
rect 115492 91158 115907 91160
rect 117958 91158 118004 91218
rect 118068 91216 118115 91220
rect 118110 91160 118115 91216
rect 115492 91156 115498 91158
rect 115841 91155 115907 91158
rect 117998 91156 118004 91158
rect 118068 91156 118115 91160
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118601 91218 118667 91221
rect 119889 91220 119955 91221
rect 119838 91218 119844 91220
rect 118252 91216 118667 91218
rect 118252 91160 118606 91216
rect 118662 91160 118667 91216
rect 118252 91158 118667 91160
rect 119798 91158 119844 91218
rect 119908 91216 119955 91220
rect 119950 91160 119955 91216
rect 118252 91156 118258 91158
rect 118049 91155 118115 91156
rect 118601 91155 118667 91158
rect 119838 91156 119844 91158
rect 119908 91156 119955 91160
rect 120574 91156 120580 91220
rect 120644 91218 120650 91220
rect 121361 91218 121427 91221
rect 120644 91216 121427 91218
rect 120644 91160 121366 91216
rect 121422 91160 121427 91216
rect 120644 91158 121427 91160
rect 120644 91156 120650 91158
rect 119889 91155 119955 91156
rect 121361 91155 121427 91158
rect 121678 91156 121684 91220
rect 121748 91218 121754 91220
rect 121913 91218 121979 91221
rect 121748 91216 121979 91218
rect 121748 91160 121918 91216
rect 121974 91160 121979 91216
rect 121748 91158 121979 91160
rect 121748 91156 121754 91158
rect 121913 91155 121979 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122741 91218 122807 91221
rect 122116 91216 122807 91218
rect 122116 91160 122746 91216
rect 122802 91160 122807 91216
rect 122116 91158 122807 91160
rect 122116 91156 122122 91158
rect 122741 91155 122807 91158
rect 122966 91156 122972 91220
rect 123036 91218 123042 91220
rect 124121 91218 124187 91221
rect 123036 91216 124187 91218
rect 123036 91160 124126 91216
rect 124182 91160 124187 91216
rect 123036 91158 124187 91160
rect 123036 91156 123042 91158
rect 124121 91155 124187 91158
rect 125358 91156 125364 91220
rect 125428 91218 125434 91220
rect 125501 91218 125567 91221
rect 125428 91216 125567 91218
rect 125428 91160 125506 91216
rect 125562 91160 125567 91216
rect 125428 91158 125567 91160
rect 125428 91156 125434 91158
rect 125501 91155 125567 91158
rect 126646 91156 126652 91220
rect 126716 91218 126722 91220
rect 126881 91218 126947 91221
rect 126716 91216 126947 91218
rect 126716 91160 126886 91216
rect 126942 91160 126947 91216
rect 126716 91158 126947 91160
rect 126716 91156 126722 91158
rect 126881 91155 126947 91158
rect 134374 91156 134380 91220
rect 134444 91218 134450 91220
rect 134793 91218 134859 91221
rect 134444 91216 134859 91218
rect 134444 91160 134798 91216
rect 134854 91160 134859 91216
rect 134444 91158 134859 91160
rect 134444 91156 134450 91158
rect 134793 91155 134859 91158
rect 166390 91082 166396 91084
rect 106046 91022 166396 91082
rect 166390 91020 166396 91022
rect 166460 91020 166466 91084
rect 380566 91020 380572 91084
rect 380636 91082 380642 91084
rect 427721 91082 427787 91085
rect 380636 91080 427787 91082
rect 380636 91024 427726 91080
rect 427782 91024 427787 91080
rect 380636 91022 427787 91024
rect 380636 91020 380642 91022
rect 427721 91019 427787 91022
rect 67357 89722 67423 89725
rect 215017 89722 215083 89725
rect 67357 89720 215083 89722
rect 67357 89664 67362 89720
rect 67418 89664 215022 89720
rect 215078 89664 215083 89720
rect 67357 89662 215083 89664
rect 67357 89659 67423 89662
rect 215017 89659 215083 89662
rect 214557 89042 214623 89045
rect 307150 89042 307156 89044
rect 214557 89040 307156 89042
rect 214557 88984 214562 89040
rect 214618 88984 307156 89040
rect 214557 88982 307156 88984
rect 214557 88979 214623 88982
rect 307150 88980 307156 88982
rect 307220 88980 307226 89044
rect 109769 88226 109835 88229
rect 170397 88226 170463 88229
rect 109769 88224 170463 88226
rect 109769 88168 109774 88224
rect 109830 88168 170402 88224
rect 170458 88168 170463 88224
rect 109769 88166 170463 88168
rect 109769 88163 109835 88166
rect 170397 88163 170463 88166
rect 179086 86124 179092 86188
rect 179156 86186 179162 86188
rect 245653 86186 245719 86189
rect 179156 86184 245719 86186
rect 179156 86128 245658 86184
rect 245714 86128 245719 86184
rect 179156 86126 245719 86128
rect 179156 86124 179162 86126
rect 245653 86123 245719 86126
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 101673 85506 101739 85509
rect 169150 85506 169156 85508
rect 101673 85504 169156 85506
rect 101673 85448 101678 85504
rect 101734 85448 169156 85504
rect 101673 85446 169156 85448
rect 101673 85443 101739 85446
rect 169150 85444 169156 85446
rect 169220 85444 169226 85508
rect -960 84690 480 84780
rect 176326 84764 176332 84828
rect 176396 84826 176402 84828
rect 313733 84826 313799 84829
rect 176396 84824 313799 84826
rect 176396 84768 313738 84824
rect 313794 84768 313799 84824
rect 176396 84766 313799 84768
rect 176396 84764 176402 84766
rect 313733 84763 313799 84766
rect 332041 84826 332107 84829
rect 449382 84826 449388 84828
rect 332041 84824 449388 84826
rect 332041 84768 332046 84824
rect 332102 84768 449388 84824
rect 332041 84766 449388 84768
rect 332041 84763 332107 84766
rect 449382 84764 449388 84766
rect 449452 84764 449458 84828
rect 2773 84690 2839 84693
rect -960 84688 2839 84690
rect -960 84632 2778 84688
rect 2834 84632 2839 84688
rect -960 84630 2839 84632
rect -960 84540 480 84630
rect 2773 84627 2839 84630
rect 295333 84284 295399 84285
rect 295333 84282 295380 84284
rect 295288 84280 295380 84282
rect 295288 84224 295338 84280
rect 295288 84222 295380 84224
rect 295333 84220 295380 84222
rect 295444 84220 295450 84284
rect 295333 84219 295399 84220
rect 102041 80066 102107 80069
rect 167494 80066 167500 80068
rect 102041 80064 167500 80066
rect 102041 80008 102046 80064
rect 102102 80008 167500 80064
rect 102041 80006 167500 80008
rect 102041 80003 102107 80006
rect 167494 80004 167500 80006
rect 167564 80004 167570 80068
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 16573 72450 16639 72453
rect 304206 72450 304212 72452
rect 16573 72448 304212 72450
rect 16573 72392 16578 72448
rect 16634 72392 304212 72448
rect 16573 72390 304212 72392
rect 16573 72387 16639 72390
rect 304206 72388 304212 72390
rect 304276 72388 304282 72452
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 31753 68234 31819 68237
rect 301630 68234 301636 68236
rect 31753 68232 301636 68234
rect 31753 68176 31758 68232
rect 31814 68176 301636 68232
rect 31753 68174 301636 68176
rect 31753 68171 31819 68174
rect 301630 68172 301636 68174
rect 301700 68172 301706 68236
rect 177062 65452 177068 65516
rect 177132 65514 177138 65516
rect 333237 65514 333303 65517
rect 177132 65512 333303 65514
rect 177132 65456 333242 65512
rect 333298 65456 333303 65512
rect 177132 65454 333303 65456
rect 177132 65452 177138 65454
rect 333237 65451 333303 65454
rect 269113 60076 269179 60077
rect 269062 60012 269068 60076
rect 269132 60074 269179 60076
rect 269132 60072 269224 60074
rect 269174 60016 269224 60072
rect 269132 60014 269224 60016
rect 269132 60012 269179 60014
rect 269113 60011 269179 60012
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 271086 46820 271092 46884
rect 271156 46882 271162 46884
rect 271689 46882 271755 46885
rect 271156 46880 271755 46882
rect 271156 46824 271694 46880
rect 271750 46824 271755 46880
rect 271156 46822 271755 46824
rect 271156 46820 271162 46822
rect 271689 46819 271755 46822
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 333237 45522 333303 45525
rect 448462 45522 448468 45524
rect 333237 45520 448468 45522
rect 333237 45464 333242 45520
rect 333298 45464 448468 45520
rect 333237 45462 448468 45464
rect 333237 45459 333303 45462
rect 448462 45460 448468 45462
rect 448532 45460 448538 45524
rect 332685 44298 332751 44301
rect 333237 44298 333303 44301
rect 332685 44296 333303 44298
rect 332685 44240 332690 44296
rect 332746 44240 333242 44296
rect 333298 44240 333303 44296
rect 332685 44238 333303 44240
rect 332685 44235 332751 44238
rect 333237 44235 333303 44238
rect 340086 42740 340092 42804
rect 340156 42802 340162 42804
rect 451038 42802 451044 42804
rect 340156 42742 451044 42802
rect 340156 42740 340162 42742
rect 451038 42740 451044 42742
rect 451108 42740 451114 42804
rect 307753 42122 307819 42125
rect 340086 42122 340092 42124
rect 307753 42120 340092 42122
rect 307753 42064 307758 42120
rect 307814 42064 340092 42120
rect 307753 42062 340092 42064
rect 307753 42059 307819 42062
rect 340086 42060 340092 42062
rect 340156 42060 340162 42124
rect 579889 33146 579955 33149
rect 583520 33146 584960 33236
rect 579889 33144 584960 33146
rect 579889 33088 579894 33144
rect 579950 33088 584960 33144
rect 579889 33086 584960 33088
rect 579889 33083 579955 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 179822 32404 179828 32468
rect 179892 32466 179898 32468
rect 287973 32466 288039 32469
rect 179892 32464 288039 32466
rect 179892 32408 287978 32464
rect 288034 32408 288039 32464
rect 179892 32406 288039 32408
rect 179892 32404 179898 32406
rect 287973 32403 288039 32406
rect 17953 29610 18019 29613
rect 305678 29610 305684 29612
rect 17953 29608 305684 29610
rect 17953 29552 17958 29608
rect 18014 29552 305684 29608
rect 17953 29550 305684 29552
rect 17953 29547 18019 29550
rect 305678 29548 305684 29550
rect 305748 29548 305754 29612
rect 340137 28930 340203 28933
rect 342897 28930 342963 28933
rect 340137 28928 342963 28930
rect 340137 28872 340142 28928
rect 340198 28872 342902 28928
rect 342958 28872 342963 28928
rect 340137 28870 342963 28872
rect 340137 28867 340203 28870
rect 342897 28867 342963 28870
rect 176510 28188 176516 28252
rect 176580 28250 176586 28252
rect 340137 28250 340203 28253
rect 176580 28248 340203 28250
rect 176580 28192 340142 28248
rect 340198 28192 340203 28248
rect 176580 28190 340203 28192
rect 176580 28188 176586 28190
rect 340137 28187 340203 28190
rect 336825 26212 336891 26213
rect 336774 26210 336780 26212
rect 336734 26150 336780 26210
rect 336844 26208 336891 26212
rect 336886 26152 336891 26208
rect 336774 26148 336780 26150
rect 336844 26148 336891 26152
rect 336825 26147 336891 26148
rect 302233 25530 302299 25533
rect 336825 25530 336891 25533
rect 302233 25528 336891 25530
rect 302233 25472 302238 25528
rect 302294 25472 336830 25528
rect 336886 25472 336891 25528
rect 302233 25470 336891 25472
rect 302233 25467 302299 25470
rect 336825 25467 336891 25470
rect 8293 24170 8359 24173
rect 299974 24170 299980 24172
rect 8293 24168 299980 24170
rect 8293 24112 8298 24168
rect 8354 24112 299980 24168
rect 8293 24110 299980 24112
rect 8293 24107 8359 24110
rect 299974 24108 299980 24110
rect 300044 24108 300050 24172
rect 297357 22674 297423 22677
rect 449934 22674 449940 22676
rect 297357 22672 449940 22674
rect 297357 22616 297362 22672
rect 297418 22616 449940 22672
rect 297357 22614 449940 22616
rect 297357 22611 297423 22614
rect 449934 22612 449940 22614
rect 450004 22612 450010 22676
rect 175038 21932 175044 21996
rect 175108 21994 175114 21996
rect 262121 21994 262187 21997
rect 175108 21992 262187 21994
rect 175108 21936 262126 21992
rect 262182 21936 262187 21992
rect 175108 21934 262187 21936
rect 175108 21932 175114 21934
rect 262121 21931 262187 21934
rect 579889 19818 579955 19821
rect 583520 19818 584960 19908
rect 579889 19816 584960 19818
rect 579889 19760 579894 19816
rect 579950 19760 584960 19816
rect 579889 19758 584960 19760
rect 579889 19755 579955 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 289486 19212 289492 19276
rect 289556 19274 289562 19276
rect 289721 19274 289787 19277
rect 289556 19272 289787 19274
rect 289556 19216 289726 19272
rect 289782 19216 289787 19272
rect 289556 19214 289787 19216
rect 289556 19212 289562 19214
rect 289721 19211 289787 19214
rect 179270 15132 179276 15196
rect 179340 15194 179346 15196
rect 240133 15194 240199 15197
rect 240777 15194 240843 15197
rect 179340 15192 240843 15194
rect 179340 15136 240138 15192
rect 240194 15136 240782 15192
rect 240838 15136 240843 15192
rect 179340 15134 240843 15136
rect 179340 15132 179346 15134
rect 240133 15131 240199 15134
rect 240777 15131 240843 15134
rect 64638 12956 64644 13020
rect 64708 13018 64714 13020
rect 135253 13018 135319 13021
rect 64708 13016 135319 13018
rect 64708 12960 135258 13016
rect 135314 12960 135319 13016
rect 64708 12958 135319 12960
rect 64708 12956 64714 12958
rect 135253 12955 135319 12958
rect 269062 11732 269068 11796
rect 269132 11794 269138 11796
rect 270401 11794 270467 11797
rect 269132 11792 270467 11794
rect 269132 11736 270406 11792
rect 270462 11736 270467 11792
rect 269132 11734 270467 11736
rect 269132 11732 269138 11734
rect 270401 11731 270467 11734
rect 297214 11732 297220 11796
rect 297284 11794 297290 11796
rect 299565 11794 299631 11797
rect 297284 11792 299631 11794
rect 297284 11736 299570 11792
rect 299626 11736 299631 11792
rect 297284 11734 299631 11736
rect 297284 11732 297290 11734
rect 299565 11731 299631 11734
rect 9673 10298 9739 10301
rect 301446 10298 301452 10300
rect 9673 10296 301452 10298
rect 9673 10240 9678 10296
rect 9734 10240 301452 10296
rect 9673 10238 301452 10240
rect 9673 10235 9739 10238
rect 301446 10236 301452 10238
rect 301516 10236 301522 10300
rect 174854 8196 174860 8260
rect 174924 8258 174930 8260
rect 297357 8258 297423 8261
rect 174924 8256 297423 8258
rect 174924 8200 297362 8256
rect 297418 8200 297423 8256
rect 174924 8198 297423 8200
rect 174924 8196 174930 8198
rect 297357 8195 297423 8198
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3509 6490 3575 6493
rect -960 6488 3575 6490
rect -960 6432 3514 6488
rect 3570 6432 3575 6488
rect 583520 6476 584960 6566
rect -960 6430 3575 6432
rect -960 6340 480 6430
rect 3509 6427 3575 6430
rect 179454 5476 179460 5540
rect 179524 5538 179530 5540
rect 305637 5538 305703 5541
rect 179524 5536 305703 5538
rect 179524 5480 305642 5536
rect 305698 5480 305703 5536
rect 179524 5478 305703 5480
rect 179524 5476 179530 5478
rect 305637 5475 305703 5478
rect 251214 3436 251220 3500
rect 251284 3498 251290 3500
rect 252369 3498 252435 3501
rect 251284 3496 252435 3498
rect 251284 3440 252374 3496
rect 252430 3440 252435 3496
rect 251284 3438 252435 3440
rect 251284 3436 251290 3438
rect 252369 3435 252435 3438
rect 258257 3498 258323 3501
rect 265566 3498 265572 3500
rect 258257 3496 265572 3498
rect 258257 3440 258262 3496
rect 258318 3440 265572 3496
rect 258257 3438 265572 3440
rect 258257 3435 258323 3438
rect 265566 3436 265572 3438
rect 265636 3436 265642 3500
rect 125869 3362 125935 3365
rect 169702 3362 169708 3364
rect 125869 3360 169708 3362
rect 125869 3304 125874 3360
rect 125930 3304 169708 3360
rect 125869 3302 169708 3304
rect 125869 3299 125935 3302
rect 169702 3300 169708 3302
rect 169772 3300 169778 3364
rect 16297 2682 16363 2685
rect 306966 2682 306972 2684
rect 16297 2680 306972 2682
rect 16297 2624 16302 2680
rect 16358 2624 306972 2680
rect 16297 2622 306972 2624
rect 16297 2619 16363 2622
rect 306966 2620 306972 2622
rect 307036 2620 307042 2684
<< obsm3 >>
rect 68800 171594 164756 174600
rect 68800 171534 164694 171594
rect 68800 129304 164756 171534
rect 68816 129244 164756 129304
rect 68800 128080 164756 129244
rect 68816 128020 164756 128080
rect 68800 126312 164756 128020
rect 68816 126252 164756 126312
rect 68800 125224 164756 126252
rect 68816 125164 164756 125224
rect 68800 123592 164756 125164
rect 68816 123532 164756 123592
rect 68800 122640 164756 123532
rect 68816 122580 164756 122640
rect 68800 120872 164756 122580
rect 68816 120812 164756 120872
rect 68800 111754 164756 120812
rect 68800 111694 164694 111754
rect 68800 110122 164756 111694
rect 68800 110062 164694 110122
rect 68800 108762 164756 110062
rect 68800 108702 164694 108762
rect 68800 102376 164756 108702
rect 68816 102316 164756 102376
rect 68800 100744 164756 102316
rect 68816 100684 164756 100744
rect 68800 95100 164756 100684
<< via3 >>
rect 63356 702476 63420 702540
rect 243492 670652 243556 670716
rect 336044 604420 336108 604484
rect 340092 603196 340156 603260
rect 337332 603060 337396 603124
rect 335860 600340 335924 600404
rect 539548 598980 539612 599044
rect 313780 597756 313844 597820
rect 340644 597756 340708 597820
rect 534028 597620 534092 597684
rect 311020 596396 311084 596460
rect 338620 596260 338684 596324
rect 55076 593404 55140 593468
rect 50844 592180 50908 592244
rect 59124 592044 59188 592108
rect 340644 592588 340708 592652
rect 535500 589052 535564 589116
rect 60044 586740 60108 586804
rect 533660 586332 533724 586396
rect 243676 585108 243740 585172
rect 64644 584564 64708 584628
rect 337516 584020 337580 584084
rect 337332 582932 337396 582996
rect 61884 582524 61948 582588
rect 243492 582388 243556 582452
rect 245700 582388 245764 582452
rect 333100 565796 333164 565860
rect 57836 562124 57900 562188
rect 538444 559132 538508 559196
rect 55628 558724 55692 558788
rect 295380 558180 295444 558244
rect 243676 557364 243740 557428
rect 331812 546484 331876 546548
rect 534396 543492 534460 543556
rect 534028 541452 534092 541516
rect 338620 540228 338684 540292
rect 337332 528532 337396 528596
rect 536788 525812 536852 525876
rect 292620 524996 292684 525060
rect 336044 522276 336108 522340
rect 57652 522004 57716 522068
rect 58940 518604 59004 518668
rect 301452 517516 301516 517580
rect 245700 515884 245764 515948
rect 46612 514796 46676 514860
rect 337516 508132 337580 508196
rect 335860 502964 335924 503028
rect 535684 497932 535748 497996
rect 246252 489364 246316 489428
rect 338988 482972 339052 483036
rect 538260 480252 538324 480316
rect 243308 478892 243372 478956
rect 63172 475084 63236 475148
rect 324268 464340 324332 464404
rect 318012 462300 318076 462364
rect 542676 455092 542740 455156
rect 53604 454004 53668 454068
rect 534212 450332 534276 450396
rect 246436 449244 246500 449308
rect 339172 442852 339236 442916
rect 63356 438364 63420 438428
rect 543780 437412 543844 437476
rect 63540 436732 63604 436796
rect 541020 425172 541084 425236
rect 337516 419732 337580 419796
rect 335860 414972 335924 415036
rect 63540 411300 63604 411364
rect 63540 411164 63604 411228
rect 63356 405044 63420 405108
rect 63172 404908 63236 404972
rect 61884 404364 61948 404428
rect 59124 403548 59188 403612
rect 50844 402188 50908 402252
rect 125732 402188 125796 402252
rect 166764 402188 166828 402252
rect 138612 401644 138676 401708
rect 340276 400828 340340 400892
rect 246252 399876 246316 399940
rect 246436 399740 246500 399804
rect 55076 399468 55140 399532
rect 339172 398788 339236 398852
rect 242940 398652 243004 398716
rect 340276 398380 340340 398444
rect 539548 396612 539612 396676
rect 338988 395388 339052 395452
rect 541020 395388 541084 395452
rect 177068 395252 177132 395316
rect 536788 395252 536852 395316
rect 543780 393212 543844 393276
rect 53604 391308 53668 391372
rect 120028 391308 120092 391372
rect 46612 391172 46676 391236
rect 246436 389812 246500 389876
rect 295564 389132 295628 389196
rect 439084 387636 439148 387700
rect 63540 386956 63604 387020
rect 542676 382876 542740 382940
rect 337332 373220 337396 373284
rect 337516 371860 337580 371924
rect 57652 370500 57716 370564
rect 309180 369880 309244 369884
rect 309180 369824 309230 369880
rect 309230 369824 309244 369880
rect 309180 369820 309244 369824
rect 295380 368596 295444 368660
rect 342852 368460 342916 368524
rect 148180 366284 148244 366348
rect 58940 364924 59004 364988
rect 340092 362808 340156 362812
rect 340092 362752 340142 362808
rect 340142 362752 340156 362808
rect 340092 362748 340156 362752
rect 299612 360844 299676 360908
rect 340092 360844 340156 360908
rect 538444 360844 538508 360908
rect 336780 358804 336844 358868
rect 297956 357988 298020 358052
rect 305500 357852 305564 357916
rect 291700 357580 291764 357644
rect 157196 357444 157260 357508
rect 294092 355948 294156 356012
rect 297404 354996 297468 355060
rect 297956 354996 298020 355060
rect 292620 353228 292684 353292
rect 175044 352140 175108 352204
rect 176516 349964 176580 350028
rect 174860 336636 174924 336700
rect 295564 336636 295628 336700
rect 295932 336696 295996 336700
rect 295932 336640 295982 336696
rect 295982 336640 295996 336696
rect 295932 336636 295996 336640
rect 535684 335956 535748 336020
rect 295380 334384 295444 334388
rect 295380 334328 295430 334384
rect 295430 334328 295444 334384
rect 295380 334324 295444 334328
rect 296116 327660 296180 327724
rect 176332 323580 176396 323644
rect 149652 322900 149716 322964
rect 179276 318956 179340 319020
rect 292620 308620 292684 308684
rect 142660 307804 142724 307868
rect 161980 302228 162044 302292
rect 70532 300868 70596 300932
rect 124812 299508 124876 299572
rect 60044 298692 60108 298756
rect 121500 298692 121564 298756
rect 146892 295292 146956 295356
rect 173572 294204 173636 294268
rect 171732 294068 171796 294132
rect 119660 293932 119724 293996
rect 170260 293932 170324 293996
rect 126100 292708 126164 292772
rect 160692 292028 160756 292092
rect 120028 291892 120092 291956
rect 376156 291756 376220 291820
rect 70532 290804 70596 290868
rect 439452 289580 439516 289644
rect 167684 289036 167748 289100
rect 157380 287132 157444 287196
rect 293908 287132 293972 287196
rect 296116 287192 296180 287196
rect 296116 287136 296166 287192
rect 296166 287136 296180 287192
rect 296116 287132 296180 287136
rect 295932 286316 295996 286380
rect 373212 286316 373276 286380
rect 55628 284820 55692 284884
rect 120580 284820 120644 284884
rect 138612 284820 138676 284884
rect 126100 283460 126164 283524
rect 121500 280876 121564 280940
rect 297220 278836 297284 278900
rect 54340 275844 54404 275908
rect 295932 270404 295996 270468
rect 120764 269180 120828 269244
rect 378732 269180 378796 269244
rect 63172 265100 63236 265164
rect 341380 264964 341444 265028
rect 179092 263876 179156 263940
rect 295380 263468 295444 263532
rect 377996 263196 378060 263260
rect 171916 262788 171980 262852
rect 59124 256804 59188 256868
rect 378916 256940 378980 257004
rect 66852 252452 66916 252516
rect 57836 251092 57900 251156
rect 166212 249052 166276 249116
rect 119660 248644 119724 248708
rect 177068 248236 177132 248300
rect 120028 246332 120092 246396
rect 166948 246332 167012 246396
rect 297404 246196 297468 246260
rect 148180 244292 148244 244356
rect 179460 244088 179524 244152
rect 179828 243476 179892 243540
rect 293172 243340 293236 243404
rect 292620 242388 292684 242452
rect 294092 242388 294156 242452
rect 382780 241708 382844 241772
rect 70532 241572 70596 241636
rect 120028 241164 120092 241228
rect 291700 241164 291764 241228
rect 289492 240756 289556 240820
rect 292620 240484 292684 240548
rect 293172 240484 293236 240548
rect 157380 240076 157444 240140
rect 70532 239804 70596 239868
rect 376156 238716 376220 238780
rect 63356 238580 63420 238644
rect 54340 238308 54404 238372
rect 120764 238308 120828 238372
rect 63172 237220 63236 237284
rect 299612 236948 299676 237012
rect 380572 236132 380636 236196
rect 377996 235996 378060 236060
rect 120580 235860 120644 235924
rect 171916 235180 171980 235244
rect 259500 233820 259564 233884
rect 380940 233276 381004 233340
rect 259316 233200 259380 233204
rect 259316 233144 259366 233200
rect 259366 233144 259380 233200
rect 259316 233140 259380 233144
rect 378732 233140 378796 233204
rect 311020 233004 311084 233068
rect 318012 232460 318076 232524
rect 271092 232052 271156 232116
rect 380940 231780 381004 231844
rect 288204 231236 288268 231300
rect 291884 231100 291948 231164
rect 322980 230420 323044 230484
rect 378916 227700 378980 227764
rect 161980 227020 162044 227084
rect 59124 226884 59188 226948
rect 378732 226884 378796 226948
rect 313780 225524 313844 225588
rect 454172 224904 454236 224908
rect 454172 224848 454186 224904
rect 454186 224848 454236 224904
rect 454172 224844 454236 224848
rect 342300 224436 342364 224500
rect 167684 221444 167748 221508
rect 448468 220900 448532 220964
rect 301452 220764 301516 220828
rect 309180 218588 309244 218652
rect 324820 217908 324884 217972
rect 160692 217364 160756 217428
rect 256740 217228 256804 217292
rect 255268 214508 255332 214572
rect 451044 213964 451108 214028
rect 261340 210292 261404 210356
rect 329788 209748 329852 209812
rect 323164 207028 323228 207092
rect 142660 206892 142724 206956
rect 334020 205668 334084 205732
rect 125732 205592 125796 205596
rect 125732 205536 125782 205592
rect 125782 205536 125796 205592
rect 125732 205532 125796 205536
rect 295932 202132 295996 202196
rect 331812 199956 331876 200020
rect 157196 199276 157260 199340
rect 331812 198732 331876 198796
rect 292620 198112 292684 198116
rect 292620 198056 292670 198112
rect 292670 198056 292684 198112
rect 292620 198052 292684 198056
rect 324820 196556 324884 196620
rect 332548 196012 332612 196076
rect 335676 196012 335740 196076
rect 259684 195196 259748 195260
rect 322060 192612 322124 192676
rect 320220 192476 320284 192540
rect 346348 191116 346412 191180
rect 66852 190980 66916 191044
rect 263548 189620 263612 189684
rect 166212 187172 166276 187236
rect 146892 187036 146956 187100
rect 262260 186900 262324 186964
rect 252508 185676 252572 185740
rect 124812 185540 124876 185604
rect 255452 184316 255516 184380
rect 169708 184180 169772 184244
rect 328684 184180 328748 184244
rect 327028 182820 327092 182884
rect 166212 182140 166276 182204
rect 263732 181596 263796 181660
rect 149652 181460 149716 181524
rect 251220 181324 251284 181388
rect 331260 181324 331324 181388
rect 256924 180100 256988 180164
rect 534212 179964 534276 180028
rect 249012 178876 249076 178940
rect 328500 178876 328564 178940
rect 326660 178740 326724 178804
rect 337884 178740 337948 178804
rect 167500 178604 167564 178668
rect 166396 178060 166460 178124
rect 110644 177924 110708 177988
rect 249748 177788 249812 177852
rect 99420 177516 99484 177580
rect 106044 177516 106108 177580
rect 106964 177516 107028 177580
rect 112116 177516 112180 177580
rect 114140 177516 114204 177580
rect 120764 177516 120828 177580
rect 122972 177516 123036 177580
rect 127020 177516 127084 177580
rect 249196 177516 249260 177580
rect 331444 177380 331508 177444
rect 113220 177244 113284 177308
rect 115796 177168 115860 177172
rect 115796 177112 115846 177168
rect 115846 177112 115860 177168
rect 115796 177108 115860 177112
rect 116900 177168 116964 177172
rect 116900 177112 116950 177168
rect 116950 177112 116964 177168
rect 116900 177108 116964 177112
rect 124444 177108 124508 177172
rect 148180 177168 148244 177172
rect 148180 177112 148230 177168
rect 148230 177112 148244 177168
rect 148180 177108 148244 177112
rect 101996 176972 102060 177036
rect 167684 176972 167748 177036
rect 103284 176836 103348 176900
rect 167500 176836 167564 176900
rect 97028 176700 97092 176764
rect 98316 176700 98380 176764
rect 100708 176760 100772 176764
rect 100708 176704 100758 176760
rect 100758 176704 100772 176760
rect 100708 176700 100772 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 109540 176700 109604 176764
rect 118372 176760 118436 176764
rect 118372 176704 118422 176760
rect 118422 176704 118436 176760
rect 118372 176700 118436 176704
rect 125732 176760 125796 176764
rect 125732 176704 125782 176760
rect 125782 176704 125796 176760
rect 125732 176700 125796 176704
rect 130700 176760 130764 176764
rect 130700 176704 130750 176760
rect 130750 176704 130764 176760
rect 130700 176700 130764 176704
rect 131988 176760 132052 176764
rect 131988 176704 132038 176760
rect 132038 176704 132052 176760
rect 131988 176700 132052 176704
rect 134380 176760 134444 176764
rect 134380 176704 134430 176760
rect 134430 176704 134444 176760
rect 134380 176700 134444 176704
rect 135668 176760 135732 176764
rect 135668 176704 135718 176760
rect 135718 176704 135732 176760
rect 135668 176700 135732 176704
rect 158852 176700 158916 176764
rect 260972 176564 261036 176628
rect 128124 176428 128188 176492
rect 327212 176156 327276 176220
rect 254532 175884 254596 175948
rect 265020 175884 265084 175948
rect 104572 175400 104636 175404
rect 104572 175344 104622 175400
rect 104622 175344 104636 175400
rect 104572 175340 104636 175344
rect 121868 175400 121932 175404
rect 121868 175344 121918 175400
rect 121918 175344 121932 175400
rect 121868 175340 121932 175344
rect 129412 175400 129476 175404
rect 129412 175344 129462 175400
rect 129462 175344 129476 175400
rect 129412 175340 129476 175344
rect 133092 175400 133156 175404
rect 133092 175344 133142 175400
rect 133142 175344 133156 175400
rect 133092 175340 133156 175344
rect 119398 174992 119462 174996
rect 119398 174936 119434 174992
rect 119434 174936 119462 174992
rect 119398 174932 119462 174936
rect 249196 174660 249260 174724
rect 265572 174524 265636 174588
rect 342852 174524 342916 174588
rect 533660 174524 533724 174588
rect 321324 174388 321388 174452
rect 249748 174252 249812 174316
rect 252508 173300 252572 173364
rect 326660 173164 326724 173228
rect 249196 172756 249260 172820
rect 327212 170852 327276 170916
rect 259684 170036 259748 170100
rect 335860 167044 335924 167108
rect 327028 166228 327092 166292
rect 166212 164324 166276 164388
rect 263732 163916 263796 163980
rect 166396 161468 166460 161532
rect 328684 161740 328748 161804
rect 259316 160652 259380 160716
rect 269068 160652 269132 160716
rect 337884 159972 337948 160036
rect 535500 159972 535564 160036
rect 256740 158748 256804 158812
rect 337884 158748 337948 158812
rect 167684 157524 167748 157588
rect 167500 157388 167564 157452
rect 255452 157252 255516 157316
rect 251772 152900 251836 152964
rect 260972 152628 261036 152692
rect 329052 150996 329116 151060
rect 259500 149636 259564 149700
rect 293908 149636 293972 149700
rect 458772 149092 458836 149156
rect 396580 147732 396644 147796
rect 451412 147732 451476 147796
rect 450124 146916 450188 146980
rect 292620 144060 292684 144124
rect 166212 143652 166276 143716
rect 449388 143440 449452 143444
rect 449388 143384 449402 143440
rect 449402 143384 449452 143440
rect 449388 143380 449452 143384
rect 265020 142564 265084 142628
rect 263548 142156 263612 142220
rect 262260 141748 262324 141812
rect 307340 141612 307404 141676
rect 251220 140796 251284 140860
rect 255268 140388 255332 140452
rect 256924 139844 256988 139908
rect 167684 138076 167748 138140
rect 328500 138620 328564 138684
rect 307156 136988 307220 137052
rect 254532 136580 254596 136644
rect 341380 136580 341444 136644
rect 307340 134404 307404 134468
rect 451044 133452 451108 133516
rect 166396 131412 166460 131476
rect 451412 132092 451476 132156
rect 331444 131276 331508 131340
rect 342300 131140 342364 131204
rect 167500 129780 167564 129844
rect 169156 128420 169220 128484
rect 301636 128420 301700 128484
rect 301452 126380 301516 126444
rect 251772 126244 251836 126308
rect 322980 125428 323044 125492
rect 329052 122980 329116 123044
rect 335676 122844 335740 122908
rect 451044 121484 451108 121548
rect 458772 118764 458836 118828
rect 454172 118084 454236 118148
rect 346348 117268 346412 117332
rect 323164 116996 323228 117060
rect 329788 114548 329852 114612
rect 291700 113868 291764 113932
rect 252508 113732 252572 113796
rect 305684 113596 305748 113660
rect 299980 112644 300044 112708
rect 396580 112372 396644 112436
rect 449940 112372 450004 112436
rect 331260 111828 331324 111892
rect 334020 111012 334084 111076
rect 252508 110740 252572 110804
rect 251220 109108 251284 109172
rect 324268 108564 324332 108628
rect 322060 108292 322124 108356
rect 382780 106388 382844 106452
rect 373212 102716 373276 102780
rect 449388 100948 449452 101012
rect 288204 99996 288268 100060
rect 304212 99724 304276 99788
rect 538260 100676 538324 100740
rect 449388 99724 449452 99788
rect 332548 98092 332612 98156
rect 306972 97820 307036 97884
rect 450124 96052 450188 96116
rect 261340 95372 261404 95436
rect 333100 95644 333164 95708
rect 534396 95236 534460 95300
rect 324268 95100 324332 95164
rect 106478 94828 106542 94892
rect 106780 94828 106844 94892
rect 151766 94888 151830 94892
rect 151766 94832 151782 94888
rect 151782 94832 151830 94888
rect 151766 94828 151830 94832
rect 94918 94752 94982 94756
rect 94918 94696 94962 94752
rect 94962 94696 94982 94752
rect 94918 94692 94982 94696
rect 113142 94752 113206 94756
rect 113142 94696 113178 94752
rect 113178 94696 113206 94752
rect 113142 94692 113206 94696
rect 115862 94752 115926 94756
rect 115862 94696 115902 94752
rect 115902 94696 115926 94752
rect 115862 94692 115926 94696
rect 126470 94752 126534 94756
rect 126470 94696 126518 94752
rect 126518 94696 126534 94752
rect 126470 94692 126534 94696
rect 128124 93876 128188 93940
rect 166212 93876 166276 93940
rect 171732 93740 171796 93804
rect 130700 93664 130764 93668
rect 130700 93608 130750 93664
rect 130750 93608 130764 93664
rect 130700 93604 130764 93608
rect 173572 93604 173636 93668
rect 97212 93528 97276 93532
rect 97212 93472 97262 93528
rect 97262 93472 97276 93528
rect 97212 93468 97276 93472
rect 113772 93528 113836 93532
rect 113772 93472 113822 93528
rect 113822 93472 113836 93528
rect 113772 93468 113836 93472
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 87092 92440 87156 92444
rect 87092 92384 87142 92440
rect 87142 92384 87156 92440
rect 87092 92380 87156 92384
rect 98132 92440 98196 92444
rect 98132 92384 98182 92440
rect 98182 92384 98196 92440
rect 98132 92380 98196 92384
rect 98500 92380 98564 92444
rect 106780 92380 106844 92444
rect 116716 92440 116780 92444
rect 116716 92384 116766 92440
rect 116766 92384 116780 92440
rect 116716 92380 116780 92384
rect 120212 92380 120276 92444
rect 124076 92440 124140 92444
rect 124076 92384 124090 92440
rect 124090 92384 124140 92440
rect 124076 92380 124140 92384
rect 125732 92440 125796 92444
rect 125732 92384 125782 92440
rect 125782 92384 125796 92440
rect 125732 92380 125796 92384
rect 129412 92440 129476 92444
rect 129412 92384 129462 92440
rect 129462 92384 129476 92440
rect 129412 92380 129476 92384
rect 133092 92440 133156 92444
rect 133092 92384 133142 92440
rect 133142 92384 133156 92440
rect 133092 92380 133156 92384
rect 135668 92440 135732 92444
rect 135668 92384 135718 92440
rect 135718 92384 135732 92440
rect 135668 92380 135732 92384
rect 151492 92440 151556 92444
rect 151492 92384 151542 92440
rect 151542 92384 151556 92440
rect 151492 92380 151556 92384
rect 152044 92440 152108 92444
rect 152044 92384 152094 92440
rect 152094 92384 152108 92440
rect 152044 92380 152108 92384
rect 170260 92380 170324 92444
rect 114140 92244 114204 92308
rect 119660 92108 119724 92172
rect 167684 92108 167748 92172
rect 99604 91700 99668 91764
rect 117084 91760 117148 91764
rect 117084 91704 117134 91760
rect 117134 91704 117148 91760
rect 117084 91700 117148 91704
rect 305500 91700 305564 91764
rect 109172 91564 109236 91628
rect 131988 91564 132052 91628
rect 151308 91624 151372 91628
rect 151308 91568 151358 91624
rect 151358 91568 151372 91624
rect 151308 91564 151372 91568
rect 122788 91488 122852 91492
rect 122788 91432 122838 91488
rect 122838 91432 122852 91488
rect 122788 91428 122852 91432
rect 101812 91292 101876 91356
rect 104204 91292 104268 91356
rect 107700 91292 107764 91356
rect 112300 91292 112364 91356
rect 124444 91292 124508 91356
rect 74764 91156 74828 91220
rect 84332 91156 84396 91220
rect 85620 91156 85684 91220
rect 86724 91156 86788 91220
rect 88932 91156 88996 91220
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 93900 91156 93964 91220
rect 96108 91156 96172 91220
rect 97028 91156 97092 91220
rect 99236 91216 99300 91220
rect 99236 91160 99286 91216
rect 99286 91160 99300 91216
rect 99236 91156 99300 91160
rect 100524 91156 100588 91220
rect 101628 91216 101692 91220
rect 101628 91160 101678 91216
rect 101678 91160 101692 91216
rect 101628 91156 101692 91160
rect 101996 91216 102060 91220
rect 101996 91160 102046 91216
rect 102046 91160 102060 91216
rect 101996 91156 102060 91160
rect 102916 91216 102980 91220
rect 102916 91160 102966 91216
rect 102966 91160 102980 91216
rect 102916 91156 102980 91160
rect 103284 91216 103348 91220
rect 103284 91160 103334 91216
rect 103334 91160 103348 91216
rect 103284 91156 103348 91160
rect 104572 91156 104636 91220
rect 105124 91156 105188 91220
rect 106044 91156 106108 91220
rect 106412 91156 106476 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 110644 91156 110708 91220
rect 111196 91156 111260 91220
rect 111932 91156 111996 91220
rect 115060 91156 115124 91220
rect 115428 91156 115492 91220
rect 118004 91216 118068 91220
rect 118004 91160 118054 91216
rect 118054 91160 118068 91216
rect 118004 91156 118068 91160
rect 118188 91156 118252 91220
rect 119844 91216 119908 91220
rect 119844 91160 119894 91216
rect 119894 91160 119908 91216
rect 119844 91156 119908 91160
rect 120580 91156 120644 91220
rect 121684 91156 121748 91220
rect 122052 91156 122116 91220
rect 122972 91156 123036 91220
rect 125364 91156 125428 91220
rect 126652 91156 126716 91220
rect 134380 91156 134444 91220
rect 166396 91020 166460 91084
rect 380572 91020 380636 91084
rect 307156 88980 307220 89044
rect 179092 86124 179156 86188
rect 169156 85444 169220 85508
rect 176332 84764 176396 84828
rect 449388 84764 449452 84828
rect 295380 84280 295444 84284
rect 295380 84224 295394 84280
rect 295394 84224 295444 84280
rect 295380 84220 295444 84224
rect 167500 80004 167564 80068
rect 304212 72388 304276 72452
rect 301636 68172 301700 68236
rect 177068 65452 177132 65516
rect 269068 60072 269132 60076
rect 269068 60016 269118 60072
rect 269118 60016 269132 60072
rect 269068 60012 269132 60016
rect 271092 46820 271156 46884
rect 448468 45460 448532 45524
rect 340092 42740 340156 42804
rect 451044 42740 451108 42804
rect 340092 42060 340156 42124
rect 179828 32404 179892 32468
rect 305684 29548 305748 29612
rect 176516 28188 176580 28252
rect 336780 26208 336844 26212
rect 336780 26152 336830 26208
rect 336830 26152 336844 26208
rect 336780 26148 336844 26152
rect 299980 24108 300044 24172
rect 449940 22612 450004 22676
rect 175044 21932 175108 21996
rect 289492 19212 289556 19276
rect 179276 15132 179340 15196
rect 64644 12956 64708 13020
rect 269068 11732 269132 11796
rect 297220 11732 297284 11796
rect 301452 10236 301516 10300
rect 174860 8196 174924 8260
rect 179460 5476 179524 5540
rect 251220 3436 251284 3500
rect 265572 3436 265636 3500
rect 169708 3300 169772 3364
rect 306972 2620 307036 2684
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55075 593468 55141 593469
rect 55075 593404 55076 593468
rect 55140 593404 55141 593468
rect 55075 593403 55141 593404
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 50843 592244 50909 592245
rect 50843 592180 50844 592244
rect 50908 592180 50909 592244
rect 50843 592179 50909 592180
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46611 514860 46677 514861
rect 46611 514796 46612 514860
rect 46676 514796 46677 514860
rect 46611 514795 46677 514796
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 46614 391237 46674 514795
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46611 391236 46677 391237
rect 46611 391172 46612 391236
rect 46676 391172 46677 391236
rect 46611 391171 46677 391172
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 372454 47414 407898
rect 50846 402253 50906 592179
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 53603 454068 53669 454069
rect 53603 454004 53604 454068
rect 53668 454004 53669 454068
rect 53603 454003 53669 454004
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 50843 402252 50909 402253
rect 50843 402188 50844 402252
rect 50908 402188 50909 402252
rect 50843 402187 50909 402188
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 376954 51914 412398
rect 53606 391373 53666 454003
rect 55078 399533 55138 593403
rect 55794 561454 56414 596898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 63355 702540 63421 702541
rect 63355 702476 63356 702540
rect 63420 702476 63421 702540
rect 63355 702475 63421 702476
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 59123 592108 59189 592109
rect 59123 592044 59124 592108
rect 59188 592044 59189 592108
rect 59123 592043 59189 592044
rect 57835 562188 57901 562189
rect 57835 562124 57836 562188
rect 57900 562124 57901 562188
rect 57835 562123 57901 562124
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55627 558788 55693 558789
rect 55627 558724 55628 558788
rect 55692 558724 55693 558788
rect 55627 558723 55693 558724
rect 55075 399532 55141 399533
rect 55075 399468 55076 399532
rect 55140 399468 55141 399532
rect 55075 399467 55141 399468
rect 53603 391372 53669 391373
rect 53603 391308 53604 391372
rect 53668 391308 53669 391372
rect 53603 391307 53669 391308
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 55630 284885 55690 558723
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 57651 522068 57717 522069
rect 57651 522004 57652 522068
rect 57716 522004 57717 522068
rect 57651 522003 57717 522004
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 57654 370565 57714 522003
rect 57651 370564 57717 370565
rect 57651 370500 57652 370564
rect 57716 370500 57717 370564
rect 57651 370499 57717 370500
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55627 284884 55693 284885
rect 55627 284820 55628 284884
rect 55692 284820 55693 284884
rect 55627 284819 55693 284820
rect 54339 275908 54405 275909
rect 54339 275844 54340 275908
rect 54404 275844 54405 275908
rect 54339 275843 54405 275844
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 54342 238373 54402 275843
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 54339 238372 54405 238373
rect 54339 238308 54340 238372
rect 54404 238308 54405 238372
rect 54339 238307 54405 238308
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 237454 56414 272898
rect 57838 251157 57898 562123
rect 58939 518668 59005 518669
rect 58939 518604 58940 518668
rect 59004 518604 59005 518668
rect 58939 518603 59005 518604
rect 58942 364989 59002 518603
rect 59126 403613 59186 592043
rect 60043 586804 60109 586805
rect 60043 586740 60044 586804
rect 60108 586740 60109 586804
rect 60043 586739 60109 586740
rect 59123 403612 59189 403613
rect 59123 403548 59124 403612
rect 59188 403548 59189 403612
rect 59123 403547 59189 403548
rect 58939 364988 59005 364989
rect 58939 364924 58940 364988
rect 59004 364924 59005 364988
rect 58939 364923 59005 364924
rect 60046 298757 60106 586739
rect 60294 565954 60914 601398
rect 61883 582588 61949 582589
rect 61883 582524 61884 582588
rect 61948 582524 61949 582588
rect 61883 582523 61949 582524
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 61886 404429 61946 582523
rect 63171 475148 63237 475149
rect 63171 475084 63172 475148
rect 63236 475084 63237 475148
rect 63171 475083 63237 475084
rect 63174 404973 63234 475083
rect 63358 438429 63418 702475
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 587000 65414 605898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 587000 69914 610398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 587000 74414 614898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 587000 78914 619398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 587000 83414 587898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 587000 87914 592398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 587000 92414 596898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 587000 96914 601398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 587000 101414 605898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 587000 105914 610398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 587000 110414 614898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 587000 114914 619398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 587000 119414 587898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 587000 123914 592398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 587000 128414 596898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 587000 132914 601398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 587000 137414 605898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 587000 141914 610398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 587000 146414 614898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 587000 150914 619398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 587000 155414 587898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 587000 159914 592398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 587000 164414 596898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 587000 168914 601398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 587000 173414 605898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 587000 177914 610398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 587000 182414 614898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 587000 186914 619398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 587000 191414 587898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 587000 195914 592398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 587000 200414 596898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 587000 204914 601398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 587000 209414 605898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 587000 213914 610398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 587000 218414 614898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 587000 222914 619398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 587000 227414 587898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 587000 231914 592398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 587000 236414 596898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 243491 670716 243557 670717
rect 243491 670652 243492 670716
rect 243556 670652 243557 670716
rect 243491 670651 243557 670652
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 587000 240914 601398
rect 64643 584628 64709 584629
rect 64643 584564 64644 584628
rect 64708 584564 64709 584628
rect 64643 584563 64709 584564
rect 63355 438428 63421 438429
rect 63355 438364 63356 438428
rect 63420 438364 63421 438428
rect 63355 438363 63421 438364
rect 63358 405109 63418 438363
rect 63539 436796 63605 436797
rect 63539 436732 63540 436796
rect 63604 436732 63605 436796
rect 63539 436731 63605 436732
rect 63542 411365 63602 436731
rect 63539 411364 63605 411365
rect 63539 411300 63540 411364
rect 63604 411300 63605 411364
rect 63539 411299 63605 411300
rect 63539 411228 63605 411229
rect 63539 411164 63540 411228
rect 63604 411164 63605 411228
rect 63539 411163 63605 411164
rect 63355 405108 63421 405109
rect 63355 405044 63356 405108
rect 63420 405044 63421 405108
rect 63355 405043 63421 405044
rect 63171 404972 63237 404973
rect 63171 404908 63172 404972
rect 63236 404908 63237 404972
rect 63171 404907 63237 404908
rect 61883 404428 61949 404429
rect 61883 404364 61884 404428
rect 61948 404364 61949 404428
rect 61883 404363 61949 404364
rect 63174 402990 63234 404907
rect 63174 402930 63418 402990
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60043 298756 60109 298757
rect 60043 298692 60044 298756
rect 60108 298692 60109 298756
rect 60043 298691 60109 298692
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 59123 256868 59189 256869
rect 59123 256804 59124 256868
rect 59188 256804 59189 256868
rect 59123 256803 59189 256804
rect 57835 251156 57901 251157
rect 57835 251092 57836 251156
rect 57900 251092 57901 251156
rect 57835 251091 57901 251092
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 59126 226949 59186 256803
rect 60294 241954 60914 277398
rect 63171 265164 63237 265165
rect 63171 265100 63172 265164
rect 63236 265100 63237 265164
rect 63171 265099 63237 265100
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 59123 226948 59189 226949
rect 59123 226884 59124 226948
rect 59188 226884 59189 226948
rect 59123 226883 59189 226884
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 241398
rect 63174 237285 63234 265099
rect 63358 238645 63418 402930
rect 63542 387021 63602 411163
rect 63539 387020 63605 387021
rect 63539 386956 63540 387020
rect 63604 386956 63605 387020
rect 63539 386955 63605 386956
rect 63355 238644 63421 238645
rect 63355 238580 63356 238644
rect 63420 238580 63421 238644
rect 63355 238579 63421 238580
rect 63171 237284 63237 237285
rect 63171 237220 63172 237284
rect 63236 237220 63237 237284
rect 63171 237219 63237 237220
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 64646 13021 64706 584563
rect 243494 582453 243554 670651
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 587000 245414 605898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 243675 585172 243741 585173
rect 243675 585108 243676 585172
rect 243740 585108 243741 585172
rect 243675 585107 243741 585108
rect 243491 582452 243557 582453
rect 243491 582388 243492 582452
rect 243556 582388 243557 582452
rect 243491 582387 243557 582388
rect 68208 579454 68528 579486
rect 68208 579218 68250 579454
rect 68486 579218 68528 579454
rect 68208 579134 68528 579218
rect 68208 578898 68250 579134
rect 68486 578898 68528 579134
rect 68208 578866 68528 578898
rect 98928 579454 99248 579486
rect 98928 579218 98970 579454
rect 99206 579218 99248 579454
rect 98928 579134 99248 579218
rect 98928 578898 98970 579134
rect 99206 578898 99248 579134
rect 98928 578866 99248 578898
rect 129648 579454 129968 579486
rect 129648 579218 129690 579454
rect 129926 579218 129968 579454
rect 129648 579134 129968 579218
rect 129648 578898 129690 579134
rect 129926 578898 129968 579134
rect 129648 578866 129968 578898
rect 160368 579454 160688 579486
rect 160368 579218 160410 579454
rect 160646 579218 160688 579454
rect 160368 579134 160688 579218
rect 160368 578898 160410 579134
rect 160646 578898 160688 579134
rect 160368 578866 160688 578898
rect 191088 579454 191408 579486
rect 191088 579218 191130 579454
rect 191366 579218 191408 579454
rect 191088 579134 191408 579218
rect 191088 578898 191130 579134
rect 191366 578898 191408 579134
rect 191088 578866 191408 578898
rect 221808 579454 222128 579486
rect 221808 579218 221850 579454
rect 222086 579218 222128 579454
rect 221808 579134 222128 579218
rect 221808 578898 221850 579134
rect 222086 578898 222128 579134
rect 221808 578866 222128 578898
rect 243678 557429 243738 585107
rect 245699 582452 245765 582453
rect 245699 582388 245700 582452
rect 245764 582388 245765 582452
rect 245699 582387 245765 582388
rect 243675 557428 243741 557429
rect 243675 557364 243676 557428
rect 243740 557364 243741 557428
rect 243675 557363 243741 557364
rect 83568 547954 83888 547986
rect 83568 547718 83610 547954
rect 83846 547718 83888 547954
rect 83568 547634 83888 547718
rect 83568 547398 83610 547634
rect 83846 547398 83888 547634
rect 83568 547366 83888 547398
rect 114288 547954 114608 547986
rect 114288 547718 114330 547954
rect 114566 547718 114608 547954
rect 114288 547634 114608 547718
rect 114288 547398 114330 547634
rect 114566 547398 114608 547634
rect 114288 547366 114608 547398
rect 145008 547954 145328 547986
rect 145008 547718 145050 547954
rect 145286 547718 145328 547954
rect 145008 547634 145328 547718
rect 145008 547398 145050 547634
rect 145286 547398 145328 547634
rect 145008 547366 145328 547398
rect 175728 547954 176048 547986
rect 175728 547718 175770 547954
rect 176006 547718 176048 547954
rect 175728 547634 176048 547718
rect 175728 547398 175770 547634
rect 176006 547398 176048 547634
rect 175728 547366 176048 547398
rect 206448 547954 206768 547986
rect 206448 547718 206490 547954
rect 206726 547718 206768 547954
rect 206448 547634 206768 547718
rect 206448 547398 206490 547634
rect 206726 547398 206768 547634
rect 206448 547366 206768 547398
rect 237168 547954 237488 547986
rect 237168 547718 237210 547954
rect 237446 547718 237488 547954
rect 237168 547634 237488 547718
rect 237168 547398 237210 547634
rect 237446 547398 237488 547634
rect 237168 547366 237488 547398
rect 68208 543454 68528 543486
rect 68208 543218 68250 543454
rect 68486 543218 68528 543454
rect 68208 543134 68528 543218
rect 68208 542898 68250 543134
rect 68486 542898 68528 543134
rect 68208 542866 68528 542898
rect 98928 543454 99248 543486
rect 98928 543218 98970 543454
rect 99206 543218 99248 543454
rect 98928 543134 99248 543218
rect 98928 542898 98970 543134
rect 99206 542898 99248 543134
rect 98928 542866 99248 542898
rect 129648 543454 129968 543486
rect 129648 543218 129690 543454
rect 129926 543218 129968 543454
rect 129648 543134 129968 543218
rect 129648 542898 129690 543134
rect 129926 542898 129968 543134
rect 129648 542866 129968 542898
rect 160368 543454 160688 543486
rect 160368 543218 160410 543454
rect 160646 543218 160688 543454
rect 160368 543134 160688 543218
rect 160368 542898 160410 543134
rect 160646 542898 160688 543134
rect 160368 542866 160688 542898
rect 191088 543454 191408 543486
rect 191088 543218 191130 543454
rect 191366 543218 191408 543454
rect 191088 543134 191408 543218
rect 191088 542898 191130 543134
rect 191366 542898 191408 543134
rect 191088 542866 191408 542898
rect 221808 543454 222128 543486
rect 221808 543218 221850 543454
rect 222086 543218 222128 543454
rect 221808 543134 222128 543218
rect 221808 542898 221850 543134
rect 222086 542898 222128 543134
rect 221808 542866 222128 542898
rect 245702 515949 245762 582387
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 245699 515948 245765 515949
rect 245699 515884 245700 515948
rect 245764 515884 245765 515948
rect 245699 515883 245765 515884
rect 83568 511954 83888 511986
rect 83568 511718 83610 511954
rect 83846 511718 83888 511954
rect 83568 511634 83888 511718
rect 83568 511398 83610 511634
rect 83846 511398 83888 511634
rect 83568 511366 83888 511398
rect 114288 511954 114608 511986
rect 114288 511718 114330 511954
rect 114566 511718 114608 511954
rect 114288 511634 114608 511718
rect 114288 511398 114330 511634
rect 114566 511398 114608 511634
rect 114288 511366 114608 511398
rect 145008 511954 145328 511986
rect 145008 511718 145050 511954
rect 145286 511718 145328 511954
rect 145008 511634 145328 511718
rect 145008 511398 145050 511634
rect 145286 511398 145328 511634
rect 145008 511366 145328 511398
rect 175728 511954 176048 511986
rect 175728 511718 175770 511954
rect 176006 511718 176048 511954
rect 175728 511634 176048 511718
rect 175728 511398 175770 511634
rect 176006 511398 176048 511634
rect 175728 511366 176048 511398
rect 206448 511954 206768 511986
rect 206448 511718 206490 511954
rect 206726 511718 206768 511954
rect 206448 511634 206768 511718
rect 206448 511398 206490 511634
rect 206726 511398 206768 511634
rect 206448 511366 206768 511398
rect 237168 511954 237488 511986
rect 237168 511718 237210 511954
rect 237446 511718 237488 511954
rect 237168 511634 237488 511718
rect 237168 511398 237210 511634
rect 237446 511398 237488 511634
rect 237168 511366 237488 511398
rect 68208 507454 68528 507486
rect 68208 507218 68250 507454
rect 68486 507218 68528 507454
rect 68208 507134 68528 507218
rect 68208 506898 68250 507134
rect 68486 506898 68528 507134
rect 68208 506866 68528 506898
rect 98928 507454 99248 507486
rect 98928 507218 98970 507454
rect 99206 507218 99248 507454
rect 98928 507134 99248 507218
rect 98928 506898 98970 507134
rect 99206 506898 99248 507134
rect 98928 506866 99248 506898
rect 129648 507454 129968 507486
rect 129648 507218 129690 507454
rect 129926 507218 129968 507454
rect 129648 507134 129968 507218
rect 129648 506898 129690 507134
rect 129926 506898 129968 507134
rect 129648 506866 129968 506898
rect 160368 507454 160688 507486
rect 160368 507218 160410 507454
rect 160646 507218 160688 507454
rect 160368 507134 160688 507218
rect 160368 506898 160410 507134
rect 160646 506898 160688 507134
rect 160368 506866 160688 506898
rect 191088 507454 191408 507486
rect 191088 507218 191130 507454
rect 191366 507218 191408 507454
rect 191088 507134 191408 507218
rect 191088 506898 191130 507134
rect 191366 506898 191408 507134
rect 191088 506866 191408 506898
rect 221808 507454 222128 507486
rect 221808 507218 221850 507454
rect 222086 507218 222128 507454
rect 221808 507134 222128 507218
rect 221808 506898 221850 507134
rect 222086 506898 222128 507134
rect 221808 506866 222128 506898
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 246251 489428 246317 489429
rect 246251 489364 246252 489428
rect 246316 489364 246317 489428
rect 246251 489363 246317 489364
rect 243307 478956 243373 478957
rect 243307 478892 243308 478956
rect 243372 478892 243373 478956
rect 243307 478891 243373 478892
rect 83568 475954 83888 475986
rect 83568 475718 83610 475954
rect 83846 475718 83888 475954
rect 83568 475634 83888 475718
rect 83568 475398 83610 475634
rect 83846 475398 83888 475634
rect 83568 475366 83888 475398
rect 114288 475954 114608 475986
rect 114288 475718 114330 475954
rect 114566 475718 114608 475954
rect 114288 475634 114608 475718
rect 114288 475398 114330 475634
rect 114566 475398 114608 475634
rect 114288 475366 114608 475398
rect 145008 475954 145328 475986
rect 145008 475718 145050 475954
rect 145286 475718 145328 475954
rect 145008 475634 145328 475718
rect 145008 475398 145050 475634
rect 145286 475398 145328 475634
rect 145008 475366 145328 475398
rect 175728 475954 176048 475986
rect 175728 475718 175770 475954
rect 176006 475718 176048 475954
rect 175728 475634 176048 475718
rect 175728 475398 175770 475634
rect 176006 475398 176048 475634
rect 175728 475366 176048 475398
rect 206448 475954 206768 475986
rect 206448 475718 206490 475954
rect 206726 475718 206768 475954
rect 206448 475634 206768 475718
rect 206448 475398 206490 475634
rect 206726 475398 206768 475634
rect 206448 475366 206768 475398
rect 237168 475954 237488 475986
rect 237168 475718 237210 475954
rect 237446 475718 237488 475954
rect 237168 475634 237488 475718
rect 237168 475398 237210 475634
rect 237446 475398 237488 475634
rect 237168 475366 237488 475398
rect 68208 471454 68528 471486
rect 68208 471218 68250 471454
rect 68486 471218 68528 471454
rect 68208 471134 68528 471218
rect 68208 470898 68250 471134
rect 68486 470898 68528 471134
rect 68208 470866 68528 470898
rect 98928 471454 99248 471486
rect 98928 471218 98970 471454
rect 99206 471218 99248 471454
rect 98928 471134 99248 471218
rect 98928 470898 98970 471134
rect 99206 470898 99248 471134
rect 98928 470866 99248 470898
rect 129648 471454 129968 471486
rect 129648 471218 129690 471454
rect 129926 471218 129968 471454
rect 129648 471134 129968 471218
rect 129648 470898 129690 471134
rect 129926 470898 129968 471134
rect 129648 470866 129968 470898
rect 160368 471454 160688 471486
rect 160368 471218 160410 471454
rect 160646 471218 160688 471454
rect 160368 471134 160688 471218
rect 160368 470898 160410 471134
rect 160646 470898 160688 471134
rect 160368 470866 160688 470898
rect 191088 471454 191408 471486
rect 191088 471218 191130 471454
rect 191366 471218 191408 471454
rect 191088 471134 191408 471218
rect 191088 470898 191130 471134
rect 191366 470898 191408 471134
rect 191088 470866 191408 470898
rect 221808 471454 222128 471486
rect 221808 471218 221850 471454
rect 222086 471218 222128 471454
rect 221808 471134 222128 471218
rect 221808 470898 221850 471134
rect 222086 470898 222128 471134
rect 221808 470866 222128 470898
rect 243310 470610 243370 478891
rect 242942 470550 243370 470610
rect 83568 439954 83888 439986
rect 83568 439718 83610 439954
rect 83846 439718 83888 439954
rect 83568 439634 83888 439718
rect 83568 439398 83610 439634
rect 83846 439398 83888 439634
rect 83568 439366 83888 439398
rect 114288 439954 114608 439986
rect 114288 439718 114330 439954
rect 114566 439718 114608 439954
rect 114288 439634 114608 439718
rect 114288 439398 114330 439634
rect 114566 439398 114608 439634
rect 114288 439366 114608 439398
rect 145008 439954 145328 439986
rect 145008 439718 145050 439954
rect 145286 439718 145328 439954
rect 145008 439634 145328 439718
rect 145008 439398 145050 439634
rect 145286 439398 145328 439634
rect 145008 439366 145328 439398
rect 175728 439954 176048 439986
rect 175728 439718 175770 439954
rect 176006 439718 176048 439954
rect 175728 439634 176048 439718
rect 175728 439398 175770 439634
rect 176006 439398 176048 439634
rect 175728 439366 176048 439398
rect 206448 439954 206768 439986
rect 206448 439718 206490 439954
rect 206726 439718 206768 439954
rect 206448 439634 206768 439718
rect 206448 439398 206490 439634
rect 206726 439398 206768 439634
rect 206448 439366 206768 439398
rect 237168 439954 237488 439986
rect 237168 439718 237210 439954
rect 237446 439718 237488 439954
rect 237168 439634 237488 439718
rect 237168 439398 237210 439634
rect 237446 439398 237488 439634
rect 237168 439366 237488 439398
rect 68208 435454 68528 435486
rect 68208 435218 68250 435454
rect 68486 435218 68528 435454
rect 68208 435134 68528 435218
rect 68208 434898 68250 435134
rect 68486 434898 68528 435134
rect 68208 434866 68528 434898
rect 98928 435454 99248 435486
rect 98928 435218 98970 435454
rect 99206 435218 99248 435454
rect 98928 435134 99248 435218
rect 98928 434898 98970 435134
rect 99206 434898 99248 435134
rect 98928 434866 99248 434898
rect 129648 435454 129968 435486
rect 129648 435218 129690 435454
rect 129926 435218 129968 435454
rect 129648 435134 129968 435218
rect 129648 434898 129690 435134
rect 129926 434898 129968 435134
rect 129648 434866 129968 434898
rect 160368 435454 160688 435486
rect 160368 435218 160410 435454
rect 160646 435218 160688 435454
rect 160368 435134 160688 435218
rect 160368 434898 160410 435134
rect 160646 434898 160688 435134
rect 160368 434866 160688 434898
rect 191088 435454 191408 435486
rect 191088 435218 191130 435454
rect 191366 435218 191408 435454
rect 191088 435134 191408 435218
rect 191088 434898 191130 435134
rect 191366 434898 191408 435134
rect 191088 434866 191408 434898
rect 221808 435454 222128 435486
rect 221808 435218 221850 435454
rect 222086 435218 222128 435454
rect 221808 435134 222128 435218
rect 221808 434898 221850 435134
rect 222086 434898 222128 435134
rect 221808 434866 222128 434898
rect 64794 390454 65414 403000
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 69294 394954 69914 403000
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 294000 69914 322398
rect 73794 399454 74414 403000
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 70531 300932 70597 300933
rect 70531 300868 70532 300932
rect 70596 300868 70597 300932
rect 70531 300867 70597 300868
rect 70534 290869 70594 300867
rect 73794 294000 74414 326898
rect 78294 367954 78914 403000
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 294000 78914 295398
rect 82794 372454 83414 403000
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 294000 83414 299898
rect 87294 376954 87914 403000
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 294000 87914 304398
rect 91794 381454 92414 403000
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 96294 385954 96914 403000
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 294000 96914 313398
rect 100794 390454 101414 403000
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 294000 101414 317898
rect 105294 394954 105914 403000
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 294000 105914 322398
rect 109794 399454 110414 403000
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 114294 367954 114914 403000
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 294000 114914 295398
rect 118794 372454 119414 403000
rect 120027 391372 120093 391373
rect 120027 391308 120028 391372
rect 120092 391308 120093 391372
rect 120027 391307 120093 391308
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 294000 119414 299898
rect 119659 293996 119725 293997
rect 119659 293932 119660 293996
rect 119724 293932 119725 293996
rect 119659 293931 119725 293932
rect 70531 290868 70597 290869
rect 70531 290804 70532 290868
rect 70596 290804 70597 290868
rect 70531 290803 70597 290804
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 89568 259954 89888 259986
rect 89568 259718 89610 259954
rect 89846 259718 89888 259954
rect 89568 259634 89888 259718
rect 89568 259398 89610 259634
rect 89846 259398 89888 259634
rect 89568 259366 89888 259398
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 66851 252516 66917 252517
rect 66851 252452 66852 252516
rect 66916 252452 66917 252516
rect 66851 252451 66917 252452
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 66854 191045 66914 252451
rect 119662 248709 119722 293931
rect 120030 291957 120090 391307
rect 123294 376954 123914 403000
rect 125731 402252 125797 402253
rect 125731 402188 125732 402252
rect 125796 402188 125797 402252
rect 125731 402187 125797 402188
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 121499 298756 121565 298757
rect 121499 298692 121500 298756
rect 121564 298692 121565 298756
rect 121499 298691 121565 298692
rect 120027 291956 120093 291957
rect 120027 291892 120028 291956
rect 120092 291892 120093 291956
rect 120027 291891 120093 291892
rect 120579 284884 120645 284885
rect 120579 284820 120580 284884
rect 120644 284820 120645 284884
rect 120579 284819 120645 284820
rect 119659 248708 119725 248709
rect 119659 248644 119660 248708
rect 119724 248644 119725 248708
rect 119659 248643 119725 248644
rect 120027 246396 120093 246397
rect 120027 246332 120028 246396
rect 120092 246332 120093 246396
rect 120027 246331 120093 246332
rect 70531 241636 70597 241637
rect 70531 241572 70532 241636
rect 70596 241572 70597 241636
rect 70531 241571 70597 241572
rect 70534 239869 70594 241571
rect 120030 241229 120090 246331
rect 120027 241228 120093 241229
rect 120027 241164 120028 241228
rect 120092 241164 120093 241228
rect 120027 241163 120093 241164
rect 70531 239868 70597 239869
rect 70531 239804 70532 239868
rect 70596 239804 70597 239868
rect 70531 239803 70597 239804
rect 69294 214954 69914 238000
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 66851 191044 66917 191045
rect 66851 190980 66852 191044
rect 66916 190980 66917 191044
rect 66851 190979 66917 190980
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 176600 69914 178398
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 78294 223954 78914 238000
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 176600 78914 187398
rect 82794 228454 83414 238000
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 176600 83414 191898
rect 87294 232954 87914 238000
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 176600 87914 196398
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 105294 214954 105914 238000
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 99419 177580 99485 177581
rect 99419 177516 99420 177580
rect 99484 177516 99485 177580
rect 99419 177515 99485 177516
rect 97027 176764 97093 176765
rect 97027 176700 97028 176764
rect 97092 176700 97093 176764
rect 97027 176699 97093 176700
rect 98315 176764 98381 176765
rect 98315 176700 98316 176764
rect 98380 176700 98381 176764
rect 98315 176699 98381 176700
rect 97030 175130 97090 176699
rect 96960 175070 97090 175130
rect 98318 175130 98378 176699
rect 99422 175130 99482 177515
rect 101995 177036 102061 177037
rect 101995 176972 101996 177036
rect 102060 176972 102061 177036
rect 101995 176971 102061 176972
rect 100707 176764 100773 176765
rect 100707 176700 100708 176764
rect 100772 176700 100773 176764
rect 100707 176699 100773 176700
rect 98318 175070 98380 175130
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 176699
rect 101998 175130 102058 176971
rect 103283 176900 103349 176901
rect 103283 176836 103284 176900
rect 103348 176836 103349 176900
rect 103283 176835 103349 176836
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176835
rect 105294 176600 105914 178398
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 106043 177580 106109 177581
rect 106043 177516 106044 177580
rect 106108 177516 106109 177580
rect 106043 177515 106109 177516
rect 106963 177580 107029 177581
rect 106963 177516 106964 177580
rect 107028 177516 107029 177580
rect 106963 177515 107029 177516
rect 104571 175404 104637 175405
rect 104571 175340 104572 175404
rect 104636 175340 104637 175404
rect 104571 175339 104637 175340
rect 104574 175130 104634 175339
rect 106046 175130 106106 177515
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 106106 175130
rect 106966 175130 107026 177515
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 108070 175130 108130 176699
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 114294 223954 114914 238000
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 110643 177988 110709 177989
rect 110643 177924 110644 177988
rect 110708 177924 110709 177988
rect 110643 177923 110709 177924
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177923
rect 112115 177580 112181 177581
rect 112115 177516 112116 177580
rect 112180 177516 112181 177580
rect 112115 177515 112181 177516
rect 114139 177580 114205 177581
rect 114139 177516 114140 177580
rect 114204 177516 114205 177580
rect 114139 177515 114205 177516
rect 112118 175130 112178 177515
rect 113219 177308 113285 177309
rect 113219 177244 113220 177308
rect 113284 177244 113285 177308
rect 113219 177243 113285 177244
rect 113222 175130 113282 177243
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114142 175130 114202 177515
rect 114294 176600 114914 187398
rect 118794 228454 119414 238000
rect 120582 235925 120642 284819
rect 121502 280941 121562 298691
rect 121499 280940 121565 280941
rect 121499 280876 121500 280940
rect 121564 280876 121565 280940
rect 121499 280875 121565 280876
rect 120763 269244 120829 269245
rect 120763 269180 120764 269244
rect 120828 269180 120829 269244
rect 120763 269179 120829 269180
rect 120766 238373 120826 269179
rect 123294 268954 123914 304398
rect 124811 299572 124877 299573
rect 124811 299508 124812 299572
rect 124876 299508 124877 299572
rect 124811 299507 124877 299508
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 120763 238372 120829 238373
rect 120763 238308 120764 238372
rect 120828 238308 120829 238372
rect 120763 238307 120829 238308
rect 120579 235924 120645 235925
rect 120579 235860 120580 235924
rect 120644 235860 120645 235924
rect 120579 235859 120645 235860
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 115795 177172 115861 177173
rect 115795 177108 115796 177172
rect 115860 177108 115861 177172
rect 115795 177107 115861 177108
rect 116899 177172 116965 177173
rect 116899 177108 116900 177172
rect 116964 177108 116965 177172
rect 116899 177107 116965 177108
rect 115798 175130 115858 177107
rect 114142 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 177107
rect 118371 176764 118437 176765
rect 118371 176700 118372 176764
rect 118436 176700 118437 176764
rect 118371 176699 118437 176700
rect 118374 175130 118434 176699
rect 118794 176600 119414 191898
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 120763 177580 120829 177581
rect 120763 177516 120764 177580
rect 120828 177516 120829 177580
rect 120763 177515 120829 177516
rect 122971 177580 123037 177581
rect 122971 177516 122972 177580
rect 123036 177516 123037 177580
rect 122971 177515 123037 177516
rect 120766 175130 120826 177515
rect 121867 175404 121933 175405
rect 121867 175340 121868 175404
rect 121932 175340 121933 175404
rect 121867 175339 121933 175340
rect 121870 175130 121930 175339
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 122974 175130 123034 177515
rect 123294 176600 123914 196398
rect 124814 185605 124874 299507
rect 125734 205597 125794 402187
rect 127794 381454 128414 403000
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 126099 292772 126165 292773
rect 126099 292708 126100 292772
rect 126164 292708 126165 292772
rect 126099 292707 126165 292708
rect 126102 283525 126162 292707
rect 126099 283524 126165 283525
rect 126099 283460 126100 283524
rect 126164 283460 126165 283524
rect 126099 283459 126165 283460
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 125731 205596 125797 205597
rect 125731 205532 125732 205596
rect 125796 205532 125797 205596
rect 125731 205531 125797 205532
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 124811 185604 124877 185605
rect 124811 185540 124812 185604
rect 124876 185540 124877 185604
rect 124811 185539 124877 185540
rect 127019 177580 127085 177581
rect 127019 177516 127020 177580
rect 127084 177516 127085 177580
rect 127019 177515 127085 177516
rect 124443 177172 124509 177173
rect 124443 177108 124444 177172
rect 124508 177108 124509 177172
rect 124443 177107 124509 177108
rect 124446 175130 124506 177107
rect 125731 176764 125797 176765
rect 125731 176700 125732 176764
rect 125796 176700 125797 176764
rect 125731 176699 125797 176700
rect 125734 175130 125794 176699
rect 127022 175130 127082 177515
rect 127794 176600 128414 200898
rect 132294 385954 132914 403000
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 130699 176764 130765 176765
rect 130699 176700 130700 176764
rect 130764 176700 130765 176764
rect 130699 176699 130765 176700
rect 131987 176764 132053 176765
rect 131987 176700 131988 176764
rect 132052 176700 132053 176764
rect 131987 176699 132053 176700
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 129411 175404 129477 175405
rect 129411 175340 129412 175404
rect 129476 175340 129477 175404
rect 129411 175339 129477 175340
rect 122974 175070 123132 175130
rect 118312 174494 118372 175070
rect 119397 174996 119463 174997
rect 119397 174932 119398 174996
rect 119462 174932 119463 174996
rect 119397 174931 119463 174932
rect 119400 174494 119460 174931
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 175339
rect 130702 175130 130762 176699
rect 129414 175070 129524 175130
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 131990 175130 132050 176699
rect 132294 176600 132914 205398
rect 136794 390454 137414 403000
rect 138611 401708 138677 401709
rect 138611 401644 138612 401708
rect 138676 401644 138677 401708
rect 138611 401643 138677 401644
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 138614 284885 138674 401643
rect 141294 394954 141914 403000
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 145794 399454 146414 403000
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 150294 367954 150914 403000
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 148179 366348 148245 366349
rect 148179 366284 148180 366348
rect 148244 366284 148245 366348
rect 148179 366283 148245 366284
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 142659 307868 142725 307869
rect 142659 307804 142660 307868
rect 142724 307804 142725 307868
rect 142659 307803 142725 307804
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 138611 284884 138677 284885
rect 138611 284820 138612 284884
rect 138676 284820 138677 284884
rect 138611 284819 138677 284820
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 135667 176764 135733 176765
rect 135667 176700 135668 176764
rect 135732 176700 135733 176764
rect 135667 176699 135733 176700
rect 133091 175404 133157 175405
rect 133091 175340 133092 175404
rect 133156 175340 133157 175404
rect 133091 175339 133157 175340
rect 133094 175130 133154 175339
rect 134382 175130 134442 176699
rect 131990 175070 132108 175130
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135670 175130 135730 176699
rect 136794 176600 137414 209898
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 142662 206957 142722 307803
rect 145794 291454 146414 326898
rect 146891 295356 146957 295357
rect 146891 295292 146892 295356
rect 146956 295292 146957 295356
rect 146891 295291 146957 295292
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 142659 206956 142725 206957
rect 142659 206892 142660 206956
rect 142724 206892 142725 206956
rect 142659 206891 142725 206892
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 176600 141914 178398
rect 145794 183454 146414 218898
rect 146894 187101 146954 295291
rect 148182 244357 148242 366283
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 149651 322964 149717 322965
rect 149651 322900 149652 322964
rect 149716 322900 149717 322964
rect 149651 322899 149717 322900
rect 148179 244356 148245 244357
rect 148179 244292 148180 244356
rect 148244 244292 148245 244356
rect 148179 244291 148245 244292
rect 146891 187100 146957 187101
rect 146891 187036 146892 187100
rect 146956 187036 146957 187100
rect 146891 187035 146957 187036
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149654 181525 149714 322899
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 149651 181524 149717 181525
rect 149651 181460 149652 181524
rect 149716 181460 149717 181524
rect 149651 181459 149717 181460
rect 148179 177172 148245 177173
rect 148179 177108 148180 177172
rect 148244 177108 148245 177172
rect 148179 177107 148245 177108
rect 148182 175130 148242 177107
rect 150294 176600 150914 187398
rect 154794 372454 155414 403000
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 159294 376954 159914 403000
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 157195 357508 157261 357509
rect 157195 357444 157196 357508
rect 157260 357444 157261 357508
rect 157195 357443 157261 357444
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 157198 199341 157258 357443
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 157379 287196 157445 287197
rect 157379 287132 157380 287196
rect 157444 287132 157445 287196
rect 157379 287131 157445 287132
rect 157382 240141 157442 287131
rect 159294 268954 159914 304398
rect 163794 381454 164414 403000
rect 166763 402252 166829 402253
rect 166763 402188 166764 402252
rect 166828 402188 166829 402252
rect 166763 402187 166829 402188
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 161979 302292 162045 302293
rect 161979 302228 161980 302292
rect 162044 302228 162045 302292
rect 161979 302227 162045 302228
rect 160691 292092 160757 292093
rect 160691 292028 160692 292092
rect 160756 292028 160757 292092
rect 160691 292027 160757 292028
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 157379 240140 157445 240141
rect 157379 240076 157380 240140
rect 157444 240076 157445 240140
rect 157379 240075 157445 240076
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 157195 199340 157261 199341
rect 157195 199276 157196 199340
rect 157260 199276 157261 199340
rect 157195 199275 157261 199276
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 176600 155414 191898
rect 159294 196954 159914 232398
rect 160694 217429 160754 292027
rect 161982 227085 162042 302227
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 166766 267750 166826 402187
rect 168294 385954 168914 403000
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 167683 289100 167749 289101
rect 167683 289036 167684 289100
rect 167748 289036 167749 289100
rect 167683 289035 167749 289036
rect 166766 267690 167010 267750
rect 166211 249116 166277 249117
rect 166211 249052 166212 249116
rect 166276 249052 166277 249116
rect 166211 249051 166277 249052
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 161979 227084 162045 227085
rect 161979 227020 161980 227084
rect 162044 227020 162045 227084
rect 161979 227019 162045 227020
rect 160691 217428 160757 217429
rect 160691 217364 160692 217428
rect 160756 217364 160757 217428
rect 160691 217363 160757 217364
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 159294 176600 159914 196398
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 166214 187237 166274 249051
rect 166950 248430 167010 267690
rect 166950 248370 167562 248430
rect 167502 246530 167562 248370
rect 166950 246470 167562 246530
rect 166950 246397 167010 246470
rect 166947 246396 167013 246397
rect 166947 246332 166948 246396
rect 167012 246332 167013 246396
rect 166947 246331 167013 246332
rect 166211 187236 166277 187237
rect 166211 187172 166212 187236
rect 166276 187172 166277 187236
rect 166211 187171 166277 187172
rect 166211 182204 166277 182205
rect 166211 182140 166212 182204
rect 166276 182140 166277 182204
rect 166211 182139 166277 182140
rect 135670 175070 135780 175130
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 166214 164389 166274 182139
rect 167502 178669 167562 246470
rect 167686 221509 167746 289035
rect 168294 277954 168914 313398
rect 172794 390454 173414 403000
rect 177067 395316 177133 395317
rect 177067 395252 177068 395316
rect 177132 395252 177133 395316
rect 177067 395251 177133 395252
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 175043 352204 175109 352205
rect 175043 352140 175044 352204
rect 175108 352140 175109 352204
rect 175043 352139 175109 352140
rect 174859 336700 174925 336701
rect 174859 336636 174860 336700
rect 174924 336636 174925 336700
rect 174859 336635 174925 336636
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 171731 294132 171797 294133
rect 171731 294068 171732 294132
rect 171796 294068 171797 294132
rect 171731 294067 171797 294068
rect 170259 293996 170325 293997
rect 170259 293932 170260 293996
rect 170324 293932 170325 293996
rect 170259 293931 170325 293932
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 167683 221508 167749 221509
rect 167683 221444 167684 221508
rect 167748 221444 167749 221508
rect 167683 221443 167749 221444
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 167499 178668 167565 178669
rect 167499 178604 167500 178668
rect 167564 178604 167565 178668
rect 167499 178603 167565 178604
rect 166395 178124 166461 178125
rect 166395 178060 166396 178124
rect 166460 178060 166461 178124
rect 166395 178059 166461 178060
rect 166211 164388 166277 164389
rect 166211 164324 166212 164388
rect 166276 164324 166277 164388
rect 166211 164323 166277 164324
rect 166398 161533 166458 178059
rect 167683 177036 167749 177037
rect 167683 176972 167684 177036
rect 167748 176972 167749 177036
rect 167683 176971 167749 176972
rect 167499 176900 167565 176901
rect 167499 176836 167500 176900
rect 167564 176836 167565 176900
rect 167499 176835 167565 176836
rect 166395 161532 166461 161533
rect 166395 161468 166396 161532
rect 166460 161468 166461 161532
rect 166395 161467 166461 161468
rect 167502 157453 167562 176835
rect 167686 157589 167746 176971
rect 168294 169954 168914 205398
rect 169707 184244 169773 184245
rect 169707 184180 169708 184244
rect 169772 184180 169773 184244
rect 169707 184179 169773 184180
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 167683 157588 167749 157589
rect 167683 157524 167684 157588
rect 167748 157524 167749 157588
rect 167683 157523 167749 157524
rect 167499 157452 167565 157453
rect 167499 157388 167500 157452
rect 167564 157388 167565 157452
rect 167499 157387 167565 157388
rect 69072 151954 69420 151986
rect 69072 151718 69128 151954
rect 69364 151718 69420 151954
rect 69072 151634 69420 151718
rect 69072 151398 69128 151634
rect 69364 151398 69420 151634
rect 69072 151366 69420 151398
rect 164136 151954 164484 151986
rect 164136 151718 164192 151954
rect 164428 151718 164484 151954
rect 164136 151634 164484 151718
rect 164136 151398 164192 151634
rect 164428 151398 164484 151634
rect 164136 151366 164484 151398
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 166211 143716 166277 143717
rect 166211 143652 166212 143716
rect 166276 143652 166277 143716
rect 166211 143651 166277 143652
rect 69072 115954 69420 115986
rect 69072 115718 69128 115954
rect 69364 115718 69420 115954
rect 69072 115634 69420 115718
rect 69072 115398 69128 115634
rect 69364 115398 69420 115634
rect 69072 115366 69420 115398
rect 164136 115954 164484 115986
rect 164136 115718 164192 115954
rect 164428 115718 164484 115954
rect 164136 115634 164484 115718
rect 164136 115398 164192 115634
rect 164428 115398 164484 115634
rect 164136 115366 164484 115398
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85682 94890
rect 86624 94830 86786 94890
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64643 13020 64709 13021
rect 64643 12956 64644 13020
rect 64708 12956 64709 13020
rect 64643 12955 64709 12956
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 70954 69914 93100
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 79954 78914 93100
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 84454 83414 93100
rect 84334 91221 84394 94830
rect 85622 91221 85682 94830
rect 86726 91221 86786 94830
rect 87094 94830 88044 94890
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 87094 92445 87154 94830
rect 87091 92444 87157 92445
rect 87091 92380 87092 92444
rect 87156 92380 87157 92444
rect 87091 92379 87157 92380
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 85619 91220 85685 91221
rect 85619 91156 85620 91220
rect 85684 91156 85685 91220
rect 85619 91155 85685 91156
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 88954 87914 93100
rect 88934 91221 88994 94830
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 91326 91221 91386 94830
rect 88931 91220 88997 91221
rect 88931 91156 88932 91220
rect 88996 91156 88997 91220
rect 88931 91155 88997 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91221 93962 94830
rect 94920 94757 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 96008 94830 96170 94890
rect 96688 94830 96906 94890
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 99136 94830 99298 94890
rect 99544 94830 99666 94890
rect 94917 94756 94983 94757
rect 94917 94692 94918 94756
rect 94982 94692 94983 94756
rect 94917 94691 94983 94692
rect 96110 91221 96170 94830
rect 96846 93870 96906 94830
rect 96846 93810 97090 93870
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 93899 91220 93965 91221
rect 93899 91156 93900 91220
rect 93964 91156 93965 91220
rect 93899 91155 93965 91156
rect 96107 91220 96173 91221
rect 96107 91156 96108 91220
rect 96172 91156 96173 91220
rect 96107 91155 96173 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 61954 96914 93100
rect 97030 91221 97090 93810
rect 97214 93533 97274 94830
rect 97211 93532 97277 93533
rect 97211 93468 97212 93532
rect 97276 93468 97277 93532
rect 97211 93467 97277 93468
rect 98134 92445 98194 94830
rect 98502 92445 98562 94830
rect 98131 92444 98197 92445
rect 98131 92380 98132 92444
rect 98196 92380 98197 92444
rect 98131 92379 98197 92380
rect 98499 92444 98565 92445
rect 98499 92380 98500 92444
rect 98564 92380 98565 92444
rect 98499 92379 98565 92380
rect 99238 91221 99298 94830
rect 99606 91765 99666 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 101690 94890
rect 99603 91764 99669 91765
rect 99603 91700 99604 91764
rect 99668 91700 99669 91764
rect 99603 91699 99669 91700
rect 100526 91221 100586 94830
rect 97027 91220 97093 91221
rect 97027 91156 97028 91220
rect 97092 91156 97093 91220
rect 97027 91155 97093 91156
rect 99235 91220 99301 91221
rect 99235 91156 99236 91220
rect 99300 91156 99301 91220
rect 99235 91155 99301 91156
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 66454 101414 93100
rect 101630 91221 101690 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 91357 101874 94830
rect 101811 91356 101877 91357
rect 101811 91292 101812 91356
rect 101876 91292 101877 91356
rect 101811 91291 101877 91292
rect 101998 91221 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 103216 94830 103346 94890
rect 102918 91221 102978 94830
rect 103286 91221 103346 94830
rect 104304 94754 104364 95200
rect 104206 94694 104364 94754
rect 104440 94754 104500 95200
rect 105392 94754 105452 95200
rect 104440 94694 104634 94754
rect 104206 91357 104266 94694
rect 104203 91356 104269 91357
rect 104203 91292 104204 91356
rect 104268 91292 104269 91356
rect 104203 91291 104269 91292
rect 104574 91221 104634 94694
rect 105126 94694 105452 94754
rect 105664 94754 105724 95200
rect 106480 94893 106540 95200
rect 106477 94892 106543 94893
rect 106477 94828 106478 94892
rect 106542 94828 106543 94892
rect 106477 94827 106543 94828
rect 106616 94754 106676 95200
rect 106779 94892 106845 94893
rect 106779 94828 106780 94892
rect 106844 94828 106845 94892
rect 106779 94827 106845 94828
rect 105664 94694 106106 94754
rect 105126 91221 105186 94694
rect 101627 91220 101693 91221
rect 101627 91156 101628 91220
rect 101692 91156 101693 91220
rect 101627 91155 101693 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 102915 91220 102981 91221
rect 102915 91156 102916 91220
rect 102980 91156 102981 91220
rect 102915 91155 102981 91156
rect 103283 91220 103349 91221
rect 103283 91156 103284 91220
rect 103348 91156 103349 91220
rect 103283 91155 103349 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105123 91220 105189 91221
rect 105123 91156 105124 91220
rect 105188 91156 105189 91220
rect 105123 91155 105189 91156
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 70954 105914 93100
rect 106046 91221 106106 94694
rect 106414 94694 106676 94754
rect 106414 91221 106474 94694
rect 106782 92445 106842 94827
rect 107704 94754 107764 95200
rect 108112 94754 108172 95200
rect 107702 94694 107764 94754
rect 108070 94694 108172 94754
rect 109064 94754 109124 95200
rect 109472 94754 109532 95200
rect 110152 94754 110212 95200
rect 110696 94754 110756 95200
rect 111240 94754 111300 95200
rect 109064 94694 109234 94754
rect 109472 94694 109602 94754
rect 106779 92444 106845 92445
rect 106779 92380 106780 92444
rect 106844 92380 106845 92444
rect 106779 92379 106845 92380
rect 107702 91357 107762 94694
rect 107699 91356 107765 91357
rect 107699 91292 107700 91356
rect 107764 91292 107765 91356
rect 107699 91291 107765 91292
rect 108070 91221 108130 94694
rect 109174 91629 109234 94694
rect 109171 91628 109237 91629
rect 109171 91564 109172 91628
rect 109236 91564 109237 91628
rect 109171 91563 109237 91564
rect 109542 91221 109602 94694
rect 110094 94694 110212 94754
rect 110646 94694 110756 94754
rect 111198 94694 111300 94754
rect 111920 94754 111980 95200
rect 112328 94754 112388 95200
rect 113144 94757 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113688 94830 113834 94890
rect 111920 94694 111994 94754
rect 110094 93261 110154 94694
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 106043 91220 106109 91221
rect 106043 91156 106044 91220
rect 106108 91156 106109 91220
rect 106043 91155 106109 91156
rect 106411 91220 106477 91221
rect 106411 91156 106412 91220
rect 106476 91156 106477 91220
rect 106411 91155 106477 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 75454 110414 93100
rect 110646 91221 110706 94694
rect 111198 91221 111258 94694
rect 111934 91221 111994 94694
rect 112302 94694 112388 94754
rect 113141 94756 113207 94757
rect 112302 91357 112362 94694
rect 113141 94692 113142 94756
rect 113206 94692 113207 94756
rect 113141 94691 113207 94692
rect 113774 93533 113834 94830
rect 114142 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 114776 94830 115122 94890
rect 113771 93532 113837 93533
rect 113771 93468 113772 93532
rect 113836 93468 113837 93532
rect 113771 93467 113837 93468
rect 114142 92309 114202 94830
rect 114139 92308 114205 92309
rect 114139 92244 114140 92308
rect 114204 92244 114205 92308
rect 114139 92243 114205 92244
rect 112299 91356 112365 91357
rect 112299 91292 112300 91356
rect 112364 91292 112365 91356
rect 112299 91291 112365 91292
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 79954 114914 93100
rect 115062 91221 115122 94830
rect 115430 94830 115516 94890
rect 115430 91221 115490 94830
rect 115864 94757 115924 95200
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115861 94756 115927 94757
rect 115861 94692 115862 94756
rect 115926 94692 115927 94756
rect 115861 94691 115927 94692
rect 116718 92445 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 92444 116781 92445
rect 116715 92380 116716 92444
rect 116780 92380 116781 92444
rect 116715 92379 116781 92380
rect 117086 91765 117146 94830
rect 117083 91764 117149 91765
rect 117083 91700 117084 91764
rect 117148 91700 117149 91764
rect 117083 91699 117149 91700
rect 118006 91221 118066 94830
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119906 94890
rect 119294 93870 119354 94830
rect 119294 93810 119722 93870
rect 115059 91220 115125 91221
rect 115059 91156 115060 91220
rect 115124 91156 115125 91220
rect 115059 91155 115125 91156
rect 115427 91220 115493 91221
rect 115427 91156 115428 91220
rect 115492 91156 115493 91220
rect 115427 91155 115493 91156
rect 118003 91220 118069 91221
rect 118003 91156 118004 91220
rect 118068 91156 118069 91220
rect 118003 91155 118069 91156
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 84454 119414 93100
rect 119662 92173 119722 93810
rect 119659 92172 119725 92173
rect 119659 92108 119660 92172
rect 119724 92108 119725 92172
rect 119659 92107 119725 92108
rect 119846 91221 119906 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 121984 94830 122114 94890
rect 120214 92445 120274 94830
rect 120211 92444 120277 92445
rect 120211 92380 120212 92444
rect 120276 92380 120277 92444
rect 120211 92379 120277 92380
rect 120582 91221 120642 94830
rect 121686 91221 121746 94830
rect 122054 91221 122114 94830
rect 122800 93870 122860 95200
rect 123208 94890 123268 95200
rect 122606 93810 122860 93870
rect 122974 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 122974 91221 123034 94830
rect 119843 91220 119909 91221
rect 119843 91156 119844 91220
rect 119908 91156 119909 91220
rect 119843 91155 119909 91156
rect 120579 91220 120645 91221
rect 120579 91156 120580 91220
rect 120644 91156 120645 91220
rect 120579 91155 120645 91156
rect 121683 91220 121749 91221
rect 121683 91156 121684 91220
rect 121748 91156 121749 91220
rect 121683 91155 121749 91156
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 122971 91220 123037 91221
rect 122971 91156 122972 91220
rect 123036 91156 123037 91220
rect 122971 91155 123037 91156
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 88954 123914 93100
rect 124078 92445 124138 94830
rect 124075 92444 124141 92445
rect 124075 92380 124076 92444
rect 124140 92380 124141 92444
rect 124075 92379 124141 92380
rect 124446 91357 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 125656 94830 125794 94890
rect 124443 91356 124509 91357
rect 124443 91292 124444 91356
rect 124508 91292 124509 91356
rect 124443 91291 124509 91292
rect 125366 91221 125426 94830
rect 125734 92445 125794 94830
rect 126472 94757 126532 95200
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 126608 94830 126714 94890
rect 128104 94830 128186 94890
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132050 94890
rect 126469 94756 126535 94757
rect 126469 94692 126470 94756
rect 126534 94692 126535 94756
rect 126469 94691 126535 94692
rect 125731 92444 125797 92445
rect 125731 92380 125732 92444
rect 125796 92380 125797 92444
rect 125731 92379 125797 92380
rect 126654 91221 126714 94830
rect 128126 93941 128186 94830
rect 128123 93940 128189 93941
rect 128123 93876 128124 93940
rect 128188 93876 128189 93940
rect 128123 93875 128189 93876
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 93100
rect 129414 92445 129474 94830
rect 130702 93669 130762 94830
rect 130699 93668 130765 93669
rect 130699 93604 130700 93668
rect 130764 93604 130765 93668
rect 130699 93603 130765 93604
rect 129411 92444 129477 92445
rect 129411 92380 129412 92444
rect 129476 92380 129477 92444
rect 129411 92379 129477 92380
rect 131990 91629 132050 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 135730 94890
rect 131987 91628 132053 91629
rect 131987 91564 131988 91628
rect 132052 91564 132053 91628
rect 131987 91563 132053 91564
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 93100
rect 133094 92445 133154 94830
rect 133091 92444 133157 92445
rect 133091 92380 133092 92444
rect 133156 92380 133157 92444
rect 133091 92379 133157 92380
rect 134382 91221 134442 94830
rect 135670 92445 135730 94830
rect 151310 94830 151556 94890
rect 135667 92444 135733 92445
rect 135667 92380 135668 92444
rect 135732 92380 135733 92444
rect 135667 92379 135733 92380
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 93100
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 70954 141914 93100
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 79954 150914 93100
rect 151310 91629 151370 94830
rect 151632 94754 151692 95200
rect 151768 94893 151828 95200
rect 151765 94892 151831 94893
rect 151765 94828 151766 94892
rect 151830 94828 151831 94892
rect 151765 94827 151831 94828
rect 151494 94694 151692 94754
rect 151904 94754 151964 95200
rect 151904 94694 152106 94754
rect 151494 92445 151554 94694
rect 152046 92445 152106 94694
rect 166214 93941 166274 143651
rect 167683 138140 167749 138141
rect 167683 138076 167684 138140
rect 167748 138076 167749 138140
rect 167683 138075 167749 138076
rect 166395 131476 166461 131477
rect 166395 131412 166396 131476
rect 166460 131412 166461 131476
rect 166395 131411 166461 131412
rect 166211 93940 166277 93941
rect 166211 93876 166212 93940
rect 166276 93876 166277 93940
rect 166211 93875 166277 93876
rect 151491 92444 151557 92445
rect 151491 92380 151492 92444
rect 151556 92380 151557 92444
rect 151491 92379 151557 92380
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 151307 91628 151373 91629
rect 151307 91564 151308 91628
rect 151372 91564 151373 91628
rect 151307 91563 151373 91564
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 84454 155414 93100
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 88954 159914 93100
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 93100
rect 166398 91085 166458 131411
rect 167499 129844 167565 129845
rect 167499 129780 167500 129844
rect 167564 129780 167565 129844
rect 167499 129779 167565 129780
rect 166395 91084 166461 91085
rect 166395 91020 166396 91084
rect 166460 91020 166461 91084
rect 166395 91019 166461 91020
rect 167502 80069 167562 129779
rect 167686 92173 167746 138075
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 169155 128484 169221 128485
rect 169155 128420 169156 128484
rect 169220 128420 169221 128484
rect 169155 128419 169221 128420
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 167683 92172 167749 92173
rect 167683 92108 167684 92172
rect 167748 92108 167749 92172
rect 167683 92107 167749 92108
rect 167499 80068 167565 80069
rect 167499 80004 167500 80068
rect 167564 80004 167565 80068
rect 167499 80003 167565 80004
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 97398
rect 169158 85509 169218 128419
rect 169155 85508 169221 85509
rect 169155 85444 169156 85508
rect 169220 85444 169221 85508
rect 169155 85443 169221 85444
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 169710 3365 169770 184179
rect 170262 92445 170322 293931
rect 171734 93805 171794 294067
rect 172794 282454 173414 317898
rect 173571 294268 173637 294269
rect 173571 294204 173572 294268
rect 173636 294204 173637 294268
rect 173571 294203 173637 294204
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 171915 262852 171981 262853
rect 171915 262788 171916 262852
rect 171980 262788 171981 262852
rect 171915 262787 171981 262788
rect 171918 235245 171978 262787
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 171915 235244 171981 235245
rect 171915 235180 171916 235244
rect 171980 235180 171981 235244
rect 171915 235179 171981 235180
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 171731 93804 171797 93805
rect 171731 93740 171732 93804
rect 171796 93740 171797 93804
rect 171731 93739 171797 93740
rect 170259 92444 170325 92445
rect 170259 92380 170260 92444
rect 170324 92380 170325 92444
rect 170259 92379 170325 92380
rect 172794 66454 173414 101898
rect 173574 93669 173634 294203
rect 173571 93668 173637 93669
rect 173571 93604 173572 93668
rect 173636 93604 173637 93668
rect 173571 93603 173637 93604
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 169707 3364 169773 3365
rect 169707 3300 169708 3364
rect 169772 3300 169773 3364
rect 169707 3299 169773 3300
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 174862 8261 174922 336635
rect 175046 21997 175106 352139
rect 176515 350028 176581 350029
rect 176515 349964 176516 350028
rect 176580 349964 176581 350028
rect 176515 349963 176581 349964
rect 176331 323644 176397 323645
rect 176331 323580 176332 323644
rect 176396 323580 176397 323644
rect 176331 323579 176397 323580
rect 176334 84829 176394 323579
rect 176331 84828 176397 84829
rect 176331 84764 176332 84828
rect 176396 84764 176397 84828
rect 176331 84763 176397 84764
rect 176518 28253 176578 349963
rect 177070 248301 177130 395251
rect 177294 394954 177914 403000
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 181794 399454 182414 403000
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 357154 182414 362898
rect 213294 394954 213914 403000
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 357154 213914 358398
rect 217794 399454 218414 403000
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 242942 398717 243002 470550
rect 246254 399941 246314 489363
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 246435 449308 246501 449309
rect 246435 449244 246436 449308
rect 246500 449244 246501 449308
rect 246435 449243 246501 449244
rect 246251 399940 246317 399941
rect 246251 399876 246252 399940
rect 246316 399876 246317 399940
rect 246251 399875 246317 399876
rect 246438 399805 246498 449243
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 246435 399804 246501 399805
rect 246435 399740 246436 399804
rect 246500 399740 246501 399804
rect 246435 399739 246501 399740
rect 242939 398716 243005 398717
rect 242939 398652 242940 398716
rect 243004 398652 243005 398716
rect 242939 398651 243005 398652
rect 246438 389877 246498 399739
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 246435 389876 246501 389877
rect 246435 389812 246436 389876
rect 246500 389812 246501 389876
rect 246435 389811 246501 389812
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 357154 218414 362898
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 357154 249914 358398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 357154 254414 362898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 357154 258914 367398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 357154 263414 371898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 357154 267914 376398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 357154 272414 380898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 357154 276914 385398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 357154 281414 389898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 357154 285914 358398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 295379 558244 295445 558245
rect 295379 558180 295380 558244
rect 295444 558180 295445 558244
rect 295379 558179 295445 558180
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 292619 525060 292685 525061
rect 292619 524996 292620 525060
rect 292684 524996 292685 525060
rect 292619 524995 292685 524996
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 292622 364350 292682 524995
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 295382 368661 295442 558179
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 301451 517580 301517 517581
rect 301451 517516 301452 517580
rect 301516 517516 301517 517580
rect 301451 517515 301517 517516
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 295563 389196 295629 389197
rect 295563 389132 295564 389196
rect 295628 389132 295629 389196
rect 295563 389131 295629 389132
rect 295379 368660 295445 368661
rect 295379 368596 295380 368660
rect 295444 368596 295445 368660
rect 295379 368595 295445 368596
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 292622 364290 293050 364350
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 357154 290414 362898
rect 291699 357644 291765 357645
rect 291699 357580 291700 357644
rect 291764 357580 291765 357644
rect 291699 357579 291765 357580
rect 291702 353290 291762 357579
rect 292619 353292 292685 353293
rect 292619 353290 292620 353292
rect 291702 353230 292620 353290
rect 292619 353228 292620 353230
rect 292684 353228 292685 353292
rect 292619 353227 292685 353228
rect 292990 335370 293050 364290
rect 294294 357154 294914 367398
rect 294091 356012 294157 356013
rect 294091 355948 294092 356012
rect 294156 355948 294157 356012
rect 294091 355947 294157 355948
rect 292622 335310 293050 335370
rect 199568 331954 199888 331986
rect 199568 331718 199610 331954
rect 199846 331718 199888 331954
rect 199568 331634 199888 331718
rect 199568 331398 199610 331634
rect 199846 331398 199888 331634
rect 199568 331366 199888 331398
rect 230288 331954 230608 331986
rect 230288 331718 230330 331954
rect 230566 331718 230608 331954
rect 230288 331634 230608 331718
rect 230288 331398 230330 331634
rect 230566 331398 230608 331634
rect 230288 331366 230608 331398
rect 261008 331954 261328 331986
rect 261008 331718 261050 331954
rect 261286 331718 261328 331954
rect 261008 331634 261328 331718
rect 261008 331398 261050 331634
rect 261286 331398 261328 331634
rect 261008 331366 261328 331398
rect 184208 327454 184528 327486
rect 184208 327218 184250 327454
rect 184486 327218 184528 327454
rect 184208 327134 184528 327218
rect 184208 326898 184250 327134
rect 184486 326898 184528 327134
rect 184208 326866 184528 326898
rect 214928 327454 215248 327486
rect 214928 327218 214970 327454
rect 215206 327218 215248 327454
rect 214928 327134 215248 327218
rect 214928 326898 214970 327134
rect 215206 326898 215248 327134
rect 214928 326866 215248 326898
rect 245648 327454 245968 327486
rect 245648 327218 245690 327454
rect 245926 327218 245968 327454
rect 245648 327134 245968 327218
rect 245648 326898 245690 327134
rect 245926 326898 245968 327134
rect 245648 326866 245968 326898
rect 276368 327454 276688 327486
rect 276368 327218 276410 327454
rect 276646 327218 276688 327454
rect 276368 327134 276688 327218
rect 276368 326898 276410 327134
rect 276646 326898 276688 327134
rect 276368 326866 276688 326898
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 179275 319020 179341 319021
rect 179275 318956 179276 319020
rect 179340 318956 179341 319020
rect 179275 318955 179341 318956
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 179091 263940 179157 263941
rect 179091 263876 179092 263940
rect 179156 263876 179157 263940
rect 179091 263875 179157 263876
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177067 248300 177133 248301
rect 177067 248236 177068 248300
rect 177132 248236 177133 248300
rect 177067 248235 177133 248236
rect 177070 65517 177130 248235
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 179094 86189 179154 263875
rect 179091 86188 179157 86189
rect 179091 86124 179092 86188
rect 179156 86124 179157 86188
rect 179091 86123 179157 86124
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177067 65516 177133 65517
rect 177067 65452 177068 65516
rect 177132 65452 177133 65516
rect 177067 65451 177133 65452
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 176515 28252 176581 28253
rect 176515 28188 176516 28252
rect 176580 28188 176581 28252
rect 176515 28187 176581 28188
rect 175043 21996 175109 21997
rect 175043 21932 175044 21996
rect 175108 21932 175109 21996
rect 175043 21931 175109 21932
rect 174859 8260 174925 8261
rect 174859 8196 174860 8260
rect 174924 8196 174925 8260
rect 174859 8195 174925 8196
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 -7066 177914 34398
rect 179278 15197 179338 318955
rect 292622 308685 292682 335310
rect 292619 308684 292685 308685
rect 292619 308620 292620 308684
rect 292684 308620 292685 308684
rect 292619 308619 292685 308620
rect 199568 295954 199888 295986
rect 199568 295718 199610 295954
rect 199846 295718 199888 295954
rect 199568 295634 199888 295718
rect 199568 295398 199610 295634
rect 199846 295398 199888 295634
rect 199568 295366 199888 295398
rect 230288 295954 230608 295986
rect 230288 295718 230330 295954
rect 230566 295718 230608 295954
rect 230288 295634 230608 295718
rect 230288 295398 230330 295634
rect 230566 295398 230608 295634
rect 230288 295366 230608 295398
rect 261008 295954 261328 295986
rect 261008 295718 261050 295954
rect 261286 295718 261328 295954
rect 261008 295634 261328 295718
rect 261008 295398 261050 295634
rect 261286 295398 261328 295634
rect 261008 295366 261328 295398
rect 184208 291454 184528 291486
rect 184208 291218 184250 291454
rect 184486 291218 184528 291454
rect 184208 291134 184528 291218
rect 184208 290898 184250 291134
rect 184486 290898 184528 291134
rect 184208 290866 184528 290898
rect 214928 291454 215248 291486
rect 214928 291218 214970 291454
rect 215206 291218 215248 291454
rect 214928 291134 215248 291218
rect 214928 290898 214970 291134
rect 215206 290898 215248 291134
rect 214928 290866 215248 290898
rect 245648 291454 245968 291486
rect 245648 291218 245690 291454
rect 245926 291218 245968 291454
rect 245648 291134 245968 291218
rect 245648 290898 245690 291134
rect 245926 290898 245968 291134
rect 245648 290866 245968 290898
rect 276368 291454 276688 291486
rect 276368 291218 276410 291454
rect 276646 291218 276688 291454
rect 276368 291134 276688 291218
rect 276368 290898 276410 291134
rect 276646 290898 276688 291134
rect 276368 290866 276688 290898
rect 293907 287196 293973 287197
rect 293907 287132 293908 287196
rect 293972 287132 293973 287196
rect 293907 287131 293973 287132
rect 199568 259954 199888 259986
rect 199568 259718 199610 259954
rect 199846 259718 199888 259954
rect 199568 259634 199888 259718
rect 199568 259398 199610 259634
rect 199846 259398 199888 259634
rect 199568 259366 199888 259398
rect 230288 259954 230608 259986
rect 230288 259718 230330 259954
rect 230566 259718 230608 259954
rect 230288 259634 230608 259718
rect 230288 259398 230330 259634
rect 230566 259398 230608 259634
rect 230288 259366 230608 259398
rect 261008 259954 261328 259986
rect 261008 259718 261050 259954
rect 261286 259718 261328 259954
rect 261008 259634 261328 259718
rect 261008 259398 261050 259634
rect 261286 259398 261328 259634
rect 261008 259366 261328 259398
rect 184208 255454 184528 255486
rect 184208 255218 184250 255454
rect 184486 255218 184528 255454
rect 184208 255134 184528 255218
rect 184208 254898 184250 255134
rect 184486 254898 184528 255134
rect 184208 254866 184528 254898
rect 214928 255454 215248 255486
rect 214928 255218 214970 255454
rect 215206 255218 215248 255454
rect 214928 255134 215248 255218
rect 214928 254898 214970 255134
rect 215206 254898 215248 255134
rect 214928 254866 215248 254898
rect 245648 255454 245968 255486
rect 245648 255218 245690 255454
rect 245926 255218 245968 255454
rect 245648 255134 245968 255218
rect 245648 254898 245690 255134
rect 245926 254898 245968 255134
rect 245648 254866 245968 254898
rect 276368 255454 276688 255486
rect 276368 255218 276410 255454
rect 276646 255218 276688 255454
rect 276368 255134 276688 255218
rect 276368 254898 276410 255134
rect 276646 254898 276688 255134
rect 276368 254866 276688 254898
rect 179459 244152 179525 244153
rect 179459 244088 179460 244152
rect 179524 244088 179525 244152
rect 179459 244087 179525 244088
rect 179275 15196 179341 15197
rect 179275 15132 179276 15196
rect 179340 15132 179341 15196
rect 179275 15131 179341 15132
rect 179462 5541 179522 244087
rect 179827 243540 179893 243541
rect 179827 243476 179828 243540
rect 179892 243476 179893 243540
rect 179827 243475 179893 243476
rect 179830 32469 179890 243475
rect 293171 243404 293237 243405
rect 293171 243340 293172 243404
rect 293236 243340 293237 243404
rect 293171 243339 293237 243340
rect 292619 242452 292685 242453
rect 292619 242450 292620 242452
rect 291886 242390 292620 242450
rect 291699 241228 291765 241229
rect 291699 241164 291700 241228
rect 291764 241164 291765 241228
rect 291699 241163 291765 241164
rect 289491 240820 289557 240821
rect 289491 240756 289492 240820
rect 289556 240756 289557 240820
rect 289491 240755 289557 240756
rect 181794 219454 182414 238000
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 179827 32468 179893 32469
rect 179827 32404 179828 32468
rect 179892 32404 179893 32468
rect 179827 32403 179893 32404
rect 179459 5540 179525 5541
rect 179459 5476 179460 5540
rect 179524 5476 179525 5540
rect 179459 5475 179525 5476
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 223954 186914 238000
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228454 191414 238000
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 232954 195914 238000
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 237454 200414 238000
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 238000
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 238000
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 238000
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 217794 219454 218414 238000
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 222294 223954 222914 238000
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 178000 222914 187398
rect 226794 228454 227414 238000
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 178000 227414 191898
rect 231294 232954 231914 238000
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 178000 231914 196398
rect 235794 237454 236414 238000
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 249294 214954 249914 238000
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 253794 219454 254414 238000
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 252507 185740 252573 185741
rect 252507 185676 252508 185740
rect 252572 185676 252573 185740
rect 252507 185675 252573 185676
rect 251219 181388 251285 181389
rect 251219 181324 251220 181388
rect 251284 181324 251285 181388
rect 251219 181323 251285 181324
rect 249011 178940 249077 178941
rect 249011 178876 249012 178940
rect 249076 178876 249077 178940
rect 249011 178875 249077 178876
rect 249014 174450 249074 178875
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 178000 249914 178398
rect 249747 177852 249813 177853
rect 249747 177788 249748 177852
rect 249812 177788 249813 177852
rect 249747 177787 249813 177788
rect 249195 177580 249261 177581
rect 249195 177516 249196 177580
rect 249260 177516 249261 177580
rect 249195 177515 249261 177516
rect 249198 174725 249258 177515
rect 249195 174724 249261 174725
rect 249195 174660 249196 174724
rect 249260 174660 249261 174724
rect 249195 174659 249261 174660
rect 249014 174390 249258 174450
rect 249198 172821 249258 174390
rect 249750 174317 249810 177787
rect 249747 174316 249813 174317
rect 249747 174252 249748 174316
rect 249812 174252 249813 174316
rect 249747 174251 249813 174252
rect 249195 172820 249261 172821
rect 249195 172756 249196 172820
rect 249260 172756 249261 172820
rect 249195 172755 249261 172756
rect 227874 151954 228194 151986
rect 227874 151718 227916 151954
rect 228152 151718 228194 151954
rect 227874 151634 228194 151718
rect 227874 151398 227916 151634
rect 228152 151398 228194 151634
rect 227874 151366 228194 151398
rect 237805 151954 238125 151986
rect 237805 151718 237847 151954
rect 238083 151718 238125 151954
rect 237805 151634 238125 151718
rect 237805 151398 237847 151634
rect 238083 151398 238125 151634
rect 237805 151366 238125 151398
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 251222 140861 251282 181323
rect 252510 173365 252570 185675
rect 253794 183454 254414 218898
rect 258294 223954 258914 238000
rect 259499 233884 259565 233885
rect 259499 233820 259500 233884
rect 259564 233820 259565 233884
rect 259499 233819 259565 233820
rect 259315 233204 259381 233205
rect 259315 233140 259316 233204
rect 259380 233140 259381 233204
rect 259315 233139 259381 233140
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 256739 217292 256805 217293
rect 256739 217228 256740 217292
rect 256804 217228 256805 217292
rect 256739 217227 256805 217228
rect 255267 214572 255333 214573
rect 255267 214508 255268 214572
rect 255332 214508 255333 214572
rect 255267 214507 255333 214508
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 252507 173364 252573 173365
rect 252507 173300 252508 173364
rect 252572 173300 252573 173364
rect 252507 173299 252573 173300
rect 251771 152964 251837 152965
rect 251771 152900 251772 152964
rect 251836 152900 251837 152964
rect 251771 152899 251837 152900
rect 251219 140860 251285 140861
rect 251219 140796 251220 140860
rect 251284 140796 251285 140860
rect 251219 140795 251285 140796
rect 251774 126309 251834 152899
rect 253794 147454 254414 182898
rect 254531 175948 254597 175949
rect 254531 175884 254532 175948
rect 254596 175884 254597 175948
rect 254531 175883 254597 175884
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 251771 126308 251837 126309
rect 251771 126244 251772 126308
rect 251836 126244 251837 126308
rect 251771 126243 251837 126244
rect 227874 115954 228194 115986
rect 227874 115718 227916 115954
rect 228152 115718 228194 115954
rect 227874 115634 228194 115718
rect 227874 115398 227916 115634
rect 228152 115398 228194 115634
rect 227874 115366 228194 115398
rect 237805 115954 238125 115986
rect 237805 115718 237847 115954
rect 238083 115718 238125 115954
rect 237805 115634 238125 115718
rect 237805 115398 237847 115634
rect 238083 115398 238125 115634
rect 237805 115366 238125 115398
rect 252507 113796 252573 113797
rect 252507 113732 252508 113796
rect 252572 113732 252573 113796
rect 252507 113731 252573 113732
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 242771 110866 243091 110898
rect 252510 110805 252570 113731
rect 253794 111454 254414 146898
rect 254534 136645 254594 175883
rect 255270 140453 255330 214507
rect 255451 184380 255517 184381
rect 255451 184316 255452 184380
rect 255516 184316 255517 184380
rect 255451 184315 255517 184316
rect 255454 157317 255514 184315
rect 256742 158813 256802 217227
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 256923 180164 256989 180165
rect 256923 180100 256924 180164
rect 256988 180100 256989 180164
rect 256923 180099 256989 180100
rect 256739 158812 256805 158813
rect 256739 158748 256740 158812
rect 256804 158748 256805 158812
rect 256739 158747 256805 158748
rect 255451 157316 255517 157317
rect 255451 157252 255452 157316
rect 255516 157252 255517 157316
rect 255451 157251 255517 157252
rect 255267 140452 255333 140453
rect 255267 140388 255268 140452
rect 255332 140388 255333 140452
rect 255267 140387 255333 140388
rect 256926 139909 256986 180099
rect 258294 151954 258914 187398
rect 259318 160717 259378 233139
rect 259315 160716 259381 160717
rect 259315 160652 259316 160716
rect 259380 160652 259381 160716
rect 259315 160651 259381 160652
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 256923 139908 256989 139909
rect 256923 139844 256924 139908
rect 256988 139844 256989 139908
rect 256923 139843 256989 139844
rect 254531 136644 254597 136645
rect 254531 136580 254532 136644
rect 254596 136580 254597 136644
rect 254531 136579 254597 136580
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 252507 110804 252573 110805
rect 252507 110740 252508 110804
rect 252572 110740 252573 110804
rect 252507 110739 252573 110740
rect 251219 109172 251285 109173
rect 251219 109108 251220 109172
rect 251284 109108 251285 109172
rect 251219 109107 251285 109108
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 79954 222914 94000
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 84454 227414 94000
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 88954 231914 94000
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 61954 240914 94000
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 66454 245414 94000
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 70954 249914 94000
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 251222 3501 251282 109107
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 251219 3500 251285 3501
rect 251219 3436 251220 3500
rect 251284 3436 251285 3500
rect 251219 3435 251285 3436
rect 253794 3454 254414 38898
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 115954 258914 151398
rect 259502 149701 259562 233819
rect 262794 228454 263414 238000
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 261339 210356 261405 210357
rect 261339 210292 261340 210356
rect 261404 210292 261405 210356
rect 261339 210291 261405 210292
rect 259683 195260 259749 195261
rect 259683 195196 259684 195260
rect 259748 195196 259749 195260
rect 259683 195195 259749 195196
rect 259686 170101 259746 195195
rect 260971 176628 261037 176629
rect 260971 176564 260972 176628
rect 261036 176564 261037 176628
rect 260971 176563 261037 176564
rect 259683 170100 259749 170101
rect 259683 170036 259684 170100
rect 259748 170036 259749 170100
rect 259683 170035 259749 170036
rect 260974 152693 261034 176563
rect 260971 152692 261037 152693
rect 260971 152628 260972 152692
rect 261036 152628 261037 152692
rect 260971 152627 261037 152628
rect 259499 149700 259565 149701
rect 259499 149636 259500 149700
rect 259564 149636 259565 149700
rect 259499 149635 259565 149636
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 261342 95437 261402 210291
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262259 186964 262325 186965
rect 262259 186900 262260 186964
rect 262324 186900 262325 186964
rect 262259 186899 262325 186900
rect 262262 141813 262322 186899
rect 262794 156454 263414 191898
rect 267294 232954 267914 238000
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 271794 237454 272414 238000
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271091 232116 271157 232117
rect 271091 232052 271092 232116
rect 271156 232052 271157 232116
rect 271091 232051 271157 232052
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 263547 189684 263613 189685
rect 263547 189620 263548 189684
rect 263612 189620 263613 189684
rect 263547 189619 263613 189620
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262259 141812 262325 141813
rect 262259 141748 262260 141812
rect 262324 141748 262325 141812
rect 262259 141747 262325 141748
rect 262794 120454 263414 155898
rect 263550 142221 263610 189619
rect 263731 181660 263797 181661
rect 263731 181596 263732 181660
rect 263796 181596 263797 181660
rect 263731 181595 263797 181596
rect 263734 163981 263794 181595
rect 265019 175948 265085 175949
rect 265019 175884 265020 175948
rect 265084 175884 265085 175948
rect 265019 175883 265085 175884
rect 263731 163980 263797 163981
rect 263731 163916 263732 163980
rect 263796 163916 263797 163980
rect 263731 163915 263797 163916
rect 265022 142629 265082 175883
rect 265571 174588 265637 174589
rect 265571 174524 265572 174588
rect 265636 174524 265637 174588
rect 265571 174523 265637 174524
rect 265019 142628 265085 142629
rect 265019 142564 265020 142628
rect 265084 142564 265085 142628
rect 265019 142563 265085 142564
rect 263547 142220 263613 142221
rect 263547 142156 263548 142220
rect 263612 142156 263613 142220
rect 263547 142155 263613 142156
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 261339 95436 261405 95437
rect 261339 95372 261340 95436
rect 261404 95372 261405 95436
rect 261339 95371 261405 95372
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 265574 3501 265634 174523
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 269067 160716 269133 160717
rect 269067 160652 269068 160716
rect 269132 160652 269133 160716
rect 269067 160651 269133 160652
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 269070 60077 269130 160651
rect 269067 60076 269133 60077
rect 269067 60012 269068 60076
rect 269132 60012 269133 60076
rect 269067 60011 269133 60012
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 265571 3500 265637 3501
rect 265571 3436 265572 3500
rect 265636 3436 265637 3500
rect 265571 3435 265637 3436
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 -3226 267914 16398
rect 269070 11797 269130 60011
rect 271094 46885 271154 232051
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271091 46884 271157 46885
rect 271091 46820 271092 46884
rect 271156 46820 271157 46884
rect 271091 46819 271157 46820
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 269067 11796 269133 11797
rect 269067 11732 269068 11796
rect 269132 11732 269133 11796
rect 269067 11731 269133 11732
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 205954 276914 238000
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 238000
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 238000
rect 288203 231300 288269 231301
rect 288203 231236 288204 231300
rect 288268 231236 288269 231300
rect 288203 231235 288269 231236
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 288206 100061 288266 231235
rect 288203 100060 288269 100061
rect 288203 99996 288204 100060
rect 288268 99996 288269 100060
rect 288203 99995 288269 99996
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 289494 19277 289554 240755
rect 289794 219454 290414 238000
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 291702 113933 291762 241163
rect 291886 231165 291946 242390
rect 292619 242388 292620 242390
rect 292684 242388 292685 242452
rect 292619 242387 292685 242388
rect 293174 240549 293234 243339
rect 292619 240548 292685 240549
rect 292619 240484 292620 240548
rect 292684 240484 292685 240548
rect 292619 240483 292685 240484
rect 293171 240548 293237 240549
rect 293171 240484 293172 240548
rect 293236 240484 293237 240548
rect 293171 240483 293237 240484
rect 291883 231164 291949 231165
rect 291883 231100 291884 231164
rect 291948 231100 291949 231164
rect 291883 231099 291949 231100
rect 292622 198117 292682 240483
rect 292619 198116 292685 198117
rect 292619 198052 292620 198116
rect 292684 198052 292685 198116
rect 292619 198051 292685 198052
rect 292622 144125 292682 198051
rect 293910 149701 293970 287131
rect 294094 242453 294154 355947
rect 295382 334389 295442 368595
rect 295566 336701 295626 389131
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 297955 358052 298021 358053
rect 297955 357988 297956 358052
rect 298020 357988 298021 358052
rect 297955 357987 298021 357988
rect 297958 355061 298018 357987
rect 297403 355060 297469 355061
rect 297403 354996 297404 355060
rect 297468 354996 297469 355060
rect 297403 354995 297469 354996
rect 297955 355060 298021 355061
rect 297955 354996 297956 355060
rect 298020 354996 298021 355060
rect 297955 354995 298021 354996
rect 295563 336700 295629 336701
rect 295563 336636 295564 336700
rect 295628 336636 295629 336700
rect 295563 336635 295629 336636
rect 295931 336700 295997 336701
rect 295931 336636 295932 336700
rect 295996 336636 295997 336700
rect 295931 336635 295997 336636
rect 295379 334388 295445 334389
rect 295379 334324 295380 334388
rect 295444 334324 295445 334388
rect 295379 334323 295445 334324
rect 295934 286381 295994 336635
rect 296115 327724 296181 327725
rect 296115 327660 296116 327724
rect 296180 327660 296181 327724
rect 296115 327659 296181 327660
rect 296118 287197 296178 327659
rect 296115 287196 296181 287197
rect 296115 287132 296116 287196
rect 296180 287132 296181 287196
rect 296115 287131 296181 287132
rect 295931 286380 295997 286381
rect 295931 286316 295932 286380
rect 295996 286316 295997 286380
rect 295931 286315 295997 286316
rect 297219 278900 297285 278901
rect 297219 278836 297220 278900
rect 297284 278836 297285 278900
rect 297219 278835 297285 278836
rect 295931 270468 295997 270469
rect 295931 270404 295932 270468
rect 295996 270404 295997 270468
rect 295931 270403 295997 270404
rect 295379 263532 295445 263533
rect 295379 263468 295380 263532
rect 295444 263468 295445 263532
rect 295379 263467 295445 263468
rect 294091 242452 294157 242453
rect 294091 242388 294092 242452
rect 294156 242388 294157 242452
rect 294091 242387 294157 242388
rect 294294 223954 294914 238000
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 293907 149700 293973 149701
rect 293907 149636 293908 149700
rect 293972 149636 293973 149700
rect 293907 149635 293973 149636
rect 292619 144124 292685 144125
rect 292619 144060 292620 144124
rect 292684 144060 292685 144124
rect 292619 144059 292685 144060
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 291699 113932 291765 113933
rect 291699 113868 291700 113932
rect 291764 113868 291765 113932
rect 291699 113867 291765 113868
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289491 19276 289557 19277
rect 289491 19212 289492 19276
rect 289556 19212 289557 19276
rect 289491 19211 289557 19212
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 79954 294914 115398
rect 295382 84285 295442 263467
rect 295934 202197 295994 270403
rect 295931 202196 295997 202197
rect 295931 202132 295932 202196
rect 295996 202132 295997 202196
rect 295931 202131 295997 202132
rect 295379 84284 295445 84285
rect 295379 84220 295380 84284
rect 295444 84220 295445 84284
rect 295379 84219 295445 84220
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 297222 11797 297282 278835
rect 297406 246261 297466 354995
rect 298794 336454 299414 371898
rect 299611 360908 299677 360909
rect 299611 360844 299612 360908
rect 299676 360844 299677 360908
rect 299611 360843 299677 360844
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 297403 246260 297469 246261
rect 297403 246196 297404 246260
rect 297468 246196 297469 246260
rect 297403 246195 297469 246196
rect 298794 228454 299414 263898
rect 299614 237013 299674 360843
rect 299611 237012 299677 237013
rect 299611 236948 299612 237012
rect 299676 236948 299677 237012
rect 299611 236947 299677 236948
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 301454 220829 301514 517515
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 311019 596460 311085 596461
rect 311019 596396 311020 596460
rect 311084 596396 311085 596460
rect 311019 596395 311085 596396
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 305499 357916 305565 357917
rect 305499 357852 305500 357916
rect 305564 357852 305565 357916
rect 305499 357851 305565 357852
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 301451 220828 301517 220829
rect 301451 220764 301452 220828
rect 301516 220764 301517 220828
rect 301451 220763 301517 220764
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 301635 128484 301701 128485
rect 301635 128420 301636 128484
rect 301700 128420 301701 128484
rect 301635 128419 301701 128420
rect 301451 126444 301517 126445
rect 301451 126380 301452 126444
rect 301516 126380 301517 126444
rect 301451 126379 301517 126380
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 299979 112708 300045 112709
rect 299979 112644 299980 112708
rect 300044 112644 300045 112708
rect 299979 112643 300045 112644
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 299982 24173 300042 112643
rect 299979 24172 300045 24173
rect 299979 24108 299980 24172
rect 300044 24108 300045 24172
rect 299979 24107 300045 24108
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 297219 11796 297285 11797
rect 297219 11732 297220 11796
rect 297284 11732 297285 11796
rect 297219 11731 297285 11732
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 -2266 299414 11898
rect 301454 10301 301514 126379
rect 301638 68237 301698 128419
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 304211 99788 304277 99789
rect 304211 99724 304212 99788
rect 304276 99724 304277 99788
rect 304211 99723 304277 99724
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 301635 68236 301701 68237
rect 301635 68172 301636 68236
rect 301700 68172 301701 68236
rect 301635 68171 301701 68172
rect 303294 52954 303914 88398
rect 304214 72453 304274 99723
rect 305502 91765 305562 357851
rect 307794 345454 308414 380898
rect 309179 369884 309245 369885
rect 309179 369820 309180 369884
rect 309244 369820 309245 369884
rect 309179 369819 309245 369820
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 309182 218653 309242 369819
rect 311022 233069 311082 596395
rect 312294 565954 312914 601398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 313779 597820 313845 597821
rect 313779 597756 313780 597820
rect 313844 597756 313845 597820
rect 313779 597755 313845 597756
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 311019 233068 311085 233069
rect 311019 233004 311020 233068
rect 311084 233004 311085 233068
rect 311019 233003 311085 233004
rect 309179 218652 309245 218653
rect 309179 218588 309180 218652
rect 309244 218588 309245 218652
rect 309179 218587 309245 218588
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 178000 308414 200898
rect 312294 205954 312914 241398
rect 313782 225589 313842 597755
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 318011 462364 318077 462365
rect 318011 462300 318012 462364
rect 318076 462300 318077 462364
rect 318011 462299 318077 462300
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 313779 225588 313845 225589
rect 313779 225524 313780 225588
rect 313844 225524 313845 225588
rect 313779 225523 313845 225524
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 178000 312914 205398
rect 316794 210454 317414 245898
rect 318014 232525 318074 462299
rect 321294 430954 321914 466398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 324267 464404 324333 464405
rect 324267 464340 324268 464404
rect 324332 464340 324333 464404
rect 324267 464339 324333 464340
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 318011 232524 318077 232525
rect 318011 232460 318012 232524
rect 318076 232460 318077 232524
rect 318011 232459 318077 232460
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 178000 317414 209898
rect 321294 214954 321914 250398
rect 322979 230484 323045 230485
rect 322979 230420 322980 230484
rect 323044 230420 323045 230484
rect 322979 230419 323045 230420
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 320219 192540 320285 192541
rect 320219 192476 320220 192540
rect 320284 192476 320285 192540
rect 320219 192475 320285 192476
rect 320222 174450 320282 192475
rect 321294 178954 321914 214398
rect 322059 192676 322125 192677
rect 322059 192612 322060 192676
rect 322124 192612 322125 192676
rect 322059 192611 322125 192612
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 178000 321914 178398
rect 321323 174452 321389 174453
rect 321323 174450 321324 174452
rect 320222 174390 321324 174450
rect 321323 174388 321324 174390
rect 321388 174388 321389 174452
rect 321323 174387 321389 174388
rect 314208 151954 314528 151986
rect 314208 151718 314250 151954
rect 314486 151718 314528 151954
rect 314208 151634 314528 151718
rect 314208 151398 314250 151634
rect 314486 151398 314528 151634
rect 314208 151366 314528 151398
rect 317472 151954 317792 151986
rect 317472 151718 317514 151954
rect 317750 151718 317792 151954
rect 317472 151634 317792 151718
rect 317472 151398 317514 151634
rect 317750 151398 317792 151634
rect 317472 151366 317792 151398
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 307339 141676 307405 141677
rect 307339 141612 307340 141676
rect 307404 141612 307405 141676
rect 307339 141611 307405 141612
rect 307155 137052 307221 137053
rect 307155 136988 307156 137052
rect 307220 136988 307221 137052
rect 307155 136987 307221 136988
rect 305683 113660 305749 113661
rect 305683 113596 305684 113660
rect 305748 113596 305749 113660
rect 305683 113595 305749 113596
rect 305499 91764 305565 91765
rect 305499 91700 305500 91764
rect 305564 91700 305565 91764
rect 305499 91699 305565 91700
rect 304211 72452 304277 72453
rect 304211 72388 304212 72452
rect 304276 72388 304277 72452
rect 304211 72387 304277 72388
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 305686 29613 305746 113595
rect 306971 97884 307037 97885
rect 306971 97820 306972 97884
rect 307036 97820 307037 97884
rect 306971 97819 307037 97820
rect 305683 29612 305749 29613
rect 305683 29548 305684 29612
rect 305748 29548 305749 29612
rect 305683 29547 305749 29548
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 301451 10300 301517 10301
rect 301451 10236 301452 10300
rect 301516 10236 301517 10300
rect 301451 10235 301517 10236
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 -3226 303914 16398
rect 306974 2685 307034 97819
rect 307158 89045 307218 136987
rect 307342 134469 307402 141611
rect 307339 134468 307405 134469
rect 307339 134404 307340 134468
rect 307404 134404 307405 134468
rect 307339 134403 307405 134404
rect 314208 115954 314528 115986
rect 314208 115718 314250 115954
rect 314486 115718 314528 115954
rect 314208 115634 314528 115718
rect 314208 115398 314250 115634
rect 314486 115398 314528 115634
rect 314208 115366 314528 115398
rect 317472 115954 317792 115986
rect 317472 115718 317514 115954
rect 317750 115718 317792 115954
rect 317472 115634 317792 115718
rect 317472 115398 317514 115634
rect 317750 115398 317792 115634
rect 317472 115366 317792 115398
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 322062 108357 322122 192611
rect 322982 125493 323042 230419
rect 324270 229110 324330 464339
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 324270 229050 324882 229110
rect 324822 217973 324882 229050
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 324819 217972 324885 217973
rect 324819 217908 324820 217972
rect 324884 217908 324885 217972
rect 324819 217907 324885 217908
rect 323163 207092 323229 207093
rect 323163 207028 323164 207092
rect 323228 207028 323229 207092
rect 323163 207027 323229 207028
rect 322979 125492 323045 125493
rect 322979 125428 322980 125492
rect 323044 125428 323045 125492
rect 322979 125427 323045 125428
rect 323166 117061 323226 207027
rect 324822 196621 324882 217907
rect 324819 196620 324885 196621
rect 324819 196556 324820 196620
rect 324884 196556 324885 196620
rect 324819 196555 324885 196556
rect 325794 183454 326414 218898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 336043 604484 336109 604485
rect 336043 604420 336044 604484
rect 336108 604420 336109 604484
rect 336043 604419 336109 604420
rect 335859 600404 335925 600405
rect 335859 600340 335860 600404
rect 335924 600340 335925 600404
rect 335859 600339 335925 600340
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 333099 565860 333165 565861
rect 333099 565796 333100 565860
rect 333164 565796 333165 565860
rect 333099 565795 333165 565796
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 331811 546548 331877 546549
rect 331811 546484 331812 546548
rect 331876 546484 331877 546548
rect 331811 546483 331877 546484
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 329787 209812 329853 209813
rect 329787 209748 329788 209812
rect 329852 209748 329853 209812
rect 329787 209747 329853 209748
rect 328683 184244 328749 184245
rect 328683 184180 328684 184244
rect 328748 184180 328749 184244
rect 328683 184179 328749 184180
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 327027 182884 327093 182885
rect 327027 182820 327028 182884
rect 327092 182820 327093 182884
rect 327027 182819 327093 182820
rect 326659 178804 326725 178805
rect 326659 178740 326660 178804
rect 326724 178740 326725 178804
rect 326659 178739 326725 178740
rect 326662 173229 326722 178739
rect 326659 173228 326725 173229
rect 326659 173164 326660 173228
rect 326724 173164 326725 173228
rect 326659 173163 326725 173164
rect 327030 166293 327090 182819
rect 328499 178940 328565 178941
rect 328499 178876 328500 178940
rect 328564 178876 328565 178940
rect 328499 178875 328565 178876
rect 327211 176220 327277 176221
rect 327211 176156 327212 176220
rect 327276 176156 327277 176220
rect 327211 176155 327277 176156
rect 327214 170917 327274 176155
rect 327211 170916 327277 170917
rect 327211 170852 327212 170916
rect 327276 170852 327277 170916
rect 327211 170851 327277 170852
rect 327027 166292 327093 166293
rect 327027 166228 327028 166292
rect 327092 166228 327093 166292
rect 327027 166227 327093 166228
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 323163 117060 323229 117061
rect 323163 116996 323164 117060
rect 323228 116996 323229 117060
rect 323163 116995 323229 116996
rect 325794 111454 326414 146898
rect 328502 138685 328562 178875
rect 328686 161805 328746 184179
rect 328683 161804 328749 161805
rect 328683 161740 328684 161804
rect 328748 161740 328749 161804
rect 328683 161739 328749 161740
rect 329051 151060 329117 151061
rect 329051 150996 329052 151060
rect 329116 150996 329117 151060
rect 329051 150995 329117 150996
rect 328499 138684 328565 138685
rect 328499 138620 328500 138684
rect 328564 138620 328565 138684
rect 328499 138619 328565 138620
rect 329054 123045 329114 150995
rect 329051 123044 329117 123045
rect 329051 122980 329052 123044
rect 329116 122980 329117 123044
rect 329051 122979 329117 122980
rect 329790 114613 329850 209747
rect 330294 187954 330914 223398
rect 331814 200021 331874 546483
rect 331811 200020 331877 200021
rect 331811 199956 331812 200020
rect 331876 199956 331877 200020
rect 331811 199955 331877 199956
rect 331814 198797 331874 199955
rect 331811 198796 331877 198797
rect 331811 198732 331812 198796
rect 331876 198732 331877 198796
rect 331811 198731 331877 198732
rect 332547 196076 332613 196077
rect 332547 196012 332548 196076
rect 332612 196012 332613 196076
rect 332547 196011 332613 196012
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 331259 181388 331325 181389
rect 331259 181324 331260 181388
rect 331324 181324 331325 181388
rect 331259 181323 331325 181324
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 329787 114612 329853 114613
rect 329787 114548 329788 114612
rect 329852 114548 329853 114612
rect 329787 114547 329853 114548
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 324267 108628 324333 108629
rect 324267 108564 324268 108628
rect 324332 108564 324333 108628
rect 324267 108563 324333 108564
rect 322059 108356 322125 108357
rect 322059 108292 322060 108356
rect 322124 108292 322125 108356
rect 322059 108291 322125 108292
rect 324270 95165 324330 108563
rect 324267 95164 324333 95165
rect 324267 95100 324268 95164
rect 324332 95100 324333 95164
rect 324267 95099 324333 95100
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307155 89044 307221 89045
rect 307155 88980 307156 89044
rect 307220 88980 307221 89044
rect 307155 88979 307221 88980
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 306971 2684 307037 2685
rect 306971 2620 306972 2684
rect 307036 2620 307037 2684
rect 306971 2619 307037 2620
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 61954 312914 94000
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 66454 317414 94000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 70954 321914 94000
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 79954 330914 115398
rect 331262 111893 331322 181323
rect 331443 177444 331509 177445
rect 331443 177380 331444 177444
rect 331508 177380 331509 177444
rect 331443 177379 331509 177380
rect 331446 131341 331506 177379
rect 331443 131340 331509 131341
rect 331443 131276 331444 131340
rect 331508 131276 331509 131340
rect 331443 131275 331509 131276
rect 331259 111892 331325 111893
rect 331259 111828 331260 111892
rect 331324 111828 331325 111892
rect 331259 111827 331325 111828
rect 332550 98157 332610 196011
rect 332547 98156 332613 98157
rect 332547 98092 332548 98156
rect 332612 98092 332613 98156
rect 332547 98091 332613 98092
rect 333102 95709 333162 565795
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 335862 503029 335922 600339
rect 336046 522341 336106 604419
rect 337331 603124 337397 603125
rect 337331 603060 337332 603124
rect 337396 603060 337397 603124
rect 337331 603059 337397 603060
rect 337334 582997 337394 603059
rect 339294 597438 339914 628398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 340091 603260 340157 603261
rect 340091 603196 340092 603260
rect 340156 603196 340157 603260
rect 340091 603195 340157 603196
rect 338619 596324 338685 596325
rect 338619 596260 338620 596324
rect 338684 596260 338685 596324
rect 338619 596259 338685 596260
rect 337515 584084 337581 584085
rect 337515 584020 337516 584084
rect 337580 584020 337581 584084
rect 337515 584019 337581 584020
rect 337331 582996 337397 582997
rect 337331 582932 337332 582996
rect 337396 582932 337397 582996
rect 337331 582931 337397 582932
rect 337331 528596 337397 528597
rect 337331 528532 337332 528596
rect 337396 528532 337397 528596
rect 337331 528531 337397 528532
rect 336043 522340 336109 522341
rect 336043 522276 336044 522340
rect 336108 522276 336109 522340
rect 336043 522275 336109 522276
rect 335859 503028 335925 503029
rect 335859 502964 335860 503028
rect 335924 502964 335925 503028
rect 335859 502963 335925 502964
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 335859 415036 335925 415037
rect 335859 414972 335860 415036
rect 335924 414972 335925 415036
rect 335859 414971 335925 414972
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334019 205732 334085 205733
rect 334019 205668 334020 205732
rect 334084 205668 334085 205732
rect 334019 205667 334085 205668
rect 334022 111077 334082 205667
rect 334794 192454 335414 227898
rect 335675 196076 335741 196077
rect 335675 196012 335676 196076
rect 335740 196012 335741 196076
rect 335675 196011 335741 196012
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 335678 180810 335738 196011
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 335494 180750 335738 180810
rect 335494 132510 335554 180750
rect 335862 167109 335922 414971
rect 337334 373285 337394 528531
rect 337518 508197 337578 584019
rect 338622 540293 338682 596259
rect 338619 540292 338685 540293
rect 338619 540228 338620 540292
rect 338684 540228 338685 540292
rect 338619 540227 338685 540228
rect 337515 508196 337581 508197
rect 337515 508132 337516 508196
rect 337580 508132 337581 508196
rect 337515 508131 337581 508132
rect 338987 483036 339053 483037
rect 338987 482972 338988 483036
rect 339052 482972 339053 483036
rect 338987 482971 339053 482972
rect 337515 419796 337581 419797
rect 337515 419732 337516 419796
rect 337580 419732 337581 419796
rect 337515 419731 337581 419732
rect 337331 373284 337397 373285
rect 337331 373220 337332 373284
rect 337396 373220 337397 373284
rect 337331 373219 337397 373220
rect 337518 371925 337578 419731
rect 338990 395453 339050 482971
rect 339171 442916 339237 442917
rect 339171 442852 339172 442916
rect 339236 442852 339237 442916
rect 339171 442851 339237 442852
rect 339174 398853 339234 442851
rect 339171 398852 339237 398853
rect 339171 398788 339172 398852
rect 339236 398788 339237 398852
rect 339171 398787 339237 398788
rect 338987 395452 339053 395453
rect 338987 395388 338988 395452
rect 339052 395388 339053 395452
rect 338987 395387 339053 395388
rect 339294 376954 339914 398000
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 337515 371924 337581 371925
rect 337515 371860 337516 371924
rect 337580 371860 337581 371924
rect 337515 371859 337581 371860
rect 336779 358868 336845 358869
rect 336779 358804 336780 358868
rect 336844 358804 336845 358868
rect 336779 358803 336845 358804
rect 335859 167108 335925 167109
rect 335859 167044 335860 167108
rect 335924 167044 335925 167108
rect 335859 167043 335925 167044
rect 335494 132450 335738 132510
rect 335678 122909 335738 132450
rect 335675 122908 335741 122909
rect 335675 122844 335676 122908
rect 335740 122844 335741 122908
rect 335675 122843 335741 122844
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334019 111076 334085 111077
rect 334019 111012 334020 111076
rect 334084 111012 334085 111076
rect 334019 111011 334085 111012
rect 333099 95708 333165 95709
rect 333099 95644 333100 95708
rect 333164 95644 333165 95708
rect 333099 95643 333165 95644
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 336782 26213 336842 358803
rect 339294 340954 339914 376398
rect 340094 362813 340154 603195
rect 340643 597820 340709 597821
rect 340643 597756 340644 597820
rect 340708 597756 340709 597820
rect 340643 597755 340709 597756
rect 340646 592653 340706 597755
rect 343794 597438 344414 632898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 597438 348914 601398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 597438 353414 605898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 597438 357914 610398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 597438 362414 614898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 597438 366914 619398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 597438 371414 623898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 597438 375914 628398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597438 380414 632898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 597438 384914 601398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 597438 389414 605898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 597438 393914 610398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 597438 398414 614898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 597438 402914 619398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 597438 407414 623898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 597438 411914 628398
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597438 416414 632898
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 597438 420914 601398
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 597438 425414 605898
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 597438 429914 610398
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 597438 434414 614898
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 597438 438914 619398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 597438 443414 623898
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 597438 447914 628398
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597438 452414 632898
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 597438 456914 601398
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 597438 461414 605898
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 597438 465914 610398
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 597438 470414 614898
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 597438 474914 619398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 597438 479414 623898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 597438 483914 628398
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597438 488414 632898
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 597438 492914 601398
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 597438 497414 605898
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 597438 501914 610398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 597438 506414 614898
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 597438 510914 619398
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 597438 515414 623898
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 597438 519914 628398
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597438 524414 632898
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 597438 528914 601398
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 597438 533414 605898
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 534027 597684 534093 597685
rect 534027 597620 534028 597684
rect 534092 597620 534093 597684
rect 534027 597619 534093 597620
rect 340643 592652 340709 592653
rect 340643 592588 340644 592652
rect 340708 592588 340709 592652
rect 340643 592587 340709 592588
rect 533659 586396 533725 586397
rect 533659 586332 533660 586396
rect 533724 586332 533725 586396
rect 533659 586331 533725 586332
rect 359568 583954 359888 583986
rect 359568 583718 359610 583954
rect 359846 583718 359888 583954
rect 359568 583634 359888 583718
rect 359568 583398 359610 583634
rect 359846 583398 359888 583634
rect 359568 583366 359888 583398
rect 390288 583954 390608 583986
rect 390288 583718 390330 583954
rect 390566 583718 390608 583954
rect 390288 583634 390608 583718
rect 390288 583398 390330 583634
rect 390566 583398 390608 583634
rect 390288 583366 390608 583398
rect 421008 583954 421328 583986
rect 421008 583718 421050 583954
rect 421286 583718 421328 583954
rect 421008 583634 421328 583718
rect 421008 583398 421050 583634
rect 421286 583398 421328 583634
rect 421008 583366 421328 583398
rect 451728 583954 452048 583986
rect 451728 583718 451770 583954
rect 452006 583718 452048 583954
rect 451728 583634 452048 583718
rect 451728 583398 451770 583634
rect 452006 583398 452048 583634
rect 451728 583366 452048 583398
rect 482448 583954 482768 583986
rect 482448 583718 482490 583954
rect 482726 583718 482768 583954
rect 482448 583634 482768 583718
rect 482448 583398 482490 583634
rect 482726 583398 482768 583634
rect 482448 583366 482768 583398
rect 513168 583954 513488 583986
rect 513168 583718 513210 583954
rect 513446 583718 513488 583954
rect 513168 583634 513488 583718
rect 513168 583398 513210 583634
rect 513446 583398 513488 583634
rect 513168 583366 513488 583398
rect 344208 579454 344528 579486
rect 344208 579218 344250 579454
rect 344486 579218 344528 579454
rect 344208 579134 344528 579218
rect 344208 578898 344250 579134
rect 344486 578898 344528 579134
rect 344208 578866 344528 578898
rect 374928 579454 375248 579486
rect 374928 579218 374970 579454
rect 375206 579218 375248 579454
rect 374928 579134 375248 579218
rect 374928 578898 374970 579134
rect 375206 578898 375248 579134
rect 374928 578866 375248 578898
rect 405648 579454 405968 579486
rect 405648 579218 405690 579454
rect 405926 579218 405968 579454
rect 405648 579134 405968 579218
rect 405648 578898 405690 579134
rect 405926 578898 405968 579134
rect 405648 578866 405968 578898
rect 436368 579454 436688 579486
rect 436368 579218 436410 579454
rect 436646 579218 436688 579454
rect 436368 579134 436688 579218
rect 436368 578898 436410 579134
rect 436646 578898 436688 579134
rect 436368 578866 436688 578898
rect 467088 579454 467408 579486
rect 467088 579218 467130 579454
rect 467366 579218 467408 579454
rect 467088 579134 467408 579218
rect 467088 578898 467130 579134
rect 467366 578898 467408 579134
rect 467088 578866 467408 578898
rect 497808 579454 498128 579486
rect 497808 579218 497850 579454
rect 498086 579218 498128 579454
rect 497808 579134 498128 579218
rect 497808 578898 497850 579134
rect 498086 578898 498128 579134
rect 497808 578866 498128 578898
rect 528528 579454 528848 579486
rect 528528 579218 528570 579454
rect 528806 579218 528848 579454
rect 528528 579134 528848 579218
rect 528528 578898 528570 579134
rect 528806 578898 528848 579134
rect 528528 578866 528848 578898
rect 359568 547954 359888 547986
rect 359568 547718 359610 547954
rect 359846 547718 359888 547954
rect 359568 547634 359888 547718
rect 359568 547398 359610 547634
rect 359846 547398 359888 547634
rect 359568 547366 359888 547398
rect 390288 547954 390608 547986
rect 390288 547718 390330 547954
rect 390566 547718 390608 547954
rect 390288 547634 390608 547718
rect 390288 547398 390330 547634
rect 390566 547398 390608 547634
rect 390288 547366 390608 547398
rect 421008 547954 421328 547986
rect 421008 547718 421050 547954
rect 421286 547718 421328 547954
rect 421008 547634 421328 547718
rect 421008 547398 421050 547634
rect 421286 547398 421328 547634
rect 421008 547366 421328 547398
rect 451728 547954 452048 547986
rect 451728 547718 451770 547954
rect 452006 547718 452048 547954
rect 451728 547634 452048 547718
rect 451728 547398 451770 547634
rect 452006 547398 452048 547634
rect 451728 547366 452048 547398
rect 482448 547954 482768 547986
rect 482448 547718 482490 547954
rect 482726 547718 482768 547954
rect 482448 547634 482768 547718
rect 482448 547398 482490 547634
rect 482726 547398 482768 547634
rect 482448 547366 482768 547398
rect 513168 547954 513488 547986
rect 513168 547718 513210 547954
rect 513446 547718 513488 547954
rect 513168 547634 513488 547718
rect 513168 547398 513210 547634
rect 513446 547398 513488 547634
rect 513168 547366 513488 547398
rect 344208 543454 344528 543486
rect 344208 543218 344250 543454
rect 344486 543218 344528 543454
rect 344208 543134 344528 543218
rect 344208 542898 344250 543134
rect 344486 542898 344528 543134
rect 344208 542866 344528 542898
rect 374928 543454 375248 543486
rect 374928 543218 374970 543454
rect 375206 543218 375248 543454
rect 374928 543134 375248 543218
rect 374928 542898 374970 543134
rect 375206 542898 375248 543134
rect 374928 542866 375248 542898
rect 405648 543454 405968 543486
rect 405648 543218 405690 543454
rect 405926 543218 405968 543454
rect 405648 543134 405968 543218
rect 405648 542898 405690 543134
rect 405926 542898 405968 543134
rect 405648 542866 405968 542898
rect 436368 543454 436688 543486
rect 436368 543218 436410 543454
rect 436646 543218 436688 543454
rect 436368 543134 436688 543218
rect 436368 542898 436410 543134
rect 436646 542898 436688 543134
rect 436368 542866 436688 542898
rect 467088 543454 467408 543486
rect 467088 543218 467130 543454
rect 467366 543218 467408 543454
rect 467088 543134 467408 543218
rect 467088 542898 467130 543134
rect 467366 542898 467408 543134
rect 467088 542866 467408 542898
rect 497808 543454 498128 543486
rect 497808 543218 497850 543454
rect 498086 543218 498128 543454
rect 497808 543134 498128 543218
rect 497808 542898 497850 543134
rect 498086 542898 498128 543134
rect 497808 542866 498128 542898
rect 528528 543454 528848 543486
rect 528528 543218 528570 543454
rect 528806 543218 528848 543454
rect 528528 543134 528848 543218
rect 528528 542898 528570 543134
rect 528806 542898 528848 543134
rect 528528 542866 528848 542898
rect 359568 511954 359888 511986
rect 359568 511718 359610 511954
rect 359846 511718 359888 511954
rect 359568 511634 359888 511718
rect 359568 511398 359610 511634
rect 359846 511398 359888 511634
rect 359568 511366 359888 511398
rect 390288 511954 390608 511986
rect 390288 511718 390330 511954
rect 390566 511718 390608 511954
rect 390288 511634 390608 511718
rect 390288 511398 390330 511634
rect 390566 511398 390608 511634
rect 390288 511366 390608 511398
rect 421008 511954 421328 511986
rect 421008 511718 421050 511954
rect 421286 511718 421328 511954
rect 421008 511634 421328 511718
rect 421008 511398 421050 511634
rect 421286 511398 421328 511634
rect 421008 511366 421328 511398
rect 451728 511954 452048 511986
rect 451728 511718 451770 511954
rect 452006 511718 452048 511954
rect 451728 511634 452048 511718
rect 451728 511398 451770 511634
rect 452006 511398 452048 511634
rect 451728 511366 452048 511398
rect 482448 511954 482768 511986
rect 482448 511718 482490 511954
rect 482726 511718 482768 511954
rect 482448 511634 482768 511718
rect 482448 511398 482490 511634
rect 482726 511398 482768 511634
rect 482448 511366 482768 511398
rect 513168 511954 513488 511986
rect 513168 511718 513210 511954
rect 513446 511718 513488 511954
rect 513168 511634 513488 511718
rect 513168 511398 513210 511634
rect 513446 511398 513488 511634
rect 513168 511366 513488 511398
rect 344208 507454 344528 507486
rect 344208 507218 344250 507454
rect 344486 507218 344528 507454
rect 344208 507134 344528 507218
rect 344208 506898 344250 507134
rect 344486 506898 344528 507134
rect 344208 506866 344528 506898
rect 374928 507454 375248 507486
rect 374928 507218 374970 507454
rect 375206 507218 375248 507454
rect 374928 507134 375248 507218
rect 374928 506898 374970 507134
rect 375206 506898 375248 507134
rect 374928 506866 375248 506898
rect 405648 507454 405968 507486
rect 405648 507218 405690 507454
rect 405926 507218 405968 507454
rect 405648 507134 405968 507218
rect 405648 506898 405690 507134
rect 405926 506898 405968 507134
rect 405648 506866 405968 506898
rect 436368 507454 436688 507486
rect 436368 507218 436410 507454
rect 436646 507218 436688 507454
rect 436368 507134 436688 507218
rect 436368 506898 436410 507134
rect 436646 506898 436688 507134
rect 436368 506866 436688 506898
rect 467088 507454 467408 507486
rect 467088 507218 467130 507454
rect 467366 507218 467408 507454
rect 467088 507134 467408 507218
rect 467088 506898 467130 507134
rect 467366 506898 467408 507134
rect 467088 506866 467408 506898
rect 497808 507454 498128 507486
rect 497808 507218 497850 507454
rect 498086 507218 498128 507454
rect 497808 507134 498128 507218
rect 497808 506898 497850 507134
rect 498086 506898 498128 507134
rect 497808 506866 498128 506898
rect 528528 507454 528848 507486
rect 528528 507218 528570 507454
rect 528806 507218 528848 507454
rect 528528 507134 528848 507218
rect 528528 506898 528570 507134
rect 528806 506898 528848 507134
rect 528528 506866 528848 506898
rect 359568 475954 359888 475986
rect 359568 475718 359610 475954
rect 359846 475718 359888 475954
rect 359568 475634 359888 475718
rect 359568 475398 359610 475634
rect 359846 475398 359888 475634
rect 359568 475366 359888 475398
rect 390288 475954 390608 475986
rect 390288 475718 390330 475954
rect 390566 475718 390608 475954
rect 390288 475634 390608 475718
rect 390288 475398 390330 475634
rect 390566 475398 390608 475634
rect 390288 475366 390608 475398
rect 421008 475954 421328 475986
rect 421008 475718 421050 475954
rect 421286 475718 421328 475954
rect 421008 475634 421328 475718
rect 421008 475398 421050 475634
rect 421286 475398 421328 475634
rect 421008 475366 421328 475398
rect 451728 475954 452048 475986
rect 451728 475718 451770 475954
rect 452006 475718 452048 475954
rect 451728 475634 452048 475718
rect 451728 475398 451770 475634
rect 452006 475398 452048 475634
rect 451728 475366 452048 475398
rect 482448 475954 482768 475986
rect 482448 475718 482490 475954
rect 482726 475718 482768 475954
rect 482448 475634 482768 475718
rect 482448 475398 482490 475634
rect 482726 475398 482768 475634
rect 482448 475366 482768 475398
rect 513168 475954 513488 475986
rect 513168 475718 513210 475954
rect 513446 475718 513488 475954
rect 513168 475634 513488 475718
rect 513168 475398 513210 475634
rect 513446 475398 513488 475634
rect 513168 475366 513488 475398
rect 344208 471454 344528 471486
rect 344208 471218 344250 471454
rect 344486 471218 344528 471454
rect 344208 471134 344528 471218
rect 344208 470898 344250 471134
rect 344486 470898 344528 471134
rect 344208 470866 344528 470898
rect 374928 471454 375248 471486
rect 374928 471218 374970 471454
rect 375206 471218 375248 471454
rect 374928 471134 375248 471218
rect 374928 470898 374970 471134
rect 375206 470898 375248 471134
rect 374928 470866 375248 470898
rect 405648 471454 405968 471486
rect 405648 471218 405690 471454
rect 405926 471218 405968 471454
rect 405648 471134 405968 471218
rect 405648 470898 405690 471134
rect 405926 470898 405968 471134
rect 405648 470866 405968 470898
rect 436368 471454 436688 471486
rect 436368 471218 436410 471454
rect 436646 471218 436688 471454
rect 436368 471134 436688 471218
rect 436368 470898 436410 471134
rect 436646 470898 436688 471134
rect 436368 470866 436688 470898
rect 467088 471454 467408 471486
rect 467088 471218 467130 471454
rect 467366 471218 467408 471454
rect 467088 471134 467408 471218
rect 467088 470898 467130 471134
rect 467366 470898 467408 471134
rect 467088 470866 467408 470898
rect 497808 471454 498128 471486
rect 497808 471218 497850 471454
rect 498086 471218 498128 471454
rect 497808 471134 498128 471218
rect 497808 470898 497850 471134
rect 498086 470898 498128 471134
rect 497808 470866 498128 470898
rect 528528 471454 528848 471486
rect 528528 471218 528570 471454
rect 528806 471218 528848 471454
rect 528528 471134 528848 471218
rect 528528 470898 528570 471134
rect 528806 470898 528848 471134
rect 528528 470866 528848 470898
rect 359568 439954 359888 439986
rect 359568 439718 359610 439954
rect 359846 439718 359888 439954
rect 359568 439634 359888 439718
rect 359568 439398 359610 439634
rect 359846 439398 359888 439634
rect 359568 439366 359888 439398
rect 390288 439954 390608 439986
rect 390288 439718 390330 439954
rect 390566 439718 390608 439954
rect 390288 439634 390608 439718
rect 390288 439398 390330 439634
rect 390566 439398 390608 439634
rect 390288 439366 390608 439398
rect 421008 439954 421328 439986
rect 421008 439718 421050 439954
rect 421286 439718 421328 439954
rect 421008 439634 421328 439718
rect 421008 439398 421050 439634
rect 421286 439398 421328 439634
rect 421008 439366 421328 439398
rect 451728 439954 452048 439986
rect 451728 439718 451770 439954
rect 452006 439718 452048 439954
rect 451728 439634 452048 439718
rect 451728 439398 451770 439634
rect 452006 439398 452048 439634
rect 451728 439366 452048 439398
rect 482448 439954 482768 439986
rect 482448 439718 482490 439954
rect 482726 439718 482768 439954
rect 482448 439634 482768 439718
rect 482448 439398 482490 439634
rect 482726 439398 482768 439634
rect 482448 439366 482768 439398
rect 513168 439954 513488 439986
rect 513168 439718 513210 439954
rect 513446 439718 513488 439954
rect 513168 439634 513488 439718
rect 513168 439398 513210 439634
rect 513446 439398 513488 439634
rect 513168 439366 513488 439398
rect 344208 435454 344528 435486
rect 344208 435218 344250 435454
rect 344486 435218 344528 435454
rect 344208 435134 344528 435218
rect 344208 434898 344250 435134
rect 344486 434898 344528 435134
rect 344208 434866 344528 434898
rect 374928 435454 375248 435486
rect 374928 435218 374970 435454
rect 375206 435218 375248 435454
rect 374928 435134 375248 435218
rect 374928 434898 374970 435134
rect 375206 434898 375248 435134
rect 374928 434866 375248 434898
rect 405648 435454 405968 435486
rect 405648 435218 405690 435454
rect 405926 435218 405968 435454
rect 405648 435134 405968 435218
rect 405648 434898 405690 435134
rect 405926 434898 405968 435134
rect 405648 434866 405968 434898
rect 436368 435454 436688 435486
rect 436368 435218 436410 435454
rect 436646 435218 436688 435454
rect 436368 435134 436688 435218
rect 436368 434898 436410 435134
rect 436646 434898 436688 435134
rect 436368 434866 436688 434898
rect 467088 435454 467408 435486
rect 467088 435218 467130 435454
rect 467366 435218 467408 435454
rect 467088 435134 467408 435218
rect 467088 434898 467130 435134
rect 467366 434898 467408 435134
rect 467088 434866 467408 434898
rect 497808 435454 498128 435486
rect 497808 435218 497850 435454
rect 498086 435218 498128 435454
rect 497808 435134 498128 435218
rect 497808 434898 497850 435134
rect 498086 434898 498128 435134
rect 497808 434866 498128 434898
rect 528528 435454 528848 435486
rect 528528 435218 528570 435454
rect 528806 435218 528848 435454
rect 528528 435134 528848 435218
rect 528528 434898 528570 435134
rect 528806 434898 528848 435134
rect 528528 434866 528848 434898
rect 359568 403954 359888 403986
rect 359568 403718 359610 403954
rect 359846 403718 359888 403954
rect 359568 403634 359888 403718
rect 359568 403398 359610 403634
rect 359846 403398 359888 403634
rect 359568 403366 359888 403398
rect 390288 403954 390608 403986
rect 390288 403718 390330 403954
rect 390566 403718 390608 403954
rect 390288 403634 390608 403718
rect 390288 403398 390330 403634
rect 390566 403398 390608 403634
rect 390288 403366 390608 403398
rect 421008 403954 421328 403986
rect 421008 403718 421050 403954
rect 421286 403718 421328 403954
rect 421008 403634 421328 403718
rect 421008 403398 421050 403634
rect 421286 403398 421328 403634
rect 421008 403366 421328 403398
rect 451728 403954 452048 403986
rect 451728 403718 451770 403954
rect 452006 403718 452048 403954
rect 451728 403634 452048 403718
rect 451728 403398 451770 403634
rect 452006 403398 452048 403634
rect 451728 403366 452048 403398
rect 482448 403954 482768 403986
rect 482448 403718 482490 403954
rect 482726 403718 482768 403954
rect 482448 403634 482768 403718
rect 482448 403398 482490 403634
rect 482726 403398 482768 403634
rect 482448 403366 482768 403398
rect 513168 403954 513488 403986
rect 513168 403718 513210 403954
rect 513446 403718 513488 403954
rect 513168 403634 513488 403718
rect 513168 403398 513210 403634
rect 513446 403398 513488 403634
rect 513168 403366 513488 403398
rect 340275 400892 340341 400893
rect 340275 400828 340276 400892
rect 340340 400828 340341 400892
rect 340275 400827 340341 400828
rect 340278 398445 340338 400827
rect 340275 398444 340341 398445
rect 340275 398380 340276 398444
rect 340340 398380 340341 398444
rect 340275 398379 340341 398380
rect 343794 381454 344414 398000
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 342851 368524 342917 368525
rect 342851 368460 342852 368524
rect 342916 368460 342917 368524
rect 342851 368459 342917 368460
rect 340091 362812 340157 362813
rect 340091 362748 340092 362812
rect 340156 362748 340157 362812
rect 340091 362747 340157 362748
rect 340091 360908 340157 360909
rect 340091 360844 340092 360908
rect 340156 360844 340157 360908
rect 340091 360843 340157 360844
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 337883 178804 337949 178805
rect 337883 178740 337884 178804
rect 337948 178740 337949 178804
rect 337883 178739 337949 178740
rect 337886 160037 337946 178739
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 337883 160036 337949 160037
rect 337883 159972 337884 160036
rect 337948 159972 337949 160036
rect 337883 159971 337949 159972
rect 337886 158813 337946 159971
rect 337883 158812 337949 158813
rect 337883 158748 337884 158812
rect 337948 158748 337949 158812
rect 337883 158747 337949 158748
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 336779 26212 336845 26213
rect 336779 26148 336780 26212
rect 336844 26148 336845 26212
rect 336779 26147 336845 26148
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 16954 339914 52398
rect 340094 42805 340154 360843
rect 341379 265028 341445 265029
rect 341379 264964 341380 265028
rect 341444 264964 341445 265028
rect 341379 264963 341445 264964
rect 341382 136645 341442 264963
rect 342299 224500 342365 224501
rect 342299 224436 342300 224500
rect 342364 224436 342365 224500
rect 342299 224435 342365 224436
rect 341379 136644 341445 136645
rect 341379 136580 341380 136644
rect 341444 136580 341445 136644
rect 341379 136579 341445 136580
rect 342302 131205 342362 224435
rect 342854 174589 342914 368459
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 342851 174588 342917 174589
rect 342851 174524 342852 174588
rect 342916 174524 342917 174588
rect 342851 174523 342917 174524
rect 343794 165454 344414 200898
rect 348294 385954 348914 398000
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 346347 191180 346413 191181
rect 346347 191116 346348 191180
rect 346412 191116 346413 191180
rect 346347 191115 346413 191116
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 342299 131204 342365 131205
rect 342299 131140 342300 131204
rect 342364 131140 342365 131204
rect 342299 131139 342365 131140
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 346350 117333 346410 191115
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 346347 117332 346413 117333
rect 346347 117268 346348 117332
rect 346412 117268 346413 117332
rect 346347 117267 346413 117268
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 340091 42804 340157 42805
rect 340091 42740 340092 42804
rect 340156 42740 340157 42804
rect 340091 42739 340157 42740
rect 340094 42125 340154 42739
rect 340091 42124 340157 42125
rect 340091 42060 340092 42124
rect 340156 42060 340157 42124
rect 340091 42059 340157 42060
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 390454 353414 398000
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 394954 357914 398000
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 363454 362414 398000
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 367954 366914 398000
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 372454 371414 398000
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 375294 376954 375914 398000
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 373211 286380 373277 286381
rect 373211 286316 373212 286380
rect 373276 286316 373277 286380
rect 373211 286315 373277 286316
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 373214 102781 373274 286315
rect 375294 268954 375914 304398
rect 379794 381454 380414 398000
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 302000 380414 308898
rect 384294 385954 384914 398000
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 302000 384914 313398
rect 388794 390454 389414 398000
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 302000 389414 317898
rect 393294 394954 393914 398000
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 302000 393914 322398
rect 397794 363454 398414 398000
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 302000 398414 326898
rect 402294 367954 402914 398000
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 302000 402914 331398
rect 406794 372454 407414 398000
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 302000 407414 335898
rect 411294 376954 411914 398000
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 302000 411914 304398
rect 415794 381454 416414 398000
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 302000 416414 308898
rect 420294 385954 420914 398000
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 302000 420914 313398
rect 424794 390454 425414 398000
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 302000 425414 317898
rect 429294 394954 429914 398000
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 302000 429914 322398
rect 433794 363454 434414 398000
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 302000 434414 326898
rect 438294 367954 438914 398000
rect 439083 387700 439149 387701
rect 439083 387636 439084 387700
rect 439148 387636 439149 387700
rect 439083 387635 439149 387636
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 302000 438914 331398
rect 439086 306390 439146 387635
rect 442794 372454 443414 398000
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 439086 306330 439514 306390
rect 399568 295954 399888 295986
rect 399568 295718 399610 295954
rect 399846 295718 399888 295954
rect 399568 295634 399888 295718
rect 399568 295398 399610 295634
rect 399846 295398 399888 295634
rect 399568 295366 399888 295398
rect 430288 295954 430608 295986
rect 430288 295718 430330 295954
rect 430566 295718 430608 295954
rect 430288 295634 430608 295718
rect 430288 295398 430330 295634
rect 430566 295398 430608 295634
rect 430288 295366 430608 295398
rect 376155 291820 376221 291821
rect 376155 291756 376156 291820
rect 376220 291756 376221 291820
rect 376155 291755 376221 291756
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 376158 238781 376218 291755
rect 384208 291454 384528 291486
rect 384208 291218 384250 291454
rect 384486 291218 384528 291454
rect 384208 291134 384528 291218
rect 384208 290898 384250 291134
rect 384486 290898 384528 291134
rect 384208 290866 384528 290898
rect 414928 291454 415248 291486
rect 414928 291218 414970 291454
rect 415206 291218 415248 291454
rect 414928 291134 415248 291218
rect 414928 290898 414970 291134
rect 415206 290898 415248 291134
rect 414928 290866 415248 290898
rect 439454 289645 439514 306330
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 439451 289644 439517 289645
rect 439451 289580 439452 289644
rect 439516 289580 439517 289644
rect 439451 289579 439517 289580
rect 378731 269244 378797 269245
rect 378731 269180 378732 269244
rect 378796 269180 378797 269244
rect 378731 269179 378797 269180
rect 377995 263260 378061 263261
rect 377995 263196 377996 263260
rect 378060 263196 378061 263260
rect 377995 263195 378061 263196
rect 376155 238780 376221 238781
rect 376155 238716 376156 238780
rect 376220 238716 376221 238780
rect 376155 238715 376221 238716
rect 377998 236061 378058 263195
rect 377995 236060 378061 236061
rect 377995 235996 377996 236060
rect 378060 235996 378061 236060
rect 377995 235995 378061 235996
rect 378734 233205 378794 269179
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 399568 259954 399888 259986
rect 399568 259718 399610 259954
rect 399846 259718 399888 259954
rect 399568 259634 399888 259718
rect 399568 259398 399610 259634
rect 399846 259398 399888 259634
rect 399568 259366 399888 259398
rect 430288 259954 430608 259986
rect 430288 259718 430330 259954
rect 430566 259718 430608 259954
rect 430288 259634 430608 259718
rect 430288 259398 430330 259634
rect 430566 259398 430608 259634
rect 430288 259366 430608 259398
rect 378915 257004 378981 257005
rect 378915 256940 378916 257004
rect 378980 256940 378981 257004
rect 378915 256939 378981 256940
rect 378731 233204 378797 233205
rect 378731 233140 378732 233204
rect 378796 233140 378797 233204
rect 378731 233139 378797 233140
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 378734 226949 378794 233139
rect 378918 227765 378978 256939
rect 384208 255454 384528 255486
rect 384208 255218 384250 255454
rect 384486 255218 384528 255454
rect 384208 255134 384528 255218
rect 384208 254898 384250 255134
rect 384486 254898 384528 255134
rect 384208 254866 384528 254898
rect 414928 255454 415248 255486
rect 414928 255218 414970 255454
rect 415206 255218 415248 255454
rect 414928 255134 415248 255218
rect 414928 254898 414970 255134
rect 415206 254898 415248 255134
rect 414928 254866 415248 254898
rect 382779 241772 382845 241773
rect 382779 241708 382780 241772
rect 382844 241708 382845 241772
rect 382779 241707 382845 241708
rect 379794 237454 380414 238000
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 378915 227764 378981 227765
rect 378915 227700 378916 227764
rect 378980 227700 378981 227764
rect 378915 227699 378981 227700
rect 378731 226948 378797 226949
rect 378731 226884 378732 226948
rect 378796 226884 378797 226948
rect 378731 226883 378797 226884
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 373211 102780 373277 102781
rect 373211 102716 373212 102780
rect 373276 102716 373277 102780
rect 373211 102715 373277 102716
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 201454 380414 236898
rect 380571 236196 380637 236197
rect 380571 236132 380572 236196
rect 380636 236132 380637 236196
rect 380571 236131 380637 236132
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 380574 91085 380634 236131
rect 380939 233340 381005 233341
rect 380939 233276 380940 233340
rect 381004 233276 381005 233340
rect 380939 233275 381005 233276
rect 380942 231845 381002 233275
rect 380939 231844 381005 231845
rect 380939 231780 380940 231844
rect 381004 231780 381005 231844
rect 380939 231779 381005 231780
rect 382782 106453 382842 241707
rect 384294 205954 384914 238000
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 382779 106452 382845 106453
rect 382779 106388 382780 106452
rect 382844 106388 382845 106452
rect 382779 106387 382845 106388
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 380571 91084 380637 91085
rect 380571 91020 380572 91084
rect 380636 91020 380637 91084
rect 380571 91019 380637 91020
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 210454 389414 238000
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 214954 393914 238000
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 397794 219454 398414 238000
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 148000 398414 182898
rect 402294 223954 402914 238000
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 148000 402914 151398
rect 406794 228454 407414 238000
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 148000 407414 155898
rect 411294 232954 411914 238000
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 148000 411914 160398
rect 415794 237454 416414 238000
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 148000 416414 164898
rect 420294 205954 420914 238000
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 148000 420914 169398
rect 424794 210454 425414 238000
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 148000 425414 173898
rect 429294 214954 429914 238000
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 148000 429914 178398
rect 433794 219454 434414 238000
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 148000 434414 182898
rect 438294 223954 438914 238000
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 148000 438914 151398
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 148000 443414 155898
rect 447294 376954 447914 398000
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 451794 381454 452414 398000
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 448467 220964 448533 220965
rect 448467 220900 448468 220964
rect 448532 220900 448533 220964
rect 448467 220899 448533 220900
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 148000 447914 160398
rect 448470 151830 448530 220899
rect 451043 214028 451109 214029
rect 451043 213964 451044 214028
rect 451108 213964 451109 214028
rect 451043 213963 451109 213964
rect 448470 151770 449450 151830
rect 396579 147796 396645 147797
rect 396579 147732 396580 147796
rect 396644 147732 396645 147796
rect 396579 147731 396645 147732
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 396582 112437 396642 147731
rect 449390 143445 449450 151770
rect 450123 146980 450189 146981
rect 450123 146916 450124 146980
rect 450188 146916 450189 146980
rect 450123 146915 450189 146916
rect 449387 143444 449453 143445
rect 449387 143380 449388 143444
rect 449452 143380 449453 143444
rect 449387 143379 449453 143380
rect 419568 115954 419888 115986
rect 419568 115718 419610 115954
rect 419846 115718 419888 115954
rect 419568 115634 419888 115718
rect 419568 115398 419610 115634
rect 419846 115398 419888 115634
rect 419568 115366 419888 115398
rect 396579 112436 396645 112437
rect 396579 112372 396580 112436
rect 396644 112372 396645 112436
rect 396579 112371 396645 112372
rect 449939 112436 450005 112437
rect 449939 112372 449940 112436
rect 450004 112372 450005 112436
rect 449939 112371 450005 112372
rect 404208 111454 404528 111486
rect 404208 111218 404250 111454
rect 404486 111218 404528 111454
rect 404208 111134 404528 111218
rect 404208 110898 404250 111134
rect 404486 110898 404528 111134
rect 404208 110866 404528 110898
rect 434928 111454 435248 111486
rect 434928 111218 434970 111454
rect 435206 111218 435248 111454
rect 434928 111134 435248 111218
rect 434928 110898 434970 111134
rect 435206 110898 435248 111134
rect 434928 110866 435248 110898
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 449387 101012 449453 101013
rect 449387 101010 449388 101012
rect 448470 100950 449388 101010
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 75454 398414 94000
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 79954 402914 94000
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 84454 407414 94000
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 88954 411914 94000
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 93454 416414 94000
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 61954 420914 94000
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 66454 425414 94000
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 70954 429914 94000
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 75454 434414 94000
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 79954 438914 94000
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 84454 443414 94000
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 88954 447914 94000
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 448470 45525 448530 100950
rect 449387 100948 449388 100950
rect 449452 100948 449453 101012
rect 449387 100947 449453 100948
rect 449387 99788 449453 99789
rect 449387 99724 449388 99788
rect 449452 99724 449453 99788
rect 449387 99723 449453 99724
rect 449390 84829 449450 99723
rect 449387 84828 449453 84829
rect 449387 84764 449388 84828
rect 449452 84764 449453 84828
rect 449387 84763 449453 84764
rect 448467 45524 448533 45525
rect 448467 45460 448468 45524
rect 448532 45460 448533 45524
rect 448467 45459 448533 45460
rect 449942 22677 450002 112371
rect 450126 96117 450186 146915
rect 451046 133517 451106 213963
rect 451794 201454 452414 236898
rect 456294 385954 456914 398000
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 454171 224908 454237 224909
rect 454171 224844 454172 224908
rect 454236 224844 454237 224908
rect 454171 224843 454237 224844
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 148000 452414 164898
rect 451411 147796 451477 147797
rect 451411 147732 451412 147796
rect 451476 147732 451477 147796
rect 451411 147731 451477 147732
rect 451043 133516 451109 133517
rect 451043 133452 451044 133516
rect 451108 133452 451109 133516
rect 451043 133451 451109 133452
rect 451414 132157 451474 147731
rect 451411 132156 451477 132157
rect 451411 132092 451412 132156
rect 451476 132092 451477 132156
rect 451411 132091 451477 132092
rect 451043 121548 451109 121549
rect 451043 121484 451044 121548
rect 451108 121484 451109 121548
rect 451043 121483 451109 121484
rect 450123 96116 450189 96117
rect 450123 96052 450124 96116
rect 450188 96052 450189 96116
rect 450123 96051 450189 96052
rect 451046 42805 451106 121483
rect 454174 118149 454234 224843
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 460794 390454 461414 398000
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 458771 149156 458837 149157
rect 458771 149092 458772 149156
rect 458836 149092 458837 149156
rect 458771 149091 458837 149092
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 454171 118148 454237 118149
rect 454171 118084 454172 118148
rect 454236 118084 454237 118148
rect 454171 118083 454237 118084
rect 456294 97954 456914 133398
rect 458774 118829 458834 149091
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 458771 118828 458837 118829
rect 458771 118764 458772 118828
rect 458836 118764 458837 118828
rect 458771 118763 458837 118764
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 451794 93454 452414 94000
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451043 42804 451109 42805
rect 451043 42740 451044 42804
rect 451108 42740 451109 42804
rect 451043 42739 451109 42740
rect 449939 22676 450005 22677
rect 449939 22612 449940 22676
rect 450004 22612 450005 22676
rect 449939 22611 450005 22612
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 394954 465914 398000
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 363454 470414 398000
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 367954 474914 398000
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 372454 479414 398000
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 376954 483914 398000
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 381454 488414 398000
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 385954 492914 398000
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 390454 497414 398000
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 394954 501914 398000
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 363454 506414 398000
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 367954 510914 398000
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 372454 515414 398000
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 376954 519914 398000
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 381454 524414 398000
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 385954 528914 398000
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 390454 533414 398000
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 533662 174589 533722 586331
rect 534030 541517 534090 597619
rect 535499 589116 535565 589117
rect 535499 589052 535500 589116
rect 535564 589052 535565 589116
rect 535499 589051 535565 589052
rect 534395 543556 534461 543557
rect 534395 543492 534396 543556
rect 534460 543492 534461 543556
rect 534395 543491 534461 543492
rect 534027 541516 534093 541517
rect 534027 541452 534028 541516
rect 534092 541452 534093 541516
rect 534027 541451 534093 541452
rect 534211 450396 534277 450397
rect 534211 450332 534212 450396
rect 534276 450332 534277 450396
rect 534211 450331 534277 450332
rect 534214 180029 534274 450331
rect 534211 180028 534277 180029
rect 534211 179964 534212 180028
rect 534276 179964 534277 180028
rect 534211 179963 534277 179964
rect 533659 174588 533725 174589
rect 533659 174524 533660 174588
rect 533724 174524 533725 174588
rect 533659 174523 533725 174524
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 534398 95301 534458 543491
rect 535502 160037 535562 589051
rect 537294 574954 537914 610398
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 539547 599044 539613 599045
rect 539547 598980 539548 599044
rect 539612 598980 539613 599044
rect 539547 598979 539613 598980
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 538443 559196 538509 559197
rect 538443 559132 538444 559196
rect 538508 559132 538509 559196
rect 538443 559131 538509 559132
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 536787 525876 536853 525877
rect 536787 525812 536788 525876
rect 536852 525812 536853 525876
rect 536787 525811 536853 525812
rect 535683 497996 535749 497997
rect 535683 497932 535684 497996
rect 535748 497932 535749 497996
rect 535683 497931 535749 497932
rect 535686 336021 535746 497931
rect 536790 395317 536850 525811
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 538259 480316 538325 480317
rect 538259 480252 538260 480316
rect 538324 480252 538325 480316
rect 538259 480251 538325 480252
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 536787 395316 536853 395317
rect 536787 395252 536788 395316
rect 536852 395252 536853 395316
rect 536787 395251 536853 395252
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 535683 336020 535749 336021
rect 535683 335956 535684 336020
rect 535748 335956 535749 336020
rect 535683 335955 535749 335956
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 535499 160036 535565 160037
rect 535499 159972 535500 160036
rect 535564 159972 535565 160036
rect 535499 159971 535565 159972
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 534395 95300 534461 95301
rect 534395 95236 534396 95300
rect 534460 95236 534461 95300
rect 534395 95235 534461 95236
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 70954 537914 106398
rect 538262 100741 538322 480251
rect 538446 360909 538506 559131
rect 539550 396677 539610 598979
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 542675 455156 542741 455157
rect 542675 455092 542676 455156
rect 542740 455092 542741 455156
rect 542675 455091 542741 455092
rect 542678 451290 542738 455091
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541019 425236 541085 425237
rect 541019 425172 541020 425236
rect 541084 425172 541085 425236
rect 541019 425171 541085 425172
rect 539547 396676 539613 396677
rect 539547 396612 539548 396676
rect 539612 396612 539613 396676
rect 539547 396611 539613 396612
rect 541022 395453 541082 425171
rect 541794 399454 542414 434898
rect 542494 451230 542738 451290
rect 542494 402990 542554 451230
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 543779 437476 543845 437477
rect 543779 437412 543780 437476
rect 543844 437412 543845 437476
rect 543779 437411 543845 437412
rect 542494 402930 542738 402990
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541019 395452 541085 395453
rect 541019 395388 541020 395452
rect 541084 395388 541085 395452
rect 541019 395387 541085 395388
rect 541794 363454 542414 398898
rect 542678 382941 542738 402930
rect 543782 393277 543842 437411
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 543779 393276 543845 393277
rect 543779 393212 543780 393276
rect 543844 393212 543845 393276
rect 543779 393211 543845 393212
rect 542675 382940 542741 382941
rect 542675 382876 542676 382940
rect 542740 382876 542741 382940
rect 542675 382875 542741 382876
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 538443 360908 538509 360909
rect 538443 360844 538444 360908
rect 538508 360844 538509 360908
rect 538443 360843 538509 360844
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 538259 100740 538325 100741
rect 538259 100676 538260 100740
rect 538324 100676 538325 100740
rect 538259 100675 538325 100676
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< obsm4 >>
rect 68800 174494 96960 174600
rect 97020 174494 98320 174600
rect 98380 174494 99408 174600
rect 99468 174494 100768 174600
rect 100828 174494 101992 174600
rect 102052 174494 103352 174600
rect 103412 174494 104576 174600
rect 104636 174494 105664 174600
rect 105724 174494 107024 174600
rect 107084 174494 108112 174600
rect 108172 174494 109472 174600
rect 109532 174494 110696 174600
rect 110756 174494 112056 174600
rect 112116 174494 113144 174600
rect 113204 174494 114368 174600
rect 114428 174494 115728 174600
rect 115788 174494 116952 174600
rect 117012 174494 118312 174600
rect 118372 174494 119400 174600
rect 119460 174494 120760 174600
rect 120820 174494 121848 174600
rect 121908 174494 123072 174600
rect 123132 174494 124432 174600
rect 124492 174494 125656 174600
rect 125716 174494 127016 174600
rect 127076 174494 128104 174600
rect 128164 174494 129464 174600
rect 129524 174494 130688 174600
rect 130748 174494 132048 174600
rect 132108 174494 133136 174600
rect 133196 174494 134360 174600
rect 134420 174494 135720 174600
rect 135780 174494 148232 174600
rect 148292 174494 158840 174600
rect 158900 174494 164756 174600
rect 68800 151986 164756 174494
rect 68800 151366 69072 151986
rect 69420 151366 164136 151986
rect 164484 151366 164756 151986
rect 68800 147486 164756 151366
rect 68800 146866 69752 147486
rect 70100 146866 163456 147486
rect 163804 146866 164756 147486
rect 68800 115986 164756 146866
rect 68800 115366 69072 115986
rect 69420 115366 164136 115986
rect 164484 115366 164756 115986
rect 68800 111486 164756 115366
rect 68800 110866 69752 111486
rect 70100 110866 163456 111486
rect 163804 110866 164756 111486
rect 68800 95200 164756 110866
rect 68800 95100 74656 95200
rect 74716 95100 84312 95200
rect 84372 95100 85536 95200
rect 85596 95100 86624 95200
rect 86684 95100 87984 95200
rect 88044 95100 88936 95200
rect 88996 95100 90160 95200
rect 90220 95100 91384 95200
rect 91444 95100 92472 95200
rect 92532 95100 93832 95200
rect 93892 95100 94920 95200
rect 94980 95100 96008 95200
rect 96068 95100 96688 95200
rect 96748 95100 97096 95200
rect 97156 95100 98048 95200
rect 98108 95100 98456 95200
rect 98516 95100 99136 95200
rect 99196 95100 99544 95200
rect 99604 95100 100632 95200
rect 100692 95100 100768 95200
rect 100828 95100 101856 95200
rect 101916 95100 101992 95200
rect 102052 95100 102944 95200
rect 103004 95100 103216 95200
rect 103276 95100 104304 95200
rect 104364 95100 104440 95200
rect 104500 95100 105392 95200
rect 105452 95100 105664 95200
rect 105724 95100 106480 95200
rect 106540 95100 106616 95200
rect 106676 95100 107704 95200
rect 107764 95100 108112 95200
rect 108172 95100 109064 95200
rect 109124 95100 109472 95200
rect 109532 95100 110152 95200
rect 110212 95100 110696 95200
rect 110756 95100 111240 95200
rect 111300 95100 111920 95200
rect 111980 95100 112328 95200
rect 112388 95100 113144 95200
rect 113204 95100 113688 95200
rect 113748 95100 114368 95200
rect 114428 95100 114776 95200
rect 114836 95100 115456 95200
rect 115516 95100 115864 95200
rect 115924 95100 116680 95200
rect 116740 95100 117088 95200
rect 117148 95100 117904 95200
rect 117964 95100 118176 95200
rect 118236 95100 119400 95200
rect 119460 95100 119536 95200
rect 119596 95100 120216 95200
rect 120276 95100 120624 95200
rect 120684 95100 121712 95200
rect 121772 95100 121984 95200
rect 122044 95100 122800 95200
rect 122860 95100 123208 95200
rect 123268 95100 124024 95200
rect 124084 95100 124432 95200
rect 124492 95100 125384 95200
rect 125444 95100 125656 95200
rect 125716 95100 126472 95200
rect 126532 95100 126608 95200
rect 126668 95100 128104 95200
rect 128164 95100 129328 95200
rect 129388 95100 130688 95200
rect 130748 95100 131912 95200
rect 131972 95100 133136 95200
rect 133196 95100 134360 95200
rect 134420 95100 135584 95200
rect 135644 95100 151496 95200
rect 151556 95100 151632 95200
rect 151692 95100 151768 95200
rect 151828 95100 151904 95200
rect 151964 95100 164756 95200
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 68250 579218 68486 579454
rect 68250 578898 68486 579134
rect 98970 579218 99206 579454
rect 98970 578898 99206 579134
rect 129690 579218 129926 579454
rect 129690 578898 129926 579134
rect 160410 579218 160646 579454
rect 160410 578898 160646 579134
rect 191130 579218 191366 579454
rect 191130 578898 191366 579134
rect 221850 579218 222086 579454
rect 221850 578898 222086 579134
rect 83610 547718 83846 547954
rect 83610 547398 83846 547634
rect 114330 547718 114566 547954
rect 114330 547398 114566 547634
rect 145050 547718 145286 547954
rect 145050 547398 145286 547634
rect 175770 547718 176006 547954
rect 175770 547398 176006 547634
rect 206490 547718 206726 547954
rect 206490 547398 206726 547634
rect 237210 547718 237446 547954
rect 237210 547398 237446 547634
rect 68250 543218 68486 543454
rect 68250 542898 68486 543134
rect 98970 543218 99206 543454
rect 98970 542898 99206 543134
rect 129690 543218 129926 543454
rect 129690 542898 129926 543134
rect 160410 543218 160646 543454
rect 160410 542898 160646 543134
rect 191130 543218 191366 543454
rect 191130 542898 191366 543134
rect 221850 543218 222086 543454
rect 221850 542898 222086 543134
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 83610 511718 83846 511954
rect 83610 511398 83846 511634
rect 114330 511718 114566 511954
rect 114330 511398 114566 511634
rect 145050 511718 145286 511954
rect 145050 511398 145286 511634
rect 175770 511718 176006 511954
rect 175770 511398 176006 511634
rect 206490 511718 206726 511954
rect 206490 511398 206726 511634
rect 237210 511718 237446 511954
rect 237210 511398 237446 511634
rect 68250 507218 68486 507454
rect 68250 506898 68486 507134
rect 98970 507218 99206 507454
rect 98970 506898 99206 507134
rect 129690 507218 129926 507454
rect 129690 506898 129926 507134
rect 160410 507218 160646 507454
rect 160410 506898 160646 507134
rect 191130 507218 191366 507454
rect 191130 506898 191366 507134
rect 221850 507218 222086 507454
rect 221850 506898 222086 507134
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 83610 475718 83846 475954
rect 83610 475398 83846 475634
rect 114330 475718 114566 475954
rect 114330 475398 114566 475634
rect 145050 475718 145286 475954
rect 145050 475398 145286 475634
rect 175770 475718 176006 475954
rect 175770 475398 176006 475634
rect 206490 475718 206726 475954
rect 206490 475398 206726 475634
rect 237210 475718 237446 475954
rect 237210 475398 237446 475634
rect 68250 471218 68486 471454
rect 68250 470898 68486 471134
rect 98970 471218 99206 471454
rect 98970 470898 99206 471134
rect 129690 471218 129926 471454
rect 129690 470898 129926 471134
rect 160410 471218 160646 471454
rect 160410 470898 160646 471134
rect 191130 471218 191366 471454
rect 191130 470898 191366 471134
rect 221850 471218 222086 471454
rect 221850 470898 222086 471134
rect 83610 439718 83846 439954
rect 83610 439398 83846 439634
rect 114330 439718 114566 439954
rect 114330 439398 114566 439634
rect 145050 439718 145286 439954
rect 145050 439398 145286 439634
rect 175770 439718 176006 439954
rect 175770 439398 176006 439634
rect 206490 439718 206726 439954
rect 206490 439398 206726 439634
rect 237210 439718 237446 439954
rect 237210 439398 237446 439634
rect 68250 435218 68486 435454
rect 68250 434898 68486 435134
rect 98970 435218 99206 435454
rect 98970 434898 99206 435134
rect 129690 435218 129926 435454
rect 129690 434898 129926 435134
rect 160410 435218 160646 435454
rect 160410 434898 160646 435134
rect 191130 435218 191366 435454
rect 191130 434898 191366 435134
rect 221850 435218 222086 435454
rect 221850 434898 222086 435134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 89610 259718 89846 259954
rect 89610 259398 89846 259634
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 69128 151718 69364 151954
rect 69128 151398 69364 151634
rect 164192 151718 164428 151954
rect 164192 151398 164428 151634
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 115718 69364 115954
rect 69128 115398 69364 115634
rect 164192 115718 164428 115954
rect 164192 115398 164428 115634
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 199610 331718 199846 331954
rect 199610 331398 199846 331634
rect 230330 331718 230566 331954
rect 230330 331398 230566 331634
rect 261050 331718 261286 331954
rect 261050 331398 261286 331634
rect 184250 327218 184486 327454
rect 184250 326898 184486 327134
rect 214970 327218 215206 327454
rect 214970 326898 215206 327134
rect 245690 327218 245926 327454
rect 245690 326898 245926 327134
rect 276410 327218 276646 327454
rect 276410 326898 276646 327134
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 199610 295718 199846 295954
rect 199610 295398 199846 295634
rect 230330 295718 230566 295954
rect 230330 295398 230566 295634
rect 261050 295718 261286 295954
rect 261050 295398 261286 295634
rect 184250 291218 184486 291454
rect 184250 290898 184486 291134
rect 214970 291218 215206 291454
rect 214970 290898 215206 291134
rect 245690 291218 245926 291454
rect 245690 290898 245926 291134
rect 276410 291218 276646 291454
rect 276410 290898 276646 291134
rect 199610 259718 199846 259954
rect 199610 259398 199846 259634
rect 230330 259718 230566 259954
rect 230330 259398 230566 259634
rect 261050 259718 261286 259954
rect 261050 259398 261286 259634
rect 184250 255218 184486 255454
rect 184250 254898 184486 255134
rect 214970 255218 215206 255454
rect 214970 254898 215206 255134
rect 245690 255218 245926 255454
rect 245690 254898 245926 255134
rect 276410 255218 276646 255454
rect 276410 254898 276646 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 227916 151718 228152 151954
rect 227916 151398 228152 151634
rect 237847 151718 238083 151954
rect 237847 151398 238083 151634
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 227916 115718 228152 115954
rect 227916 115398 228152 115634
rect 237847 115718 238083 115954
rect 237847 115398 238083 115634
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 242813 110898 243049 111134
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 314250 151718 314486 151954
rect 314250 151398 314486 151634
rect 317514 151718 317750 151954
rect 317514 151398 317750 151634
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 314250 115718 314486 115954
rect 314250 115398 314486 115634
rect 317514 115718 317750 115954
rect 317514 115398 317750 115634
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 359610 583718 359846 583954
rect 359610 583398 359846 583634
rect 390330 583718 390566 583954
rect 390330 583398 390566 583634
rect 421050 583718 421286 583954
rect 421050 583398 421286 583634
rect 451770 583718 452006 583954
rect 451770 583398 452006 583634
rect 482490 583718 482726 583954
rect 482490 583398 482726 583634
rect 513210 583718 513446 583954
rect 513210 583398 513446 583634
rect 344250 579218 344486 579454
rect 344250 578898 344486 579134
rect 374970 579218 375206 579454
rect 374970 578898 375206 579134
rect 405690 579218 405926 579454
rect 405690 578898 405926 579134
rect 436410 579218 436646 579454
rect 436410 578898 436646 579134
rect 467130 579218 467366 579454
rect 467130 578898 467366 579134
rect 497850 579218 498086 579454
rect 497850 578898 498086 579134
rect 528570 579218 528806 579454
rect 528570 578898 528806 579134
rect 359610 547718 359846 547954
rect 359610 547398 359846 547634
rect 390330 547718 390566 547954
rect 390330 547398 390566 547634
rect 421050 547718 421286 547954
rect 421050 547398 421286 547634
rect 451770 547718 452006 547954
rect 451770 547398 452006 547634
rect 482490 547718 482726 547954
rect 482490 547398 482726 547634
rect 513210 547718 513446 547954
rect 513210 547398 513446 547634
rect 344250 543218 344486 543454
rect 344250 542898 344486 543134
rect 374970 543218 375206 543454
rect 374970 542898 375206 543134
rect 405690 543218 405926 543454
rect 405690 542898 405926 543134
rect 436410 543218 436646 543454
rect 436410 542898 436646 543134
rect 467130 543218 467366 543454
rect 467130 542898 467366 543134
rect 497850 543218 498086 543454
rect 497850 542898 498086 543134
rect 528570 543218 528806 543454
rect 528570 542898 528806 543134
rect 359610 511718 359846 511954
rect 359610 511398 359846 511634
rect 390330 511718 390566 511954
rect 390330 511398 390566 511634
rect 421050 511718 421286 511954
rect 421050 511398 421286 511634
rect 451770 511718 452006 511954
rect 451770 511398 452006 511634
rect 482490 511718 482726 511954
rect 482490 511398 482726 511634
rect 513210 511718 513446 511954
rect 513210 511398 513446 511634
rect 344250 507218 344486 507454
rect 344250 506898 344486 507134
rect 374970 507218 375206 507454
rect 374970 506898 375206 507134
rect 405690 507218 405926 507454
rect 405690 506898 405926 507134
rect 436410 507218 436646 507454
rect 436410 506898 436646 507134
rect 467130 507218 467366 507454
rect 467130 506898 467366 507134
rect 497850 507218 498086 507454
rect 497850 506898 498086 507134
rect 528570 507218 528806 507454
rect 528570 506898 528806 507134
rect 359610 475718 359846 475954
rect 359610 475398 359846 475634
rect 390330 475718 390566 475954
rect 390330 475398 390566 475634
rect 421050 475718 421286 475954
rect 421050 475398 421286 475634
rect 451770 475718 452006 475954
rect 451770 475398 452006 475634
rect 482490 475718 482726 475954
rect 482490 475398 482726 475634
rect 513210 475718 513446 475954
rect 513210 475398 513446 475634
rect 344250 471218 344486 471454
rect 344250 470898 344486 471134
rect 374970 471218 375206 471454
rect 374970 470898 375206 471134
rect 405690 471218 405926 471454
rect 405690 470898 405926 471134
rect 436410 471218 436646 471454
rect 436410 470898 436646 471134
rect 467130 471218 467366 471454
rect 467130 470898 467366 471134
rect 497850 471218 498086 471454
rect 497850 470898 498086 471134
rect 528570 471218 528806 471454
rect 528570 470898 528806 471134
rect 359610 439718 359846 439954
rect 359610 439398 359846 439634
rect 390330 439718 390566 439954
rect 390330 439398 390566 439634
rect 421050 439718 421286 439954
rect 421050 439398 421286 439634
rect 451770 439718 452006 439954
rect 451770 439398 452006 439634
rect 482490 439718 482726 439954
rect 482490 439398 482726 439634
rect 513210 439718 513446 439954
rect 513210 439398 513446 439634
rect 344250 435218 344486 435454
rect 344250 434898 344486 435134
rect 374970 435218 375206 435454
rect 374970 434898 375206 435134
rect 405690 435218 405926 435454
rect 405690 434898 405926 435134
rect 436410 435218 436646 435454
rect 436410 434898 436646 435134
rect 467130 435218 467366 435454
rect 467130 434898 467366 435134
rect 497850 435218 498086 435454
rect 497850 434898 498086 435134
rect 528570 435218 528806 435454
rect 528570 434898 528806 435134
rect 359610 403718 359846 403954
rect 359610 403398 359846 403634
rect 390330 403718 390566 403954
rect 390330 403398 390566 403634
rect 421050 403718 421286 403954
rect 421050 403398 421286 403634
rect 451770 403718 452006 403954
rect 451770 403398 452006 403634
rect 482490 403718 482726 403954
rect 482490 403398 482726 403634
rect 513210 403718 513446 403954
rect 513210 403398 513446 403634
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 399610 295718 399846 295954
rect 399610 295398 399846 295634
rect 430330 295718 430566 295954
rect 430330 295398 430566 295634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 384250 291218 384486 291454
rect 384250 290898 384486 291134
rect 414970 291218 415206 291454
rect 414970 290898 415206 291134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 399610 259718 399846 259954
rect 399610 259398 399846 259634
rect 430330 259718 430566 259954
rect 430330 259398 430566 259634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 384250 255218 384486 255454
rect 384250 254898 384486 255134
rect 414970 255218 415206 255454
rect 414970 254898 415206 255134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 419610 115718 419846 115954
rect 419610 115398 419846 115634
rect 404250 111218 404486 111454
rect 404250 110898 404486 111134
rect 434970 111218 435206 111454
rect 434970 110898 435206 111134
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 359610 583954
rect 359846 583718 390330 583954
rect 390566 583718 421050 583954
rect 421286 583718 451770 583954
rect 452006 583718 482490 583954
rect 482726 583718 513210 583954
rect 513446 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 359610 583634
rect 359846 583398 390330 583634
rect 390566 583398 421050 583634
rect 421286 583398 451770 583634
rect 452006 583398 482490 583634
rect 482726 583398 513210 583634
rect 513446 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 68250 579454
rect 68486 579218 98970 579454
rect 99206 579218 129690 579454
rect 129926 579218 160410 579454
rect 160646 579218 191130 579454
rect 191366 579218 221850 579454
rect 222086 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 344250 579454
rect 344486 579218 374970 579454
rect 375206 579218 405690 579454
rect 405926 579218 436410 579454
rect 436646 579218 467130 579454
rect 467366 579218 497850 579454
rect 498086 579218 528570 579454
rect 528806 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 68250 579134
rect 68486 578898 98970 579134
rect 99206 578898 129690 579134
rect 129926 578898 160410 579134
rect 160646 578898 191130 579134
rect 191366 578898 221850 579134
rect 222086 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 344250 579134
rect 344486 578898 374970 579134
rect 375206 578898 405690 579134
rect 405926 578898 436410 579134
rect 436646 578898 467130 579134
rect 467366 578898 497850 579134
rect 498086 578898 528570 579134
rect 528806 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 83610 547954
rect 83846 547718 114330 547954
rect 114566 547718 145050 547954
rect 145286 547718 175770 547954
rect 176006 547718 206490 547954
rect 206726 547718 237210 547954
rect 237446 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 359610 547954
rect 359846 547718 390330 547954
rect 390566 547718 421050 547954
rect 421286 547718 451770 547954
rect 452006 547718 482490 547954
rect 482726 547718 513210 547954
rect 513446 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 83610 547634
rect 83846 547398 114330 547634
rect 114566 547398 145050 547634
rect 145286 547398 175770 547634
rect 176006 547398 206490 547634
rect 206726 547398 237210 547634
rect 237446 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 359610 547634
rect 359846 547398 390330 547634
rect 390566 547398 421050 547634
rect 421286 547398 451770 547634
rect 452006 547398 482490 547634
rect 482726 547398 513210 547634
rect 513446 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 68250 543454
rect 68486 543218 98970 543454
rect 99206 543218 129690 543454
rect 129926 543218 160410 543454
rect 160646 543218 191130 543454
rect 191366 543218 221850 543454
rect 222086 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 344250 543454
rect 344486 543218 374970 543454
rect 375206 543218 405690 543454
rect 405926 543218 436410 543454
rect 436646 543218 467130 543454
rect 467366 543218 497850 543454
rect 498086 543218 528570 543454
rect 528806 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 68250 543134
rect 68486 542898 98970 543134
rect 99206 542898 129690 543134
rect 129926 542898 160410 543134
rect 160646 542898 191130 543134
rect 191366 542898 221850 543134
rect 222086 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 344250 543134
rect 344486 542898 374970 543134
rect 375206 542898 405690 543134
rect 405926 542898 436410 543134
rect 436646 542898 467130 543134
rect 467366 542898 497850 543134
rect 498086 542898 528570 543134
rect 528806 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 83610 511954
rect 83846 511718 114330 511954
rect 114566 511718 145050 511954
rect 145286 511718 175770 511954
rect 176006 511718 206490 511954
rect 206726 511718 237210 511954
rect 237446 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 359610 511954
rect 359846 511718 390330 511954
rect 390566 511718 421050 511954
rect 421286 511718 451770 511954
rect 452006 511718 482490 511954
rect 482726 511718 513210 511954
rect 513446 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 83610 511634
rect 83846 511398 114330 511634
rect 114566 511398 145050 511634
rect 145286 511398 175770 511634
rect 176006 511398 206490 511634
rect 206726 511398 237210 511634
rect 237446 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 359610 511634
rect 359846 511398 390330 511634
rect 390566 511398 421050 511634
rect 421286 511398 451770 511634
rect 452006 511398 482490 511634
rect 482726 511398 513210 511634
rect 513446 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 68250 507454
rect 68486 507218 98970 507454
rect 99206 507218 129690 507454
rect 129926 507218 160410 507454
rect 160646 507218 191130 507454
rect 191366 507218 221850 507454
rect 222086 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 344250 507454
rect 344486 507218 374970 507454
rect 375206 507218 405690 507454
rect 405926 507218 436410 507454
rect 436646 507218 467130 507454
rect 467366 507218 497850 507454
rect 498086 507218 528570 507454
rect 528806 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 68250 507134
rect 68486 506898 98970 507134
rect 99206 506898 129690 507134
rect 129926 506898 160410 507134
rect 160646 506898 191130 507134
rect 191366 506898 221850 507134
rect 222086 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 344250 507134
rect 344486 506898 374970 507134
rect 375206 506898 405690 507134
rect 405926 506898 436410 507134
rect 436646 506898 467130 507134
rect 467366 506898 497850 507134
rect 498086 506898 528570 507134
rect 528806 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 83610 475954
rect 83846 475718 114330 475954
rect 114566 475718 145050 475954
rect 145286 475718 175770 475954
rect 176006 475718 206490 475954
rect 206726 475718 237210 475954
rect 237446 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 359610 475954
rect 359846 475718 390330 475954
rect 390566 475718 421050 475954
rect 421286 475718 451770 475954
rect 452006 475718 482490 475954
rect 482726 475718 513210 475954
rect 513446 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 83610 475634
rect 83846 475398 114330 475634
rect 114566 475398 145050 475634
rect 145286 475398 175770 475634
rect 176006 475398 206490 475634
rect 206726 475398 237210 475634
rect 237446 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 359610 475634
rect 359846 475398 390330 475634
rect 390566 475398 421050 475634
rect 421286 475398 451770 475634
rect 452006 475398 482490 475634
rect 482726 475398 513210 475634
rect 513446 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 68250 471454
rect 68486 471218 98970 471454
rect 99206 471218 129690 471454
rect 129926 471218 160410 471454
rect 160646 471218 191130 471454
rect 191366 471218 221850 471454
rect 222086 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 344250 471454
rect 344486 471218 374970 471454
rect 375206 471218 405690 471454
rect 405926 471218 436410 471454
rect 436646 471218 467130 471454
rect 467366 471218 497850 471454
rect 498086 471218 528570 471454
rect 528806 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 68250 471134
rect 68486 470898 98970 471134
rect 99206 470898 129690 471134
rect 129926 470898 160410 471134
rect 160646 470898 191130 471134
rect 191366 470898 221850 471134
rect 222086 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 344250 471134
rect 344486 470898 374970 471134
rect 375206 470898 405690 471134
rect 405926 470898 436410 471134
rect 436646 470898 467130 471134
rect 467366 470898 497850 471134
rect 498086 470898 528570 471134
rect 528806 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 83610 439954
rect 83846 439718 114330 439954
rect 114566 439718 145050 439954
rect 145286 439718 175770 439954
rect 176006 439718 206490 439954
rect 206726 439718 237210 439954
rect 237446 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 359610 439954
rect 359846 439718 390330 439954
rect 390566 439718 421050 439954
rect 421286 439718 451770 439954
rect 452006 439718 482490 439954
rect 482726 439718 513210 439954
rect 513446 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 83610 439634
rect 83846 439398 114330 439634
rect 114566 439398 145050 439634
rect 145286 439398 175770 439634
rect 176006 439398 206490 439634
rect 206726 439398 237210 439634
rect 237446 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 359610 439634
rect 359846 439398 390330 439634
rect 390566 439398 421050 439634
rect 421286 439398 451770 439634
rect 452006 439398 482490 439634
rect 482726 439398 513210 439634
rect 513446 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 68250 435454
rect 68486 435218 98970 435454
rect 99206 435218 129690 435454
rect 129926 435218 160410 435454
rect 160646 435218 191130 435454
rect 191366 435218 221850 435454
rect 222086 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 344250 435454
rect 344486 435218 374970 435454
rect 375206 435218 405690 435454
rect 405926 435218 436410 435454
rect 436646 435218 467130 435454
rect 467366 435218 497850 435454
rect 498086 435218 528570 435454
rect 528806 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 68250 435134
rect 68486 434898 98970 435134
rect 99206 434898 129690 435134
rect 129926 434898 160410 435134
rect 160646 434898 191130 435134
rect 191366 434898 221850 435134
rect 222086 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 344250 435134
rect 344486 434898 374970 435134
rect 375206 434898 405690 435134
rect 405926 434898 436410 435134
rect 436646 434898 467130 435134
rect 467366 434898 497850 435134
rect 498086 434898 528570 435134
rect 528806 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 359610 403954
rect 359846 403718 390330 403954
rect 390566 403718 421050 403954
rect 421286 403718 451770 403954
rect 452006 403718 482490 403954
rect 482726 403718 513210 403954
rect 513446 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 359610 403634
rect 359846 403398 390330 403634
rect 390566 403398 421050 403634
rect 421286 403398 451770 403634
rect 452006 403398 482490 403634
rect 482726 403398 513210 403634
rect 513446 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 199610 331954
rect 199846 331718 230330 331954
rect 230566 331718 261050 331954
rect 261286 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 199610 331634
rect 199846 331398 230330 331634
rect 230566 331398 261050 331634
rect 261286 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 184250 327454
rect 184486 327218 214970 327454
rect 215206 327218 245690 327454
rect 245926 327218 276410 327454
rect 276646 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 184250 327134
rect 184486 326898 214970 327134
rect 215206 326898 245690 327134
rect 245926 326898 276410 327134
rect 276646 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 199610 295954
rect 199846 295718 230330 295954
rect 230566 295718 261050 295954
rect 261286 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 399610 295954
rect 399846 295718 430330 295954
rect 430566 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 199610 295634
rect 199846 295398 230330 295634
rect 230566 295398 261050 295634
rect 261286 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 399610 295634
rect 399846 295398 430330 295634
rect 430566 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 184250 291454
rect 184486 291218 214970 291454
rect 215206 291218 245690 291454
rect 245926 291218 276410 291454
rect 276646 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 384250 291454
rect 384486 291218 414970 291454
rect 415206 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 184250 291134
rect 184486 290898 214970 291134
rect 215206 290898 245690 291134
rect 245926 290898 276410 291134
rect 276646 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 384250 291134
rect 384486 290898 414970 291134
rect 415206 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 89610 259954
rect 89846 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 199610 259954
rect 199846 259718 230330 259954
rect 230566 259718 261050 259954
rect 261286 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 399610 259954
rect 399846 259718 430330 259954
rect 430566 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 89610 259634
rect 89846 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 199610 259634
rect 199846 259398 230330 259634
rect 230566 259398 261050 259634
rect 261286 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 399610 259634
rect 399846 259398 430330 259634
rect 430566 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 184250 255454
rect 184486 255218 214970 255454
rect 215206 255218 245690 255454
rect 245926 255218 276410 255454
rect 276646 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 384250 255454
rect 384486 255218 414970 255454
rect 415206 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 184250 255134
rect 184486 254898 214970 255134
rect 215206 254898 245690 255134
rect 245926 254898 276410 255134
rect 276646 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 384250 255134
rect 384486 254898 414970 255134
rect 415206 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 69128 151954
rect 69364 151718 164192 151954
rect 164428 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 227916 151954
rect 228152 151718 237847 151954
rect 238083 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 314250 151954
rect 314486 151718 317514 151954
rect 317750 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 69128 151634
rect 69364 151398 164192 151634
rect 164428 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 227916 151634
rect 228152 151398 237847 151634
rect 238083 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 314250 151634
rect 314486 151398 317514 151634
rect 317750 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 69128 115954
rect 69364 115718 164192 115954
rect 164428 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 227916 115954
rect 228152 115718 237847 115954
rect 238083 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 314250 115954
rect 314486 115718 317514 115954
rect 317750 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 419610 115954
rect 419846 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 69128 115634
rect 69364 115398 164192 115634
rect 164428 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 227916 115634
rect 228152 115398 237847 115634
rect 238083 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 314250 115634
rect 314486 115398 317514 115634
rect 317750 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 419610 115634
rect 419846 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 404250 111454
rect 404486 111218 434970 111454
rect 435206 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 404250 111134
rect 404486 110898 434970 111134
rect 435206 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_etpu  wrapped_etpu_3
timestamp 0
transform 1 0 64000 0 1 405000
box -10 0 180000 180000
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
use wrapped_ibnalhaytham  wrapped_ibnalhaytham_1
timestamp 0
transform 1 0 180000 0 1 240000
box 0 0 113010 115154
use wrapped_mbsFSK  wrapped_mbsFSK_5
timestamp 0
transform 1 0 400000 0 1 96000
box -10 -52 50000 50000
use wrapped_silife  wrapped_silife_2
timestamp 0
transform 1 0 340000 0 1 400000
box 0 0 193294 195438
use wrapped_snn_network  wrapped_snn_network_4
timestamp 0
transform 1 0 380000 0 1 240000
box -10 -52 60000 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 176600 74414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 294000 74414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 587000 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 176600 110414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 294000 110414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 587000 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 176600 146414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 587000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 357154 182414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 587000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 178000 218414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 357154 218414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 587000 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 357154 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 357154 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 597438 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 148000 398414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 302000 398414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 597438 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 148000 434414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 302000 434414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 597438 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 597438 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 597438 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 176600 83414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 294000 83414 403000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 587000 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 176600 119414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 294000 119414 403000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 587000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 176600 155414 403000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 587000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 587000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 178000 227414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 587000 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 357154 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 597438 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 148000 407414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 302000 407414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 597438 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 148000 443414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 597438 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 597438 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 597438 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 176600 92414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 294000 92414 403000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 587000 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 176600 128414 403000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 587000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 176600 164414 403000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 587000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 587000 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 178000 236414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 587000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 357154 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 178000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 597438 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 302000 380414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 597438 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 148000 416414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 302000 416414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 597438 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 148000 452414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 597438 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 597438 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 597438 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 403000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 587000 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 294000 101414 403000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 587000 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 176600 137414 403000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 587000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 403000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 587000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 587000 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 587000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 357154 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 178000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 597438 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 302000 389414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 597438 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 148000 425414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 302000 425414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 597438 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 597438 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 597438 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 597438 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 294000 96914 403000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 587000 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 176600 132914 403000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 587000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 403000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 587000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 587000 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 587000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 357154 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 178000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 597438 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 302000 384914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 597438 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 148000 420914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 302000 420914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 597438 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 597438 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 597438 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 597438 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 176600 69914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 294000 69914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 587000 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 176600 105914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 294000 105914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 587000 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 176600 141914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 587000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 587000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 357154 213914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 587000 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 178000 249914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 357154 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 357154 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 178000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 597438 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 302000 393914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 597438 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 148000 429914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 302000 429914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 597438 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 597438 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 597438 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 176600 78914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 294000 78914 403000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 587000 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 176600 114914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 294000 114914 403000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 587000 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 176600 150914 403000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 587000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 587000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 178000 222914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 587000 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 357154 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 357154 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 597438 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 148000 402914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 302000 402914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 597438 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 148000 438914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 302000 438914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 597438 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 597438 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 597438 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 176600 87914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 294000 87914 403000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 587000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 176600 123914 403000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 587000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 176600 159914 403000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 587000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 587000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 178000 231914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 587000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 357154 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 597438 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 597438 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 148000 411914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 302000 411914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 597438 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 148000 447914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 597438 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 597438 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 597438 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
