VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_silife
  CLASS BLOCK ;
  FOREIGN wrapped_silife ;
  ORIGIN 0.000 0.000 ;
  SIZE 966.470 BY 977.190 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 907.840 966.470 908.440 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 973.190 254.750 977.190 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 973.190 303.050 977.190 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 973.190 889.090 977.190 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 894.240 966.470 894.840 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 973.190 435.070 977.190 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 265.240 966.470 265.840 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 744.640 966.470 745.240 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 112.240 966.470 112.840 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 973.190 171.030 977.190 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 973.190 505.910 977.190 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 856.840 966.470 857.440 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 377.440 966.470 378.040 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 973.190 148.490 977.190 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 973.190 686.230 977.190 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 973.190 579.970 977.190 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 973.190 135.610 977.190 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 958.840 966.470 959.440 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 973.190 818.250 977.190 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 973.190 734.530 977.190 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 768.440 966.470 769.040 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 530.440 966.470 531.040 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 37.440 966.470 38.040 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 973.190 87.310 977.190 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 353.640 966.470 354.240 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 973.190 386.770 977.190 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 973.190 267.630 977.190 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 605.240 966.470 605.840 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 136.040 966.470 136.640 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 656.240 966.470 656.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 973.190 280.510 977.190 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 973.190 805.370 977.190 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 666.440 966.470 667.040 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 149.640 966.470 150.240 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 340.040 966.470 340.640 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 973.190 377.110 977.190 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 973.190 412.530 977.190 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 74.840 966.470 75.440 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 567.840 966.470 568.440 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 973.190 183.910 977.190 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 591.640 966.470 592.240 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 972.440 966.470 973.040 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 973.190 399.650 977.190 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 754.840 966.470 755.440 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 973.190 747.410 977.190 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 973.190 937.390 977.190 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 973.190 209.670 977.190 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 312.840 966.470 313.440 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 973.190 628.270 977.190 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 973.190 950.270 977.190 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 10.240 966.470 10.840 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 326.440 966.470 327.040 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 973.190 42.230 977.190 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 452.240 966.470 452.840 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 973.190 496.250 977.190 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 973.190 663.690 977.190 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 833.040 966.470 833.640 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 973.190 518.790 977.190 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 973.190 602.510 977.190 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 618.840 966.470 619.440 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 275.440 966.470 276.040 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 973.190 232.210 977.190 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 973.190 29.350 977.190 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 88.440 966.470 89.040 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 717.440 966.470 718.040 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 973.190 914.850 977.190 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 973.190 293.390 977.190 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 973.190 196.790 977.190 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 401.240 966.470 401.840 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 931.640 966.470 932.240 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 554.240 966.470 554.840 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 973.190 447.950 977.190 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 125.840 966.470 126.440 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 47.640 966.470 48.240 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 973.190 460.830 977.190 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 200.640 966.470 201.240 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 214.240 966.470 214.840 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 973.190 769.950 977.190 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 973.190 315.930 977.190 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 642.640 966.470 643.240 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 795.640 966.470 796.240 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 973.190 422.190 977.190 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 973.190 3.590 977.190 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 973.190 161.370 977.190 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 578.040 966.470 578.640 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 629.040 966.470 629.640 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 973.190 853.670 977.190 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 479.440 966.470 480.040 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 973.190 721.650 977.190 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 693.640 966.470 694.240 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 973.190 531.670 977.190 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 251.640 966.470 252.240 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 973.190 673.350 977.190 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 391.040 966.470 391.640 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 973.190 963.150 977.190 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 289.040 966.470 289.640 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 819.440 966.470 820.040 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 973.190 866.550 977.190 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 973.190 567.090 977.190 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 973.190 64.770 977.190 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 973.190 589.630 977.190 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 884.040 966.470 884.640 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 973.190 245.090 977.190 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 973.190 77.650 977.190 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 973.190 615.390 977.190 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 965.840 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 965.840 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 23.840 966.470 24.440 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 973.190 470.490 977.190 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 187.040 966.470 187.640 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 973.190 879.430 977.190 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 973.190 699.110 977.190 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 973.190 113.070 977.190 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 973.190 100.190 977.190 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 540.640 966.470 541.240 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 489.640 966.470 490.240 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 428.440 966.470 429.040 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 176.840 966.470 177.440 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 973.190 831.130 977.190 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 870.440 966.470 871.040 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 98.640 966.470 99.240 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 973.190 351.350 977.190 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 973.190 544.550 977.190 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 442.040 966.470 442.640 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 782.040 966.470 782.640 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 973.190 924.510 977.190 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 302.640 966.470 303.240 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 163.240 966.470 163.840 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 973.190 483.370 977.190 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 973.190 51.890 977.190 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 973.190 16.470 977.190 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 414.840 966.470 415.440 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 973.190 782.830 977.190 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 945.240 966.470 945.840 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 973.190 219.330 977.190 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 921.440 966.470 922.040 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 680.040 966.470 680.640 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 973.190 901.970 977.190 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 973.190 364.230 977.190 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 516.840 966.470 517.440 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 224.440 966.470 225.040 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 363.840 966.470 364.440 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 973.190 840.790 977.190 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 805.840 966.470 806.440 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 0.040 966.470 0.640 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 503.240 966.470 503.840 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 843.240 966.470 843.840 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 973.190 795.710 977.190 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 61.240 966.470 61.840 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 973.190 757.070 977.190 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 973.190 328.810 977.190 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 973.190 554.210 977.190 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 973.190 338.470 977.190 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 973.190 711.990 977.190 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 238.040 966.470 238.640 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 731.040 966.470 731.640 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 707.240 966.470 707.840 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 973.190 650.810 977.190 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 973.190 637.930 977.190 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 973.190 125.950 977.190 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 962.470 465.840 966.470 466.440 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 960.940 965.685 ;
      LAYER met1 ;
        RECT 0.070 0.040 966.390 969.300 ;
      LAYER met2 ;
        RECT 0.100 972.910 3.030 973.490 ;
        RECT 3.870 972.910 15.910 973.490 ;
        RECT 16.750 972.910 28.790 973.490 ;
        RECT 29.630 972.910 41.670 973.490 ;
        RECT 42.510 972.910 51.330 973.490 ;
        RECT 52.170 972.910 64.210 973.490 ;
        RECT 65.050 972.910 77.090 973.490 ;
        RECT 77.930 972.910 86.750 973.490 ;
        RECT 87.590 972.910 99.630 973.490 ;
        RECT 100.470 972.910 112.510 973.490 ;
        RECT 113.350 972.910 125.390 973.490 ;
        RECT 126.230 972.910 135.050 973.490 ;
        RECT 135.890 972.910 147.930 973.490 ;
        RECT 148.770 972.910 160.810 973.490 ;
        RECT 161.650 972.910 170.470 973.490 ;
        RECT 171.310 972.910 183.350 973.490 ;
        RECT 184.190 972.910 196.230 973.490 ;
        RECT 197.070 972.910 209.110 973.490 ;
        RECT 209.950 972.910 218.770 973.490 ;
        RECT 219.610 972.910 231.650 973.490 ;
        RECT 232.490 972.910 244.530 973.490 ;
        RECT 245.370 972.910 254.190 973.490 ;
        RECT 255.030 972.910 267.070 973.490 ;
        RECT 267.910 972.910 279.950 973.490 ;
        RECT 280.790 972.910 292.830 973.490 ;
        RECT 293.670 972.910 302.490 973.490 ;
        RECT 303.330 972.910 315.370 973.490 ;
        RECT 316.210 972.910 328.250 973.490 ;
        RECT 329.090 972.910 337.910 973.490 ;
        RECT 338.750 972.910 350.790 973.490 ;
        RECT 351.630 972.910 363.670 973.490 ;
        RECT 364.510 972.910 376.550 973.490 ;
        RECT 377.390 972.910 386.210 973.490 ;
        RECT 387.050 972.910 399.090 973.490 ;
        RECT 399.930 972.910 411.970 973.490 ;
        RECT 412.810 972.910 421.630 973.490 ;
        RECT 422.470 972.910 434.510 973.490 ;
        RECT 435.350 972.910 447.390 973.490 ;
        RECT 448.230 972.910 460.270 973.490 ;
        RECT 461.110 972.910 469.930 973.490 ;
        RECT 470.770 972.910 482.810 973.490 ;
        RECT 483.650 972.910 495.690 973.490 ;
        RECT 496.530 972.910 505.350 973.490 ;
        RECT 506.190 972.910 518.230 973.490 ;
        RECT 519.070 972.910 531.110 973.490 ;
        RECT 531.950 972.910 543.990 973.490 ;
        RECT 544.830 972.910 553.650 973.490 ;
        RECT 554.490 972.910 566.530 973.490 ;
        RECT 567.370 972.910 579.410 973.490 ;
        RECT 580.250 972.910 589.070 973.490 ;
        RECT 589.910 972.910 601.950 973.490 ;
        RECT 602.790 972.910 614.830 973.490 ;
        RECT 615.670 972.910 627.710 973.490 ;
        RECT 628.550 972.910 637.370 973.490 ;
        RECT 638.210 972.910 650.250 973.490 ;
        RECT 651.090 972.910 663.130 973.490 ;
        RECT 663.970 972.910 672.790 973.490 ;
        RECT 673.630 972.910 685.670 973.490 ;
        RECT 686.510 972.910 698.550 973.490 ;
        RECT 699.390 972.910 711.430 973.490 ;
        RECT 712.270 972.910 721.090 973.490 ;
        RECT 721.930 972.910 733.970 973.490 ;
        RECT 734.810 972.910 746.850 973.490 ;
        RECT 747.690 972.910 756.510 973.490 ;
        RECT 757.350 972.910 769.390 973.490 ;
        RECT 770.230 972.910 782.270 973.490 ;
        RECT 783.110 972.910 795.150 973.490 ;
        RECT 795.990 972.910 804.810 973.490 ;
        RECT 805.650 972.910 817.690 973.490 ;
        RECT 818.530 972.910 830.570 973.490 ;
        RECT 831.410 972.910 840.230 973.490 ;
        RECT 841.070 972.910 853.110 973.490 ;
        RECT 853.950 972.910 865.990 973.490 ;
        RECT 866.830 972.910 878.870 973.490 ;
        RECT 879.710 972.910 888.530 973.490 ;
        RECT 889.370 972.910 901.410 973.490 ;
        RECT 902.250 972.910 914.290 973.490 ;
        RECT 915.130 972.910 923.950 973.490 ;
        RECT 924.790 972.910 936.830 973.490 ;
        RECT 937.670 972.910 949.710 973.490 ;
        RECT 950.550 972.910 962.590 973.490 ;
        RECT 963.430 972.910 966.370 973.490 ;
        RECT 0.100 4.280 966.370 972.910 ;
        RECT 0.650 0.010 9.470 4.280 ;
        RECT 10.310 0.010 22.350 4.280 ;
        RECT 23.190 0.010 35.230 4.280 ;
        RECT 36.070 0.010 44.890 4.280 ;
        RECT 45.730 0.010 57.770 4.280 ;
        RECT 58.610 0.010 70.650 4.280 ;
        RECT 71.490 0.010 83.530 4.280 ;
        RECT 84.370 0.010 93.190 4.280 ;
        RECT 94.030 0.010 106.070 4.280 ;
        RECT 106.910 0.010 118.950 4.280 ;
        RECT 119.790 0.010 128.610 4.280 ;
        RECT 129.450 0.010 141.490 4.280 ;
        RECT 142.330 0.010 154.370 4.280 ;
        RECT 155.210 0.010 167.250 4.280 ;
        RECT 168.090 0.010 176.910 4.280 ;
        RECT 177.750 0.010 189.790 4.280 ;
        RECT 190.630 0.010 202.670 4.280 ;
        RECT 203.510 0.010 212.330 4.280 ;
        RECT 213.170 0.010 225.210 4.280 ;
        RECT 226.050 0.010 238.090 4.280 ;
        RECT 238.930 0.010 250.970 4.280 ;
        RECT 251.810 0.010 260.630 4.280 ;
        RECT 261.470 0.010 273.510 4.280 ;
        RECT 274.350 0.010 286.390 4.280 ;
        RECT 287.230 0.010 296.050 4.280 ;
        RECT 296.890 0.010 308.930 4.280 ;
        RECT 309.770 0.010 321.810 4.280 ;
        RECT 322.650 0.010 334.690 4.280 ;
        RECT 335.530 0.010 344.350 4.280 ;
        RECT 345.190 0.010 357.230 4.280 ;
        RECT 358.070 0.010 370.110 4.280 ;
        RECT 370.950 0.010 379.770 4.280 ;
        RECT 380.610 0.010 392.650 4.280 ;
        RECT 393.490 0.010 405.530 4.280 ;
        RECT 406.370 0.010 418.410 4.280 ;
        RECT 419.250 0.010 428.070 4.280 ;
        RECT 428.910 0.010 440.950 4.280 ;
        RECT 441.790 0.010 453.830 4.280 ;
        RECT 454.670 0.010 463.490 4.280 ;
        RECT 464.330 0.010 476.370 4.280 ;
        RECT 477.210 0.010 489.250 4.280 ;
        RECT 490.090 0.010 502.130 4.280 ;
        RECT 502.970 0.010 511.790 4.280 ;
        RECT 512.630 0.010 524.670 4.280 ;
        RECT 525.510 0.010 537.550 4.280 ;
        RECT 538.390 0.010 547.210 4.280 ;
        RECT 548.050 0.010 560.090 4.280 ;
        RECT 560.930 0.010 572.970 4.280 ;
        RECT 573.810 0.010 585.850 4.280 ;
        RECT 586.690 0.010 595.510 4.280 ;
        RECT 596.350 0.010 608.390 4.280 ;
        RECT 609.230 0.010 621.270 4.280 ;
        RECT 622.110 0.010 630.930 4.280 ;
        RECT 631.770 0.010 643.810 4.280 ;
        RECT 644.650 0.010 656.690 4.280 ;
        RECT 657.530 0.010 669.570 4.280 ;
        RECT 670.410 0.010 679.230 4.280 ;
        RECT 680.070 0.010 692.110 4.280 ;
        RECT 692.950 0.010 704.990 4.280 ;
        RECT 705.830 0.010 714.650 4.280 ;
        RECT 715.490 0.010 727.530 4.280 ;
        RECT 728.370 0.010 740.410 4.280 ;
        RECT 741.250 0.010 753.290 4.280 ;
        RECT 754.130 0.010 762.950 4.280 ;
        RECT 763.790 0.010 775.830 4.280 ;
        RECT 776.670 0.010 788.710 4.280 ;
        RECT 789.550 0.010 798.370 4.280 ;
        RECT 799.210 0.010 811.250 4.280 ;
        RECT 812.090 0.010 824.130 4.280 ;
        RECT 824.970 0.010 837.010 4.280 ;
        RECT 837.850 0.010 846.670 4.280 ;
        RECT 847.510 0.010 859.550 4.280 ;
        RECT 860.390 0.010 872.430 4.280 ;
        RECT 873.270 0.010 882.090 4.280 ;
        RECT 882.930 0.010 894.970 4.280 ;
        RECT 895.810 0.010 907.850 4.280 ;
        RECT 908.690 0.010 920.730 4.280 ;
        RECT 921.570 0.010 930.390 4.280 ;
        RECT 931.230 0.010 943.270 4.280 ;
        RECT 944.110 0.010 956.150 4.280 ;
        RECT 956.990 0.010 966.370 4.280 ;
      LAYER met3 ;
        RECT 4.400 972.040 962.070 972.905 ;
        RECT 3.990 959.840 966.395 972.040 ;
        RECT 4.400 958.440 962.070 959.840 ;
        RECT 3.990 946.240 966.395 958.440 ;
        RECT 4.400 944.840 962.070 946.240 ;
        RECT 3.990 932.640 966.395 944.840 ;
        RECT 4.400 931.240 962.070 932.640 ;
        RECT 3.990 922.440 966.395 931.240 ;
        RECT 4.400 921.040 962.070 922.440 ;
        RECT 3.990 908.840 966.395 921.040 ;
        RECT 4.400 907.440 962.070 908.840 ;
        RECT 3.990 895.240 966.395 907.440 ;
        RECT 4.400 893.840 962.070 895.240 ;
        RECT 3.990 885.040 966.395 893.840 ;
        RECT 4.400 883.640 962.070 885.040 ;
        RECT 3.990 871.440 966.395 883.640 ;
        RECT 4.400 870.040 962.070 871.440 ;
        RECT 3.990 857.840 966.395 870.040 ;
        RECT 4.400 856.440 962.070 857.840 ;
        RECT 3.990 844.240 966.395 856.440 ;
        RECT 4.400 842.840 962.070 844.240 ;
        RECT 3.990 834.040 966.395 842.840 ;
        RECT 4.400 832.640 962.070 834.040 ;
        RECT 3.990 820.440 966.395 832.640 ;
        RECT 4.400 819.040 962.070 820.440 ;
        RECT 3.990 806.840 966.395 819.040 ;
        RECT 4.400 805.440 962.070 806.840 ;
        RECT 3.990 796.640 966.395 805.440 ;
        RECT 4.400 795.240 962.070 796.640 ;
        RECT 3.990 783.040 966.395 795.240 ;
        RECT 4.400 781.640 962.070 783.040 ;
        RECT 3.990 769.440 966.395 781.640 ;
        RECT 4.400 768.040 962.070 769.440 ;
        RECT 3.990 755.840 966.395 768.040 ;
        RECT 4.400 754.440 962.070 755.840 ;
        RECT 3.990 745.640 966.395 754.440 ;
        RECT 4.400 744.240 962.070 745.640 ;
        RECT 3.990 732.040 966.395 744.240 ;
        RECT 4.400 730.640 962.070 732.040 ;
        RECT 3.990 718.440 966.395 730.640 ;
        RECT 4.400 717.040 962.070 718.440 ;
        RECT 3.990 708.240 966.395 717.040 ;
        RECT 4.400 706.840 962.070 708.240 ;
        RECT 3.990 694.640 966.395 706.840 ;
        RECT 4.400 693.240 962.070 694.640 ;
        RECT 3.990 681.040 966.395 693.240 ;
        RECT 4.400 679.640 962.070 681.040 ;
        RECT 3.990 667.440 966.395 679.640 ;
        RECT 4.400 666.040 962.070 667.440 ;
        RECT 3.990 657.240 966.395 666.040 ;
        RECT 4.400 655.840 962.070 657.240 ;
        RECT 3.990 643.640 966.395 655.840 ;
        RECT 4.400 642.240 962.070 643.640 ;
        RECT 3.990 630.040 966.395 642.240 ;
        RECT 4.400 628.640 962.070 630.040 ;
        RECT 3.990 619.840 966.395 628.640 ;
        RECT 4.400 618.440 962.070 619.840 ;
        RECT 3.990 606.240 966.395 618.440 ;
        RECT 4.400 604.840 962.070 606.240 ;
        RECT 3.990 592.640 966.395 604.840 ;
        RECT 4.400 591.240 962.070 592.640 ;
        RECT 3.990 579.040 966.395 591.240 ;
        RECT 4.400 577.640 962.070 579.040 ;
        RECT 3.990 568.840 966.395 577.640 ;
        RECT 4.400 567.440 962.070 568.840 ;
        RECT 3.990 555.240 966.395 567.440 ;
        RECT 4.400 553.840 962.070 555.240 ;
        RECT 3.990 541.640 966.395 553.840 ;
        RECT 4.400 540.240 962.070 541.640 ;
        RECT 3.990 531.440 966.395 540.240 ;
        RECT 4.400 530.040 962.070 531.440 ;
        RECT 3.990 517.840 966.395 530.040 ;
        RECT 4.400 516.440 962.070 517.840 ;
        RECT 3.990 504.240 966.395 516.440 ;
        RECT 4.400 502.840 962.070 504.240 ;
        RECT 3.990 490.640 966.395 502.840 ;
        RECT 4.400 489.240 962.070 490.640 ;
        RECT 3.990 480.440 966.395 489.240 ;
        RECT 4.400 479.040 962.070 480.440 ;
        RECT 3.990 466.840 966.395 479.040 ;
        RECT 4.400 465.440 962.070 466.840 ;
        RECT 3.990 453.240 966.395 465.440 ;
        RECT 4.400 451.840 962.070 453.240 ;
        RECT 3.990 443.040 966.395 451.840 ;
        RECT 4.400 441.640 962.070 443.040 ;
        RECT 3.990 429.440 966.395 441.640 ;
        RECT 4.400 428.040 962.070 429.440 ;
        RECT 3.990 415.840 966.395 428.040 ;
        RECT 4.400 414.440 962.070 415.840 ;
        RECT 3.990 402.240 966.395 414.440 ;
        RECT 4.400 400.840 962.070 402.240 ;
        RECT 3.990 392.040 966.395 400.840 ;
        RECT 4.400 390.640 962.070 392.040 ;
        RECT 3.990 378.440 966.395 390.640 ;
        RECT 4.400 377.040 962.070 378.440 ;
        RECT 3.990 364.840 966.395 377.040 ;
        RECT 4.400 363.440 962.070 364.840 ;
        RECT 3.990 354.640 966.395 363.440 ;
        RECT 4.400 353.240 962.070 354.640 ;
        RECT 3.990 341.040 966.395 353.240 ;
        RECT 4.400 339.640 962.070 341.040 ;
        RECT 3.990 327.440 966.395 339.640 ;
        RECT 4.400 326.040 962.070 327.440 ;
        RECT 3.990 313.840 966.395 326.040 ;
        RECT 4.400 312.440 962.070 313.840 ;
        RECT 3.990 303.640 966.395 312.440 ;
        RECT 4.400 302.240 962.070 303.640 ;
        RECT 3.990 290.040 966.395 302.240 ;
        RECT 4.400 288.640 962.070 290.040 ;
        RECT 3.990 276.440 966.395 288.640 ;
        RECT 4.400 275.040 962.070 276.440 ;
        RECT 3.990 266.240 966.395 275.040 ;
        RECT 4.400 264.840 962.070 266.240 ;
        RECT 3.990 252.640 966.395 264.840 ;
        RECT 4.400 251.240 962.070 252.640 ;
        RECT 3.990 239.040 966.395 251.240 ;
        RECT 4.400 237.640 962.070 239.040 ;
        RECT 3.990 225.440 966.395 237.640 ;
        RECT 4.400 224.040 962.070 225.440 ;
        RECT 3.990 215.240 966.395 224.040 ;
        RECT 4.400 213.840 962.070 215.240 ;
        RECT 3.990 201.640 966.395 213.840 ;
        RECT 4.400 200.240 962.070 201.640 ;
        RECT 3.990 188.040 966.395 200.240 ;
        RECT 4.400 186.640 962.070 188.040 ;
        RECT 3.990 177.840 966.395 186.640 ;
        RECT 4.400 176.440 962.070 177.840 ;
        RECT 3.990 164.240 966.395 176.440 ;
        RECT 4.400 162.840 962.070 164.240 ;
        RECT 3.990 150.640 966.395 162.840 ;
        RECT 4.400 149.240 962.070 150.640 ;
        RECT 3.990 137.040 966.395 149.240 ;
        RECT 4.400 135.640 962.070 137.040 ;
        RECT 3.990 126.840 966.395 135.640 ;
        RECT 4.400 125.440 962.070 126.840 ;
        RECT 3.990 113.240 966.395 125.440 ;
        RECT 4.400 111.840 962.070 113.240 ;
        RECT 3.990 99.640 966.395 111.840 ;
        RECT 4.400 98.240 962.070 99.640 ;
        RECT 3.990 89.440 966.395 98.240 ;
        RECT 4.400 88.040 962.070 89.440 ;
        RECT 3.990 75.840 966.395 88.040 ;
        RECT 4.400 74.440 962.070 75.840 ;
        RECT 3.990 62.240 966.395 74.440 ;
        RECT 4.400 60.840 962.070 62.240 ;
        RECT 3.990 48.640 966.395 60.840 ;
        RECT 4.400 47.240 962.070 48.640 ;
        RECT 3.990 38.440 966.395 47.240 ;
        RECT 4.400 37.040 962.070 38.440 ;
        RECT 3.990 24.840 966.395 37.040 ;
        RECT 4.400 23.440 962.070 24.840 ;
        RECT 3.990 11.240 966.395 23.440 ;
        RECT 4.400 9.840 962.070 11.240 ;
        RECT 3.990 1.040 966.395 9.840 ;
        RECT 3.990 0.175 962.070 1.040 ;
      LAYER met4 ;
        RECT 10.415 15.135 20.640 964.065 ;
        RECT 23.040 15.135 97.440 964.065 ;
        RECT 99.840 15.135 174.240 964.065 ;
        RECT 176.640 15.135 251.040 964.065 ;
        RECT 253.440 15.135 327.840 964.065 ;
        RECT 330.240 15.135 404.640 964.065 ;
        RECT 407.040 15.135 481.440 964.065 ;
        RECT 483.840 15.135 558.240 964.065 ;
        RECT 560.640 15.135 635.040 964.065 ;
        RECT 637.440 15.135 711.840 964.065 ;
        RECT 714.240 15.135 788.640 964.065 ;
        RECT 791.040 15.135 865.440 964.065 ;
        RECT 867.840 15.135 942.240 964.065 ;
        RECT 944.640 15.135 962.945 964.065 ;
  END
END wrapped_silife
END LIBRARY

