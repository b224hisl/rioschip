VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO l1dcache
  CLASS BLOCK ;
  FOREIGN l1dcache ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 450.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END clk
  PIN data_chip_en_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END data_chip_en_1
  PIN data_chip_en_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END data_chip_en_2
  PIN data_in_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END data_in_1[0]
  PIN data_in_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 446.000 351.350 450.000 ;
    END
  END data_in_1[10]
  PIN data_in_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 446.000 203.230 450.000 ;
    END
  END data_in_1[11]
  PIN data_in_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 217.640 700.000 218.240 ;
    END
  END data_in_1[12]
  PIN data_in_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 446.000 348.130 450.000 ;
    END
  END data_in_1[13]
  PIN data_in_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 309.440 700.000 310.040 ;
    END
  END data_in_1[14]
  PIN data_in_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END data_in_1[15]
  PIN data_in_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 446.000 42.230 450.000 ;
    END
  END data_in_1[16]
  PIN data_in_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END data_in_1[17]
  PIN data_in_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 435.240 700.000 435.840 ;
    END
  END data_in_1[18]
  PIN data_in_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 176.840 700.000 177.440 ;
    END
  END data_in_1[19]
  PIN data_in_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END data_in_1[1]
  PIN data_in_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END data_in_1[20]
  PIN data_in_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END data_in_1[21]
  PIN data_in_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END data_in_1[22]
  PIN data_in_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 261.840 700.000 262.440 ;
    END
  END data_in_1[23]
  PIN data_in_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END data_in_1[24]
  PIN data_in_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END data_in_1[25]
  PIN data_in_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END data_in_1[26]
  PIN data_in_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END data_in_1[27]
  PIN data_in_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END data_in_1[28]
  PIN data_in_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 446.000 451.170 450.000 ;
    END
  END data_in_1[29]
  PIN data_in_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END data_in_1[2]
  PIN data_in_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 446.000 676.570 450.000 ;
    END
  END data_in_1[30]
  PIN data_in_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 446.000 528.450 450.000 ;
    END
  END data_in_1[31]
  PIN data_in_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 57.840 700.000 58.440 ;
    END
  END data_in_1[3]
  PIN data_in_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END data_in_1[4]
  PIN data_in_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 446.000 547.770 450.000 ;
    END
  END data_in_1[5]
  PIN data_in_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 446.000 389.990 450.000 ;
    END
  END data_in_1[6]
  PIN data_in_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 159.840 700.000 160.440 ;
    END
  END data_in_1[7]
  PIN data_in_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 446.000 55.110 450.000 ;
    END
  END data_in_1[8]
  PIN data_in_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END data_in_1[9]
  PIN data_in_2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 446.000 541.330 450.000 ;
    END
  END data_in_2[0]
  PIN data_in_2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 95.240 700.000 95.840 ;
    END
  END data_in_2[10]
  PIN data_in_2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 446.000 473.710 450.000 ;
    END
  END data_in_2[11]
  PIN data_in_2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 446.000 96.970 450.000 ;
    END
  END data_in_2[12]
  PIN data_in_2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END data_in_2[13]
  PIN data_in_2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 183.640 700.000 184.240 ;
    END
  END data_in_2[14]
  PIN data_in_2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END data_in_2[15]
  PIN data_in_2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 446.000 464.050 450.000 ;
    END
  END data_in_2[16]
  PIN data_in_2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END data_in_2[17]
  PIN data_in_2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END data_in_2[18]
  PIN data_in_2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END data_in_2[19]
  PIN data_in_2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 446.000 225.770 450.000 ;
    END
  END data_in_2[1]
  PIN data_in_2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 446.000 467.270 450.000 ;
    END
  END data_in_2[20]
  PIN data_in_2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 446.000 48.670 450.000 ;
    END
  END data_in_2[21]
  PIN data_in_2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 446.000 67.990 450.000 ;
    END
  END data_in_2[22]
  PIN data_in_2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 446.000 13.250 450.000 ;
    END
  END data_in_2[23]
  PIN data_in_2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END data_in_2[24]
  PIN data_in_2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END data_in_2[25]
  PIN data_in_2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END data_in_2[26]
  PIN data_in_2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 446.000 647.590 450.000 ;
    END
  END data_in_2[27]
  PIN data_in_2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END data_in_2[28]
  PIN data_in_2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 44.240 700.000 44.840 ;
    END
  END data_in_2[29]
  PIN data_in_2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END data_in_2[2]
  PIN data_in_2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END data_in_2[30]
  PIN data_in_2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 446.000 654.030 450.000 ;
    END
  END data_in_2[31]
  PIN data_in_2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 446.000 187.130 450.000 ;
    END
  END data_in_2[3]
  PIN data_in_2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END data_in_2[4]
  PIN data_in_2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 446.000 608.950 450.000 ;
    END
  END data_in_2[5]
  PIN data_in_2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END data_in_2[6]
  PIN data_in_2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 438.640 700.000 439.240 ;
    END
  END data_in_2[7]
  PIN data_in_2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END data_in_2[8]
  PIN data_in_2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END data_in_2[9]
  PIN data_index_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 289.040 700.000 289.640 ;
    END
  END data_index_1[0]
  PIN data_index_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END data_index_1[1]
  PIN data_index_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END data_index_1[2]
  PIN data_index_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 136.040 700.000 136.640 ;
    END
  END data_index_1[3]
  PIN data_index_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 446.000 309.490 450.000 ;
    END
  END data_index_1[4]
  PIN data_index_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END data_index_1[5]
  PIN data_index_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END data_index_1[6]
  PIN data_index_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 446.000 241.870 450.000 ;
    END
  END data_index_1[7]
  PIN data_index_2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END data_index_2[0]
  PIN data_index_2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 446.000 550.990 450.000 ;
    END
  END data_index_2[1]
  PIN data_index_2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 408.040 700.000 408.640 ;
    END
  END data_index_2[2]
  PIN data_index_2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 374.040 700.000 374.640 ;
    END
  END data_index_2[3]
  PIN data_index_2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END data_index_2[4]
  PIN data_index_2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END data_index_2[5]
  PIN data_index_2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END data_index_2[6]
  PIN data_index_2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END data_index_2[7]
  PIN data_out_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 295.840 700.000 296.440 ;
    END
  END data_out_1[0]
  PIN data_out_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END data_out_1[10]
  PIN data_out_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 163.240 700.000 163.840 ;
    END
  END data_out_1[11]
  PIN data_out_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 446.000 499.470 450.000 ;
    END
  END data_out_1[12]
  PIN data_out_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 370.640 700.000 371.240 ;
    END
  END data_out_1[13]
  PIN data_out_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 122.440 700.000 123.040 ;
    END
  END data_out_1[14]
  PIN data_out_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END data_out_1[15]
  PIN data_out_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 170.040 700.000 170.640 ;
    END
  END data_out_1[16]
  PIN data_out_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END data_out_1[17]
  PIN data_out_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 23.840 700.000 24.440 ;
    END
  END data_out_1[18]
  PIN data_out_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END data_out_1[19]
  PIN data_out_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END data_out_1[1]
  PIN data_out_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 446.000 525.230 450.000 ;
    END
  END data_out_1[20]
  PIN data_out_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 446.000 161.370 450.000 ;
    END
  END data_out_1[21]
  PIN data_out_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 446.000 216.110 450.000 ;
    END
  END data_out_1[22]
  PIN data_out_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END data_out_1[23]
  PIN data_out_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 190.440 700.000 191.040 ;
    END
  END data_out_1[24]
  PIN data_out_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END data_out_1[25]
  PIN data_out_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END data_out_1[26]
  PIN data_out_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 446.000 409.310 450.000 ;
    END
  END data_out_1[27]
  PIN data_out_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 37.440 700.000 38.040 ;
    END
  END data_out_1[28]
  PIN data_out_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 446.000 663.690 450.000 ;
    END
  END data_out_1[29]
  PIN data_out_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END data_out_1[2]
  PIN data_out_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 329.840 700.000 330.440 ;
    END
  END data_out_1[30]
  PIN data_out_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END data_out_1[31]
  PIN data_out_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 282.240 700.000 282.840 ;
    END
  END data_out_1[3]
  PIN data_out_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 446.000 354.570 450.000 ;
    END
  END data_out_1[4]
  PIN data_out_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END data_out_1[5]
  PIN data_out_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END data_out_1[6]
  PIN data_out_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END data_out_1[7]
  PIN data_out_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END data_out_1[8]
  PIN data_out_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END data_out_1[9]
  PIN data_out_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END data_out_2[0]
  PIN data_out_2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 446.000 341.690 450.000 ;
    END
  END data_out_2[10]
  PIN data_out_2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 387.640 700.000 388.240 ;
    END
  END data_out_2[11]
  PIN data_out_2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 446.000 441.510 450.000 ;
    END
  END data_out_2[12]
  PIN data_out_2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END data_out_2[13]
  PIN data_out_2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 446.000 248.310 450.000 ;
    END
  END data_out_2[14]
  PIN data_out_2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END data_out_2[15]
  PIN data_out_2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 446.000 489.810 450.000 ;
    END
  END data_out_2[16]
  PIN data_out_2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END data_out_2[17]
  PIN data_out_2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 446.000 174.250 450.000 ;
    END
  END data_out_2[18]
  PIN data_out_2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END data_out_2[19]
  PIN data_out_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END data_out_2[1]
  PIN data_out_2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 91.840 700.000 92.440 ;
    END
  END data_out_2[20]
  PIN data_out_2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END data_out_2[21]
  PIN data_out_2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 446.000 612.170 450.000 ;
    END
  END data_out_2[22]
  PIN data_out_2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 446.000 576.750 450.000 ;
    END
  END data_out_2[23]
  PIN data_out_2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 446.000 422.190 450.000 ;
    END
  END data_out_2[24]
  PIN data_out_2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END data_out_2[25]
  PIN data_out_2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END data_out_2[26]
  PIN data_out_2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 446.000 26.130 450.000 ;
    END
  END data_out_2[27]
  PIN data_out_2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END data_out_2[28]
  PIN data_out_2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END data_out_2[29]
  PIN data_out_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 446.000 154.930 450.000 ;
    END
  END data_out_2[2]
  PIN data_out_2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 156.440 700.000 157.040 ;
    END
  END data_out_2[30]
  PIN data_out_2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 446.000 29.350 450.000 ;
    END
  END data_out_2[31]
  PIN data_out_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 446.000 113.070 450.000 ;
    END
  END data_out_2[3]
  PIN data_out_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END data_out_2[4]
  PIN data_out_2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 446.000 454.390 450.000 ;
    END
  END data_out_2[5]
  PIN data_out_2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END data_out_2[6]
  PIN data_out_2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 446.000 325.590 450.000 ;
    END
  END data_out_2[7]
  PIN data_out_2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 446.000 51.890 450.000 ;
    END
  END data_out_2[8]
  PIN data_out_2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END data_out_2[9]
  PIN data_write_en_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END data_write_en_1
  PIN data_write_en_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END data_write_en_2
  PIN ld_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END ld_data_o[0]
  PIN ld_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 380.840 700.000 381.440 ;
    END
  END ld_data_o[10]
  PIN ld_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 108.840 700.000 109.440 ;
    END
  END ld_data_o[11]
  PIN ld_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END ld_data_o[12]
  PIN ld_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 446.000 142.050 450.000 ;
    END
  END ld_data_o[13]
  PIN ld_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END ld_data_o[14]
  PIN ld_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END ld_data_o[15]
  PIN ld_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END ld_data_o[16]
  PIN ld_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 446.000 290.170 450.000 ;
    END
  END ld_data_o[17]
  PIN ld_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 446.000 77.650 450.000 ;
    END
  END ld_data_o[18]
  PIN ld_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 446.000 74.430 450.000 ;
    END
  END ld_data_o[19]
  PIN ld_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 397.840 700.000 398.440 ;
    END
  END ld_data_o[1]
  PIN ld_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 446.000 303.050 450.000 ;
    END
  END ld_data_o[20]
  PIN ld_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 446.000 296.610 450.000 ;
    END
  END ld_data_o[21]
  PIN ld_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END ld_data_o[22]
  PIN ld_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END ld_data_o[23]
  PIN ld_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 446.000 264.410 450.000 ;
    END
  END ld_data_o[24]
  PIN ld_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 446.000 438.290 450.000 ;
    END
  END ld_data_o[25]
  PIN ld_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 446.000 579.970 450.000 ;
    END
  END ld_data_o[26]
  PIN ld_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END ld_data_o[27]
  PIN ld_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 129.240 700.000 129.840 ;
    END
  END ld_data_o[28]
  PIN ld_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END ld_data_o[29]
  PIN ld_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 204.040 700.000 204.640 ;
    END
  END ld_data_o[2]
  PIN ld_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END ld_data_o[30]
  PIN ld_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 446.000 380.330 450.000 ;
    END
  END ld_data_o[31]
  PIN ld_data_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 78.240 700.000 78.840 ;
    END
  END ld_data_o[32]
  PIN ld_data_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 446.000 428.630 450.000 ;
    END
  END ld_data_o[33]
  PIN ld_data_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END ld_data_o[34]
  PIN ld_data_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 442.040 700.000 442.640 ;
    END
  END ld_data_o[35]
  PIN ld_data_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 446.000 200.010 450.000 ;
    END
  END ld_data_o[36]
  PIN ld_data_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END ld_data_o[37]
  PIN ld_data_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END ld_data_o[38]
  PIN ld_data_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 353.640 700.000 354.240 ;
    END
  END ld_data_o[39]
  PIN ld_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 448.840 700.000 449.440 ;
    END
  END ld_data_o[3]
  PIN ld_data_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END ld_data_o[40]
  PIN ld_data_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 446.000 277.290 450.000 ;
    END
  END ld_data_o[41]
  PIN ld_data_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 394.440 700.000 395.040 ;
    END
  END ld_data_o[42]
  PIN ld_data_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 446.000 412.530 450.000 ;
    END
  END ld_data_o[43]
  PIN ld_data_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 231.240 700.000 231.840 ;
    END
  END ld_data_o[44]
  PIN ld_data_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END ld_data_o[45]
  PIN ld_data_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 446.000 164.590 450.000 ;
    END
  END ld_data_o[46]
  PIN ld_data_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END ld_data_o[47]
  PIN ld_data_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END ld_data_o[48]
  PIN ld_data_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END ld_data_o[49]
  PIN ld_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END ld_data_o[4]
  PIN ld_data_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END ld_data_o[50]
  PIN ld_data_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 446.000 386.770 450.000 ;
    END
  END ld_data_o[51]
  PIN ld_data_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 446.000 138.830 450.000 ;
    END
  END ld_data_o[52]
  PIN ld_data_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END ld_data_o[53]
  PIN ld_data_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END ld_data_o[54]
  PIN ld_data_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 446.000 673.350 450.000 ;
    END
  END ld_data_o[55]
  PIN ld_data_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END ld_data_o[56]
  PIN ld_data_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 0.040 700.000 0.640 ;
    END
  END ld_data_o[57]
  PIN ld_data_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END ld_data_o[58]
  PIN ld_data_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END ld_data_o[59]
  PIN ld_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 446.000 100.190 450.000 ;
    END
  END ld_data_o[5]
  PIN ld_data_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 446.000 328.810 450.000 ;
    END
  END ld_data_o[60]
  PIN ld_data_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END ld_data_o[61]
  PIN ld_data_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END ld_data_o[62]
  PIN ld_data_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 446.000 122.730 450.000 ;
    END
  END ld_data_o[63]
  PIN ld_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END ld_data_o[6]
  PIN ld_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END ld_data_o[7]
  PIN ld_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 446.000 377.110 450.000 ;
    END
  END ld_data_o[8]
  PIN ld_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END ld_data_o[9]
  PIN opcode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 446.000 335.250 450.000 ;
    END
  END opcode
  PIN req_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END req_addr_i[0]
  PIN req_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END req_addr_i[10]
  PIN req_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END req_addr_i[11]
  PIN req_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END req_addr_i[12]
  PIN req_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END req_addr_i[13]
  PIN req_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END req_addr_i[14]
  PIN req_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 173.440 700.000 174.040 ;
    END
  END req_addr_i[15]
  PIN req_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END req_addr_i[16]
  PIN req_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END req_addr_i[17]
  PIN req_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END req_addr_i[18]
  PIN req_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END req_addr_i[19]
  PIN req_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END req_addr_i[1]
  PIN req_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 446.000 312.710 450.000 ;
    END
  END req_addr_i[20]
  PIN req_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 446.000 238.650 450.000 ;
    END
  END req_addr_i[21]
  PIN req_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 446.000 699.110 450.000 ;
    END
  END req_addr_i[22]
  PIN req_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 446.000 364.230 450.000 ;
    END
  END req_addr_i[23]
  PIN req_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 446.000 16.470 450.000 ;
    END
  END req_addr_i[24]
  PIN req_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END req_addr_i[25]
  PIN req_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END req_addr_i[26]
  PIN req_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 446.000 621.830 450.000 ;
    END
  END req_addr_i[27]
  PIN req_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END req_addr_i[28]
  PIN req_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END req_addr_i[29]
  PIN req_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END req_addr_i[2]
  PIN req_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 13.640 700.000 14.240 ;
    END
  END req_addr_i[30]
  PIN req_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END req_addr_i[31]
  PIN req_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END req_addr_i[3]
  PIN req_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 446.000 338.470 450.000 ;
    END
  END req_addr_i[4]
  PIN req_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END req_addr_i[5]
  PIN req_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 446.000 254.750 450.000 ;
    END
  END req_addr_i[6]
  PIN req_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END req_addr_i[7]
  PIN req_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END req_addr_i[8]
  PIN req_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 446.000 628.270 450.000 ;
    END
  END req_addr_i[9]
  PIN req_ready_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END req_ready_o
  PIN req_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END req_valid_i
  PIN resp_ready_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END resp_ready_i
  PIN resp_valid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 446.000 80.870 450.000 ;
    END
  END resp_valid_o
  PIN rob_index_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 446.000 679.790 450.000 ;
    END
  END rob_index_i
  PIN rob_index_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 446.000 261.190 450.000 ;
    END
  END rob_index_o
  PIN rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 446.000 125.950 450.000 ;
    END
  END rstn
  PIN st_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 446.000 650.810 450.000 ;
    END
  END st_data_i[0]
  PIN st_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 446.000 560.650 450.000 ;
    END
  END st_data_i[10]
  PIN st_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END st_data_i[11]
  PIN st_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 446.000 641.150 450.000 ;
    END
  END st_data_i[12]
  PIN st_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END st_data_i[13]
  PIN st_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END st_data_i[14]
  PIN st_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END st_data_i[15]
  PIN st_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 446.000 103.410 450.000 ;
    END
  END st_data_i[16]
  PIN st_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END st_data_i[17]
  PIN st_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END st_data_i[18]
  PIN st_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 446.000 267.630 450.000 ;
    END
  END st_data_i[19]
  PIN st_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END st_data_i[1]
  PIN st_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END st_data_i[20]
  PIN st_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 306.040 700.000 306.640 ;
    END
  END st_data_i[21]
  PIN st_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END st_data_i[22]
  PIN st_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 265.240 700.000 265.840 ;
    END
  END st_data_i[23]
  PIN st_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END st_data_i[24]
  PIN st_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END st_data_i[25]
  PIN st_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 64.640 700.000 65.240 ;
    END
  END st_data_i[26]
  PIN st_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 446.000 586.410 450.000 ;
    END
  END st_data_i[27]
  PIN st_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 446.000 212.890 450.000 ;
    END
  END st_data_i[28]
  PIN st_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 446.000 567.090 450.000 ;
    END
  END st_data_i[29]
  PIN st_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 446.000 625.050 450.000 ;
    END
  END st_data_i[2]
  PIN st_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END st_data_i[30]
  PIN st_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 446.000 460.830 450.000 ;
    END
  END st_data_i[31]
  PIN st_data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 446.000 602.510 450.000 ;
    END
  END st_data_i[32]
  PIN st_data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 446.000 435.070 450.000 ;
    END
  END st_data_i[33]
  PIN st_data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 292.440 700.000 293.040 ;
    END
  END st_data_i[34]
  PIN st_data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END st_data_i[35]
  PIN st_data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END st_data_i[36]
  PIN st_data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 401.240 700.000 401.840 ;
    END
  END st_data_i[37]
  PIN st_data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 446.000 322.370 450.000 ;
    END
  END st_data_i[38]
  PIN st_data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END st_data_i[39]
  PIN st_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END st_data_i[3]
  PIN st_data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 446.000 209.670 450.000 ;
    END
  END st_data_i[40]
  PIN st_data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END st_data_i[41]
  PIN st_data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END st_data_i[42]
  PIN st_data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 414.840 700.000 415.440 ;
    END
  END st_data_i[43]
  PIN st_data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END st_data_i[44]
  PIN st_data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 105.440 700.000 106.040 ;
    END
  END st_data_i[45]
  PIN st_data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END st_data_i[46]
  PIN st_data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 346.840 700.000 347.440 ;
    END
  END st_data_i[47]
  PIN st_data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 98.640 700.000 99.240 ;
    END
  END st_data_i[48]
  PIN st_data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 446.000 634.710 450.000 ;
    END
  END st_data_i[49]
  PIN st_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 446.000 692.670 450.000 ;
    END
  END st_data_i[4]
  PIN st_data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END st_data_i[50]
  PIN st_data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 210.840 700.000 211.440 ;
    END
  END st_data_i[51]
  PIN st_data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END st_data_i[52]
  PIN st_data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 81.640 700.000 82.240 ;
    END
  END st_data_i[53]
  PIN st_data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END st_data_i[54]
  PIN st_data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 446.000 447.950 450.000 ;
    END
  END st_data_i[55]
  PIN st_data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END st_data_i[56]
  PIN st_data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END st_data_i[57]
  PIN st_data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 316.240 700.000 316.840 ;
    END
  END st_data_i[58]
  PIN st_data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 17.040 700.000 17.640 ;
    END
  END st_data_i[59]
  PIN st_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END st_data_i[5]
  PIN st_data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 446.000 22.910 450.000 ;
    END
  END st_data_i[60]
  PIN st_data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END st_data_i[61]
  PIN st_data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END st_data_i[62]
  PIN st_data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 446.000 235.430 450.000 ;
    END
  END st_data_i[63]
  PIN st_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 255.040 700.000 255.640 ;
    END
  END st_data_i[6]
  PIN st_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 446.000 280.510 450.000 ;
    END
  END st_data_i[7]
  PIN st_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 68.040 700.000 68.640 ;
    END
  END st_data_i[8]
  PIN st_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END st_data_i[9]
  PIN tag_chip_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END tag_chip_en
  PIN tag_data_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 187.040 700.000 187.640 ;
    END
  END tag_data_in[0]
  PIN tag_data_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 446.000 367.450 450.000 ;
    END
  END tag_data_in[10]
  PIN tag_data_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END tag_data_in[11]
  PIN tag_data_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END tag_data_in[12]
  PIN tag_data_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END tag_data_in[13]
  PIN tag_data_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END tag_data_in[14]
  PIN tag_data_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END tag_data_in[15]
  PIN tag_data_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 446.000 10.030 450.000 ;
    END
  END tag_data_in[16]
  PIN tag_data_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END tag_data_in[17]
  PIN tag_data_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 446.000 315.930 450.000 ;
    END
  END tag_data_in[18]
  PIN tag_data_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 40.840 700.000 41.440 ;
    END
  END tag_data_in[19]
  PIN tag_data_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 446.000 3.590 450.000 ;
    END
  END tag_data_in[1]
  PIN tag_data_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 3.440 700.000 4.040 ;
    END
  END tag_data_in[20]
  PIN tag_data_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END tag_data_in[21]
  PIN tag_data_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 446.000 373.890 450.000 ;
    END
  END tag_data_in[22]
  PIN tag_data_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 446.000 0.370 450.000 ;
    END
  END tag_data_in[23]
  PIN tag_data_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 119.040 700.000 119.640 ;
    END
  END tag_data_in[24]
  PIN tag_data_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 367.240 700.000 367.840 ;
    END
  END tag_data_in[25]
  PIN tag_data_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 428.440 700.000 429.040 ;
    END
  END tag_data_in[26]
  PIN tag_data_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 446.000 589.630 450.000 ;
    END
  END tag_data_in[27]
  PIN tag_data_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 360.440 700.000 361.040 ;
    END
  END tag_data_in[28]
  PIN tag_data_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 446.000 399.650 450.000 ;
    END
  END tag_data_in[29]
  PIN tag_data_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END tag_data_in[2]
  PIN tag_data_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END tag_data_in[30]
  PIN tag_data_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 446.000 177.470 450.000 ;
    END
  END tag_data_in[31]
  PIN tag_data_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 142.840 700.000 143.440 ;
    END
  END tag_data_in[3]
  PIN tag_data_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END tag_data_in[4]
  PIN tag_data_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END tag_data_in[5]
  PIN tag_data_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 268.640 700.000 269.240 ;
    END
  END tag_data_in[6]
  PIN tag_data_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 197.240 700.000 197.840 ;
    END
  END tag_data_in[7]
  PIN tag_data_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END tag_data_in[8]
  PIN tag_data_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END tag_data_in[9]
  PIN tag_index[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 446.000 151.710 450.000 ;
    END
  END tag_index[0]
  PIN tag_index[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 333.240 700.000 333.840 ;
    END
  END tag_index[1]
  PIN tag_index[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END tag_index[2]
  PIN tag_index[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END tag_index[3]
  PIN tag_index[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END tag_index[4]
  PIN tag_index[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END tag_index[5]
  PIN tag_index[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END tag_index[6]
  PIN tag_index[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END tag_index[7]
  PIN tag_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 278.840 700.000 279.440 ;
    END
  END tag_out[0]
  PIN tag_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END tag_out[10]
  PIN tag_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 446.000 480.150 450.000 ;
    END
  END tag_out[11]
  PIN tag_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 446.000 396.430 450.000 ;
    END
  END tag_out[12]
  PIN tag_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END tag_out[13]
  PIN tag_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 336.640 700.000 337.240 ;
    END
  END tag_out[14]
  PIN tag_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END tag_out[15]
  PIN tag_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 446.000 90.530 450.000 ;
    END
  END tag_out[16]
  PIN tag_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END tag_out[17]
  PIN tag_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END tag_out[18]
  PIN tag_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 446.000 599.290 450.000 ;
    END
  END tag_out[19]
  PIN tag_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 446.000 563.870 450.000 ;
    END
  END tag_out[1]
  PIN tag_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 446.000 660.470 450.000 ;
    END
  END tag_out[20]
  PIN tag_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 446.000 686.230 450.000 ;
    END
  END tag_out[21]
  PIN tag_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 446.000 689.450 450.000 ;
    END
  END tag_out[22]
  PIN tag_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END tag_out[23]
  PIN tag_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 446.000 509.130 450.000 ;
    END
  END tag_out[24]
  PIN tag_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END tag_out[25]
  PIN tag_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END tag_out[26]
  PIN tag_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 446.000 129.170 450.000 ;
    END
  END tag_out[27]
  PIN tag_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END tag_out[28]
  PIN tag_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END tag_out[29]
  PIN tag_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END tag_out[2]
  PIN tag_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END tag_out[30]
  PIN tag_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 446.000 196.790 450.000 ;
    END
  END tag_out[31]
  PIN tag_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END tag_out[3]
  PIN tag_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END tag_out[4]
  PIN tag_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END tag_out[5]
  PIN tag_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 446.000 486.590 450.000 ;
    END
  END tag_out[6]
  PIN tag_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END tag_out[7]
  PIN tag_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END tag_out[8]
  PIN tag_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END tag_out[9]
  PIN tag_write_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 227.840 700.000 228.440 ;
    END
  END tag_write_en
  PIN type_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 343.440 700.000 344.040 ;
    END
  END type_i[0]
  PIN type_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END type_i[1]
  PIN type_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 446.000 180.690 450.000 ;
    END
  END type_i[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 438.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 438.160 ;
    END
  END vssd1
  PIN wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END wb_ack_i
  PIN wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 446.000 64.770 450.000 ;
    END
  END wb_adr_o[0]
  PIN wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 446.000 402.870 450.000 ;
    END
  END wb_adr_o[10]
  PIN wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 238.040 700.000 238.640 ;
    END
  END wb_adr_o[11]
  PIN wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END wb_adr_o[12]
  PIN wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END wb_adr_o[13]
  PIN wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END wb_adr_o[14]
  PIN wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 446.000 361.010 450.000 ;
    END
  END wb_adr_o[15]
  PIN wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END wb_adr_o[16]
  PIN wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 446.000 148.490 450.000 ;
    END
  END wb_adr_o[17]
  PIN wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wb_adr_o[18]
  PIN wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 224.440 700.000 225.040 ;
    END
  END wb_adr_o[19]
  PIN wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wb_adr_o[1]
  PIN wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END wb_adr_o[20]
  PIN wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wb_adr_o[21]
  PIN wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END wb_adr_o[22]
  PIN wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wb_adr_o[23]
  PIN wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 446.000 534.890 450.000 ;
    END
  END wb_adr_o[24]
  PIN wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 384.240 700.000 384.840 ;
    END
  END wb_adr_o[25]
  PIN wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 446.000 167.810 450.000 ;
    END
  END wb_adr_o[26]
  PIN wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 446.000 222.550 450.000 ;
    END
  END wb_adr_o[27]
  PIN wb_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 6.840 700.000 7.440 ;
    END
  END wb_adr_o[28]
  PIN wb_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 446.000 135.610 450.000 ;
    END
  END wb_adr_o[29]
  PIN wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 112.240 700.000 112.840 ;
    END
  END wb_adr_o[2]
  PIN wb_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END wb_adr_o[30]
  PIN wb_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 446.000 299.830 450.000 ;
    END
  END wb_adr_o[31]
  PIN wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 446.000 61.550 450.000 ;
    END
  END wb_adr_o[3]
  PIN wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wb_adr_o[4]
  PIN wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END wb_adr_o[5]
  PIN wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END wb_adr_o[6]
  PIN wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 319.640 700.000 320.240 ;
    END
  END wb_adr_o[7]
  PIN wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END wb_adr_o[8]
  PIN wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 275.440 700.000 276.040 ;
    END
  END wb_adr_o[9]
  PIN wb_bl_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 85.040 700.000 85.640 ;
    END
  END wb_bl_o[0]
  PIN wb_bl_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END wb_bl_o[1]
  PIN wb_bl_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 446.000 425.410 450.000 ;
    END
  END wb_bl_o[2]
  PIN wb_bl_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 446.000 592.850 450.000 ;
    END
  END wb_bl_o[3]
  PIN wb_bl_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wb_bl_o[4]
  PIN wb_bl_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END wb_bl_o[5]
  PIN wb_bl_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 30.640 700.000 31.240 ;
    END
  END wb_bl_o[6]
  PIN wb_bl_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 446.000 116.290 450.000 ;
    END
  END wb_bl_o[7]
  PIN wb_bl_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wb_bl_o[8]
  PIN wb_bl_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wb_bl_o[9]
  PIN wb_bry_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END wb_bry_o
  PIN wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 251.640 700.000 252.240 ;
    END
  END wb_cyc_o
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 446.000 666.910 450.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 146.240 700.000 146.840 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 446.000 512.350 450.000 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 51.040 700.000 51.640 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 446.000 251.530 450.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 421.640 700.000 422.240 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 200.640 700.000 201.240 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 446.000 476.930 450.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 446.000 615.390 450.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 446.000 109.850 450.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 248.240 700.000 248.840 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 446.000 637.930 450.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 357.040 700.000 357.640 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 71.440 700.000 72.040 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 446.000 573.530 450.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 446.000 228.990 450.000 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 241.440 700.000 242.040 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 54.440 700.000 55.040 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 132.640 700.000 133.240 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 446.000 554.210 450.000 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 411.440 700.000 412.040 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 214.240 700.000 214.840 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 425.040 700.000 425.640 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 446.000 538.110 450.000 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 446.000 522.010 450.000 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 446.000 39.010 450.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 446.000 274.070 450.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 446.000 415.750 450.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 446.000 286.950 450.000 ;
    END
  END wb_dat_o[9]
  PIN wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END wb_sel_o[0]
  PIN wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 446.000 515.570 450.000 ;
    END
  END wb_sel_o[1]
  PIN wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 27.240 700.000 27.840 ;
    END
  END wb_sel_o[2]
  PIN wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END wb_sel_o[3]
  PIN wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 323.040 700.000 323.640 ;
    END
  END wb_stb_o
  PIN wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wb_we_o
  PIN write_data_mask_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END write_data_mask_1[0]
  PIN write_data_mask_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END write_data_mask_1[1]
  PIN write_data_mask_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 302.640 700.000 303.240 ;
    END
  END write_data_mask_1[2]
  PIN write_data_mask_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END write_data_mask_1[3]
  PIN write_data_mask_2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 446.000 502.690 450.000 ;
    END
  END write_data_mask_2[0]
  PIN write_data_mask_2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 446.000 493.030 450.000 ;
    END
  END write_data_mask_2[1]
  PIN write_data_mask_2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 446.000 87.310 450.000 ;
    END
  END write_data_mask_2[2]
  PIN write_data_mask_2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 446.000 190.350 450.000 ;
    END
  END write_data_mask_2[3]
  PIN write_tag_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END write_tag_mask[0]
  PIN write_tag_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END write_tag_mask[1]
  PIN write_tag_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 446.000 35.790 450.000 ;
    END
  END write_tag_mask[2]
  PIN write_tag_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 149.640 700.000 150.240 ;
    END
  END write_tag_mask[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 694.140 438.005 ;
      LAYER met1 ;
        RECT 0.070 6.160 699.130 441.280 ;
      LAYER met2 ;
        RECT 0.650 445.720 3.030 449.325 ;
        RECT 3.870 445.720 9.470 449.325 ;
        RECT 10.310 445.720 12.690 449.325 ;
        RECT 13.530 445.720 15.910 449.325 ;
        RECT 16.750 445.720 22.350 449.325 ;
        RECT 23.190 445.720 25.570 449.325 ;
        RECT 26.410 445.720 28.790 449.325 ;
        RECT 29.630 445.720 35.230 449.325 ;
        RECT 36.070 445.720 38.450 449.325 ;
        RECT 39.290 445.720 41.670 449.325 ;
        RECT 42.510 445.720 48.110 449.325 ;
        RECT 48.950 445.720 51.330 449.325 ;
        RECT 52.170 445.720 54.550 449.325 ;
        RECT 55.390 445.720 60.990 449.325 ;
        RECT 61.830 445.720 64.210 449.325 ;
        RECT 65.050 445.720 67.430 449.325 ;
        RECT 68.270 445.720 73.870 449.325 ;
        RECT 74.710 445.720 77.090 449.325 ;
        RECT 77.930 445.720 80.310 449.325 ;
        RECT 81.150 445.720 86.750 449.325 ;
        RECT 87.590 445.720 89.970 449.325 ;
        RECT 90.810 445.720 96.410 449.325 ;
        RECT 97.250 445.720 99.630 449.325 ;
        RECT 100.470 445.720 102.850 449.325 ;
        RECT 103.690 445.720 109.290 449.325 ;
        RECT 110.130 445.720 112.510 449.325 ;
        RECT 113.350 445.720 115.730 449.325 ;
        RECT 116.570 445.720 122.170 449.325 ;
        RECT 123.010 445.720 125.390 449.325 ;
        RECT 126.230 445.720 128.610 449.325 ;
        RECT 129.450 445.720 135.050 449.325 ;
        RECT 135.890 445.720 138.270 449.325 ;
        RECT 139.110 445.720 141.490 449.325 ;
        RECT 142.330 445.720 147.930 449.325 ;
        RECT 148.770 445.720 151.150 449.325 ;
        RECT 151.990 445.720 154.370 449.325 ;
        RECT 155.210 445.720 160.810 449.325 ;
        RECT 161.650 445.720 164.030 449.325 ;
        RECT 164.870 445.720 167.250 449.325 ;
        RECT 168.090 445.720 173.690 449.325 ;
        RECT 174.530 445.720 176.910 449.325 ;
        RECT 177.750 445.720 180.130 449.325 ;
        RECT 180.970 445.720 186.570 449.325 ;
        RECT 187.410 445.720 189.790 449.325 ;
        RECT 190.630 445.720 196.230 449.325 ;
        RECT 197.070 445.720 199.450 449.325 ;
        RECT 200.290 445.720 202.670 449.325 ;
        RECT 203.510 445.720 209.110 449.325 ;
        RECT 209.950 445.720 212.330 449.325 ;
        RECT 213.170 445.720 215.550 449.325 ;
        RECT 216.390 445.720 221.990 449.325 ;
        RECT 222.830 445.720 225.210 449.325 ;
        RECT 226.050 445.720 228.430 449.325 ;
        RECT 229.270 445.720 234.870 449.325 ;
        RECT 235.710 445.720 238.090 449.325 ;
        RECT 238.930 445.720 241.310 449.325 ;
        RECT 242.150 445.720 247.750 449.325 ;
        RECT 248.590 445.720 250.970 449.325 ;
        RECT 251.810 445.720 254.190 449.325 ;
        RECT 255.030 445.720 260.630 449.325 ;
        RECT 261.470 445.720 263.850 449.325 ;
        RECT 264.690 445.720 267.070 449.325 ;
        RECT 267.910 445.720 273.510 449.325 ;
        RECT 274.350 445.720 276.730 449.325 ;
        RECT 277.570 445.720 279.950 449.325 ;
        RECT 280.790 445.720 286.390 449.325 ;
        RECT 287.230 445.720 289.610 449.325 ;
        RECT 290.450 445.720 296.050 449.325 ;
        RECT 296.890 445.720 299.270 449.325 ;
        RECT 300.110 445.720 302.490 449.325 ;
        RECT 303.330 445.720 308.930 449.325 ;
        RECT 309.770 445.720 312.150 449.325 ;
        RECT 312.990 445.720 315.370 449.325 ;
        RECT 316.210 445.720 321.810 449.325 ;
        RECT 322.650 445.720 325.030 449.325 ;
        RECT 325.870 445.720 328.250 449.325 ;
        RECT 329.090 445.720 334.690 449.325 ;
        RECT 335.530 445.720 337.910 449.325 ;
        RECT 338.750 445.720 341.130 449.325 ;
        RECT 341.970 445.720 347.570 449.325 ;
        RECT 348.410 445.720 350.790 449.325 ;
        RECT 351.630 445.720 354.010 449.325 ;
        RECT 354.850 445.720 360.450 449.325 ;
        RECT 361.290 445.720 363.670 449.325 ;
        RECT 364.510 445.720 366.890 449.325 ;
        RECT 367.730 445.720 373.330 449.325 ;
        RECT 374.170 445.720 376.550 449.325 ;
        RECT 377.390 445.720 379.770 449.325 ;
        RECT 380.610 445.720 386.210 449.325 ;
        RECT 387.050 445.720 389.430 449.325 ;
        RECT 390.270 445.720 395.870 449.325 ;
        RECT 396.710 445.720 399.090 449.325 ;
        RECT 399.930 445.720 402.310 449.325 ;
        RECT 403.150 445.720 408.750 449.325 ;
        RECT 409.590 445.720 411.970 449.325 ;
        RECT 412.810 445.720 415.190 449.325 ;
        RECT 416.030 445.720 421.630 449.325 ;
        RECT 422.470 445.720 424.850 449.325 ;
        RECT 425.690 445.720 428.070 449.325 ;
        RECT 428.910 445.720 434.510 449.325 ;
        RECT 435.350 445.720 437.730 449.325 ;
        RECT 438.570 445.720 440.950 449.325 ;
        RECT 441.790 445.720 447.390 449.325 ;
        RECT 448.230 445.720 450.610 449.325 ;
        RECT 451.450 445.720 453.830 449.325 ;
        RECT 454.670 445.720 460.270 449.325 ;
        RECT 461.110 445.720 463.490 449.325 ;
        RECT 464.330 445.720 466.710 449.325 ;
        RECT 467.550 445.720 473.150 449.325 ;
        RECT 473.990 445.720 476.370 449.325 ;
        RECT 477.210 445.720 479.590 449.325 ;
        RECT 480.430 445.720 486.030 449.325 ;
        RECT 486.870 445.720 489.250 449.325 ;
        RECT 490.090 445.720 492.470 449.325 ;
        RECT 493.310 445.720 498.910 449.325 ;
        RECT 499.750 445.720 502.130 449.325 ;
        RECT 502.970 445.720 508.570 449.325 ;
        RECT 509.410 445.720 511.790 449.325 ;
        RECT 512.630 445.720 515.010 449.325 ;
        RECT 515.850 445.720 521.450 449.325 ;
        RECT 522.290 445.720 524.670 449.325 ;
        RECT 525.510 445.720 527.890 449.325 ;
        RECT 528.730 445.720 534.330 449.325 ;
        RECT 535.170 445.720 537.550 449.325 ;
        RECT 538.390 445.720 540.770 449.325 ;
        RECT 541.610 445.720 547.210 449.325 ;
        RECT 548.050 445.720 550.430 449.325 ;
        RECT 551.270 445.720 553.650 449.325 ;
        RECT 554.490 445.720 560.090 449.325 ;
        RECT 560.930 445.720 563.310 449.325 ;
        RECT 564.150 445.720 566.530 449.325 ;
        RECT 567.370 445.720 572.970 449.325 ;
        RECT 573.810 445.720 576.190 449.325 ;
        RECT 577.030 445.720 579.410 449.325 ;
        RECT 580.250 445.720 585.850 449.325 ;
        RECT 586.690 445.720 589.070 449.325 ;
        RECT 589.910 445.720 592.290 449.325 ;
        RECT 593.130 445.720 598.730 449.325 ;
        RECT 599.570 445.720 601.950 449.325 ;
        RECT 602.790 445.720 608.390 449.325 ;
        RECT 609.230 445.720 611.610 449.325 ;
        RECT 612.450 445.720 614.830 449.325 ;
        RECT 615.670 445.720 621.270 449.325 ;
        RECT 622.110 445.720 624.490 449.325 ;
        RECT 625.330 445.720 627.710 449.325 ;
        RECT 628.550 445.720 634.150 449.325 ;
        RECT 634.990 445.720 637.370 449.325 ;
        RECT 638.210 445.720 640.590 449.325 ;
        RECT 641.430 445.720 647.030 449.325 ;
        RECT 647.870 445.720 650.250 449.325 ;
        RECT 651.090 445.720 653.470 449.325 ;
        RECT 654.310 445.720 659.910 449.325 ;
        RECT 660.750 445.720 663.130 449.325 ;
        RECT 663.970 445.720 666.350 449.325 ;
        RECT 667.190 445.720 672.790 449.325 ;
        RECT 673.630 445.720 676.010 449.325 ;
        RECT 676.850 445.720 679.230 449.325 ;
        RECT 680.070 445.720 685.670 449.325 ;
        RECT 686.510 445.720 688.890 449.325 ;
        RECT 689.730 445.720 692.110 449.325 ;
        RECT 692.950 445.720 698.550 449.325 ;
        RECT 0.100 4.280 699.100 445.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
        RECT 119.790 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 138.270 4.280 ;
        RECT 139.110 0.155 141.490 4.280 ;
        RECT 142.330 0.155 144.710 4.280 ;
        RECT 145.550 0.155 151.150 4.280 ;
        RECT 151.990 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 164.030 4.280 ;
        RECT 164.870 0.155 167.250 4.280 ;
        RECT 168.090 0.155 170.470 4.280 ;
        RECT 171.310 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 189.790 4.280 ;
        RECT 190.630 0.155 193.010 4.280 ;
        RECT 193.850 0.155 196.230 4.280 ;
        RECT 197.070 0.155 202.670 4.280 ;
        RECT 203.510 0.155 205.890 4.280 ;
        RECT 206.730 0.155 212.330 4.280 ;
        RECT 213.170 0.155 215.550 4.280 ;
        RECT 216.390 0.155 218.770 4.280 ;
        RECT 219.610 0.155 225.210 4.280 ;
        RECT 226.050 0.155 228.430 4.280 ;
        RECT 229.270 0.155 231.650 4.280 ;
        RECT 232.490 0.155 238.090 4.280 ;
        RECT 238.930 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 250.970 4.280 ;
        RECT 251.810 0.155 254.190 4.280 ;
        RECT 255.030 0.155 257.410 4.280 ;
        RECT 258.250 0.155 263.850 4.280 ;
        RECT 264.690 0.155 267.070 4.280 ;
        RECT 267.910 0.155 270.290 4.280 ;
        RECT 271.130 0.155 276.730 4.280 ;
        RECT 277.570 0.155 279.950 4.280 ;
        RECT 280.790 0.155 283.170 4.280 ;
        RECT 284.010 0.155 289.610 4.280 ;
        RECT 290.450 0.155 292.830 4.280 ;
        RECT 293.670 0.155 296.050 4.280 ;
        RECT 296.890 0.155 302.490 4.280 ;
        RECT 303.330 0.155 305.710 4.280 ;
        RECT 306.550 0.155 312.150 4.280 ;
        RECT 312.990 0.155 315.370 4.280 ;
        RECT 316.210 0.155 318.590 4.280 ;
        RECT 319.430 0.155 325.030 4.280 ;
        RECT 325.870 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.470 4.280 ;
        RECT 332.310 0.155 337.910 4.280 ;
        RECT 338.750 0.155 341.130 4.280 ;
        RECT 341.970 0.155 344.350 4.280 ;
        RECT 345.190 0.155 350.790 4.280 ;
        RECT 351.630 0.155 354.010 4.280 ;
        RECT 354.850 0.155 357.230 4.280 ;
        RECT 358.070 0.155 363.670 4.280 ;
        RECT 364.510 0.155 366.890 4.280 ;
        RECT 367.730 0.155 370.110 4.280 ;
        RECT 370.950 0.155 376.550 4.280 ;
        RECT 377.390 0.155 379.770 4.280 ;
        RECT 380.610 0.155 382.990 4.280 ;
        RECT 383.830 0.155 389.430 4.280 ;
        RECT 390.270 0.155 392.650 4.280 ;
        RECT 393.490 0.155 395.870 4.280 ;
        RECT 396.710 0.155 402.310 4.280 ;
        RECT 403.150 0.155 405.530 4.280 ;
        RECT 406.370 0.155 411.970 4.280 ;
        RECT 412.810 0.155 415.190 4.280 ;
        RECT 416.030 0.155 418.410 4.280 ;
        RECT 419.250 0.155 424.850 4.280 ;
        RECT 425.690 0.155 428.070 4.280 ;
        RECT 428.910 0.155 431.290 4.280 ;
        RECT 432.130 0.155 437.730 4.280 ;
        RECT 438.570 0.155 440.950 4.280 ;
        RECT 441.790 0.155 444.170 4.280 ;
        RECT 445.010 0.155 450.610 4.280 ;
        RECT 451.450 0.155 453.830 4.280 ;
        RECT 454.670 0.155 457.050 4.280 ;
        RECT 457.890 0.155 463.490 4.280 ;
        RECT 464.330 0.155 466.710 4.280 ;
        RECT 467.550 0.155 469.930 4.280 ;
        RECT 470.770 0.155 476.370 4.280 ;
        RECT 477.210 0.155 479.590 4.280 ;
        RECT 480.430 0.155 482.810 4.280 ;
        RECT 483.650 0.155 489.250 4.280 ;
        RECT 490.090 0.155 492.470 4.280 ;
        RECT 493.310 0.155 495.690 4.280 ;
        RECT 496.530 0.155 502.130 4.280 ;
        RECT 502.970 0.155 505.350 4.280 ;
        RECT 506.190 0.155 508.570 4.280 ;
        RECT 509.410 0.155 515.010 4.280 ;
        RECT 515.850 0.155 518.230 4.280 ;
        RECT 519.070 0.155 524.670 4.280 ;
        RECT 525.510 0.155 527.890 4.280 ;
        RECT 528.730 0.155 531.110 4.280 ;
        RECT 531.950 0.155 537.550 4.280 ;
        RECT 538.390 0.155 540.770 4.280 ;
        RECT 541.610 0.155 543.990 4.280 ;
        RECT 544.830 0.155 550.430 4.280 ;
        RECT 551.270 0.155 553.650 4.280 ;
        RECT 554.490 0.155 556.870 4.280 ;
        RECT 557.710 0.155 563.310 4.280 ;
        RECT 564.150 0.155 566.530 4.280 ;
        RECT 567.370 0.155 569.750 4.280 ;
        RECT 570.590 0.155 576.190 4.280 ;
        RECT 577.030 0.155 579.410 4.280 ;
        RECT 580.250 0.155 582.630 4.280 ;
        RECT 583.470 0.155 589.070 4.280 ;
        RECT 589.910 0.155 592.290 4.280 ;
        RECT 593.130 0.155 595.510 4.280 ;
        RECT 596.350 0.155 601.950 4.280 ;
        RECT 602.790 0.155 605.170 4.280 ;
        RECT 606.010 0.155 608.390 4.280 ;
        RECT 609.230 0.155 614.830 4.280 ;
        RECT 615.670 0.155 618.050 4.280 ;
        RECT 618.890 0.155 624.490 4.280 ;
        RECT 625.330 0.155 627.710 4.280 ;
        RECT 628.550 0.155 630.930 4.280 ;
        RECT 631.770 0.155 637.370 4.280 ;
        RECT 638.210 0.155 640.590 4.280 ;
        RECT 641.430 0.155 643.810 4.280 ;
        RECT 644.650 0.155 650.250 4.280 ;
        RECT 651.090 0.155 653.470 4.280 ;
        RECT 654.310 0.155 656.690 4.280 ;
        RECT 657.530 0.155 663.130 4.280 ;
        RECT 663.970 0.155 666.350 4.280 ;
        RECT 667.190 0.155 669.570 4.280 ;
        RECT 670.410 0.155 676.010 4.280 ;
        RECT 676.850 0.155 679.230 4.280 ;
        RECT 680.070 0.155 682.450 4.280 ;
        RECT 683.290 0.155 688.890 4.280 ;
        RECT 689.730 0.155 692.110 4.280 ;
        RECT 692.950 0.155 695.330 4.280 ;
        RECT 696.170 0.155 699.100 4.280 ;
      LAYER met3 ;
        RECT 4.400 448.440 695.600 449.305 ;
        RECT 4.000 443.040 696.000 448.440 ;
        RECT 4.400 441.640 695.600 443.040 ;
        RECT 4.000 439.640 696.000 441.640 ;
        RECT 4.400 438.240 695.600 439.640 ;
        RECT 4.000 436.240 696.000 438.240 ;
        RECT 4.400 434.840 695.600 436.240 ;
        RECT 4.000 429.440 696.000 434.840 ;
        RECT 4.400 428.040 695.600 429.440 ;
        RECT 4.000 426.040 696.000 428.040 ;
        RECT 4.400 424.640 695.600 426.040 ;
        RECT 4.000 422.640 696.000 424.640 ;
        RECT 4.000 421.240 695.600 422.640 ;
        RECT 4.000 419.240 696.000 421.240 ;
        RECT 4.400 417.840 696.000 419.240 ;
        RECT 4.000 415.840 696.000 417.840 ;
        RECT 4.400 414.440 695.600 415.840 ;
        RECT 4.000 412.440 696.000 414.440 ;
        RECT 4.400 411.040 695.600 412.440 ;
        RECT 4.000 409.040 696.000 411.040 ;
        RECT 4.000 407.640 695.600 409.040 ;
        RECT 4.000 405.640 696.000 407.640 ;
        RECT 4.400 404.240 696.000 405.640 ;
        RECT 4.000 402.240 696.000 404.240 ;
        RECT 4.400 400.840 695.600 402.240 ;
        RECT 4.000 398.840 696.000 400.840 ;
        RECT 4.400 397.440 695.600 398.840 ;
        RECT 4.000 395.440 696.000 397.440 ;
        RECT 4.000 394.040 695.600 395.440 ;
        RECT 4.000 392.040 696.000 394.040 ;
        RECT 4.400 390.640 696.000 392.040 ;
        RECT 4.000 388.640 696.000 390.640 ;
        RECT 4.400 387.240 695.600 388.640 ;
        RECT 4.000 385.240 696.000 387.240 ;
        RECT 4.400 383.840 695.600 385.240 ;
        RECT 4.000 381.840 696.000 383.840 ;
        RECT 4.000 380.440 695.600 381.840 ;
        RECT 4.000 378.440 696.000 380.440 ;
        RECT 4.400 377.040 696.000 378.440 ;
        RECT 4.000 375.040 696.000 377.040 ;
        RECT 4.400 373.640 695.600 375.040 ;
        RECT 4.000 371.640 696.000 373.640 ;
        RECT 4.400 370.240 695.600 371.640 ;
        RECT 4.000 368.240 696.000 370.240 ;
        RECT 4.000 366.840 695.600 368.240 ;
        RECT 4.000 364.840 696.000 366.840 ;
        RECT 4.400 363.440 696.000 364.840 ;
        RECT 4.000 361.440 696.000 363.440 ;
        RECT 4.400 360.040 695.600 361.440 ;
        RECT 4.000 358.040 696.000 360.040 ;
        RECT 4.400 356.640 695.600 358.040 ;
        RECT 4.000 354.640 696.000 356.640 ;
        RECT 4.000 353.240 695.600 354.640 ;
        RECT 4.000 351.240 696.000 353.240 ;
        RECT 4.400 349.840 696.000 351.240 ;
        RECT 4.000 347.840 696.000 349.840 ;
        RECT 4.400 346.440 695.600 347.840 ;
        RECT 4.000 344.440 696.000 346.440 ;
        RECT 4.400 343.040 695.600 344.440 ;
        RECT 4.000 337.640 696.000 343.040 ;
        RECT 4.400 336.240 695.600 337.640 ;
        RECT 4.000 334.240 696.000 336.240 ;
        RECT 4.400 332.840 695.600 334.240 ;
        RECT 4.000 330.840 696.000 332.840 ;
        RECT 4.400 329.440 695.600 330.840 ;
        RECT 4.000 324.040 696.000 329.440 ;
        RECT 4.400 322.640 695.600 324.040 ;
        RECT 4.000 320.640 696.000 322.640 ;
        RECT 4.400 319.240 695.600 320.640 ;
        RECT 4.000 317.240 696.000 319.240 ;
        RECT 4.000 315.840 695.600 317.240 ;
        RECT 4.000 313.840 696.000 315.840 ;
        RECT 4.400 312.440 696.000 313.840 ;
        RECT 4.000 310.440 696.000 312.440 ;
        RECT 4.400 309.040 695.600 310.440 ;
        RECT 4.000 307.040 696.000 309.040 ;
        RECT 4.400 305.640 695.600 307.040 ;
        RECT 4.000 303.640 696.000 305.640 ;
        RECT 4.000 302.240 695.600 303.640 ;
        RECT 4.000 300.240 696.000 302.240 ;
        RECT 4.400 298.840 696.000 300.240 ;
        RECT 4.000 296.840 696.000 298.840 ;
        RECT 4.400 295.440 695.600 296.840 ;
        RECT 4.000 293.440 696.000 295.440 ;
        RECT 4.400 292.040 695.600 293.440 ;
        RECT 4.000 290.040 696.000 292.040 ;
        RECT 4.000 288.640 695.600 290.040 ;
        RECT 4.000 286.640 696.000 288.640 ;
        RECT 4.400 285.240 696.000 286.640 ;
        RECT 4.000 283.240 696.000 285.240 ;
        RECT 4.400 281.840 695.600 283.240 ;
        RECT 4.000 279.840 696.000 281.840 ;
        RECT 4.400 278.440 695.600 279.840 ;
        RECT 4.000 276.440 696.000 278.440 ;
        RECT 4.000 275.040 695.600 276.440 ;
        RECT 4.000 273.040 696.000 275.040 ;
        RECT 4.400 271.640 696.000 273.040 ;
        RECT 4.000 269.640 696.000 271.640 ;
        RECT 4.400 268.240 695.600 269.640 ;
        RECT 4.000 266.240 696.000 268.240 ;
        RECT 4.400 264.840 695.600 266.240 ;
        RECT 4.000 262.840 696.000 264.840 ;
        RECT 4.000 261.440 695.600 262.840 ;
        RECT 4.000 259.440 696.000 261.440 ;
        RECT 4.400 258.040 696.000 259.440 ;
        RECT 4.000 256.040 696.000 258.040 ;
        RECT 4.400 254.640 695.600 256.040 ;
        RECT 4.000 252.640 696.000 254.640 ;
        RECT 4.400 251.240 695.600 252.640 ;
        RECT 4.000 249.240 696.000 251.240 ;
        RECT 4.000 247.840 695.600 249.240 ;
        RECT 4.000 245.840 696.000 247.840 ;
        RECT 4.400 244.440 696.000 245.840 ;
        RECT 4.000 242.440 696.000 244.440 ;
        RECT 4.400 241.040 695.600 242.440 ;
        RECT 4.000 239.040 696.000 241.040 ;
        RECT 4.400 237.640 695.600 239.040 ;
        RECT 4.000 232.240 696.000 237.640 ;
        RECT 4.400 230.840 695.600 232.240 ;
        RECT 4.000 228.840 696.000 230.840 ;
        RECT 4.400 227.440 695.600 228.840 ;
        RECT 4.000 225.440 696.000 227.440 ;
        RECT 4.400 224.040 695.600 225.440 ;
        RECT 4.000 218.640 696.000 224.040 ;
        RECT 4.400 217.240 695.600 218.640 ;
        RECT 4.000 215.240 696.000 217.240 ;
        RECT 4.400 213.840 695.600 215.240 ;
        RECT 4.000 211.840 696.000 213.840 ;
        RECT 4.000 210.440 695.600 211.840 ;
        RECT 4.000 208.440 696.000 210.440 ;
        RECT 4.400 207.040 696.000 208.440 ;
        RECT 4.000 205.040 696.000 207.040 ;
        RECT 4.400 203.640 695.600 205.040 ;
        RECT 4.000 201.640 696.000 203.640 ;
        RECT 4.400 200.240 695.600 201.640 ;
        RECT 4.000 198.240 696.000 200.240 ;
        RECT 4.000 196.840 695.600 198.240 ;
        RECT 4.000 194.840 696.000 196.840 ;
        RECT 4.400 193.440 696.000 194.840 ;
        RECT 4.000 191.440 696.000 193.440 ;
        RECT 4.400 190.040 695.600 191.440 ;
        RECT 4.000 188.040 696.000 190.040 ;
        RECT 4.400 186.640 695.600 188.040 ;
        RECT 4.000 184.640 696.000 186.640 ;
        RECT 4.000 183.240 695.600 184.640 ;
        RECT 4.000 181.240 696.000 183.240 ;
        RECT 4.400 179.840 696.000 181.240 ;
        RECT 4.000 177.840 696.000 179.840 ;
        RECT 4.400 176.440 695.600 177.840 ;
        RECT 4.000 174.440 696.000 176.440 ;
        RECT 4.400 173.040 695.600 174.440 ;
        RECT 4.000 171.040 696.000 173.040 ;
        RECT 4.000 169.640 695.600 171.040 ;
        RECT 4.000 167.640 696.000 169.640 ;
        RECT 4.400 166.240 696.000 167.640 ;
        RECT 4.000 164.240 696.000 166.240 ;
        RECT 4.400 162.840 695.600 164.240 ;
        RECT 4.000 160.840 696.000 162.840 ;
        RECT 4.400 159.440 695.600 160.840 ;
        RECT 4.000 157.440 696.000 159.440 ;
        RECT 4.000 156.040 695.600 157.440 ;
        RECT 4.000 154.040 696.000 156.040 ;
        RECT 4.400 152.640 696.000 154.040 ;
        RECT 4.000 150.640 696.000 152.640 ;
        RECT 4.400 149.240 695.600 150.640 ;
        RECT 4.000 147.240 696.000 149.240 ;
        RECT 4.400 145.840 695.600 147.240 ;
        RECT 4.000 143.840 696.000 145.840 ;
        RECT 4.000 142.440 695.600 143.840 ;
        RECT 4.000 140.440 696.000 142.440 ;
        RECT 4.400 139.040 696.000 140.440 ;
        RECT 4.000 137.040 696.000 139.040 ;
        RECT 4.400 135.640 695.600 137.040 ;
        RECT 4.000 133.640 696.000 135.640 ;
        RECT 4.400 132.240 695.600 133.640 ;
        RECT 4.000 130.240 696.000 132.240 ;
        RECT 4.000 128.840 695.600 130.240 ;
        RECT 4.000 126.840 696.000 128.840 ;
        RECT 4.400 125.440 696.000 126.840 ;
        RECT 4.000 123.440 696.000 125.440 ;
        RECT 4.400 122.040 695.600 123.440 ;
        RECT 4.000 120.040 696.000 122.040 ;
        RECT 4.400 118.640 695.600 120.040 ;
        RECT 4.000 113.240 696.000 118.640 ;
        RECT 4.400 111.840 695.600 113.240 ;
        RECT 4.000 109.840 696.000 111.840 ;
        RECT 4.400 108.440 695.600 109.840 ;
        RECT 4.000 106.440 696.000 108.440 ;
        RECT 4.000 105.040 695.600 106.440 ;
        RECT 4.000 103.040 696.000 105.040 ;
        RECT 4.400 101.640 696.000 103.040 ;
        RECT 4.000 99.640 696.000 101.640 ;
        RECT 4.400 98.240 695.600 99.640 ;
        RECT 4.000 96.240 696.000 98.240 ;
        RECT 4.400 94.840 695.600 96.240 ;
        RECT 4.000 92.840 696.000 94.840 ;
        RECT 4.000 91.440 695.600 92.840 ;
        RECT 4.000 89.440 696.000 91.440 ;
        RECT 4.400 88.040 696.000 89.440 ;
        RECT 4.000 86.040 696.000 88.040 ;
        RECT 4.400 84.640 695.600 86.040 ;
        RECT 4.000 82.640 696.000 84.640 ;
        RECT 4.400 81.240 695.600 82.640 ;
        RECT 4.000 79.240 696.000 81.240 ;
        RECT 4.000 77.840 695.600 79.240 ;
        RECT 4.000 75.840 696.000 77.840 ;
        RECT 4.400 74.440 696.000 75.840 ;
        RECT 4.000 72.440 696.000 74.440 ;
        RECT 4.400 71.040 695.600 72.440 ;
        RECT 4.000 69.040 696.000 71.040 ;
        RECT 4.400 67.640 695.600 69.040 ;
        RECT 4.000 65.640 696.000 67.640 ;
        RECT 4.000 64.240 695.600 65.640 ;
        RECT 4.000 62.240 696.000 64.240 ;
        RECT 4.400 60.840 696.000 62.240 ;
        RECT 4.000 58.840 696.000 60.840 ;
        RECT 4.400 57.440 695.600 58.840 ;
        RECT 4.000 55.440 696.000 57.440 ;
        RECT 4.400 54.040 695.600 55.440 ;
        RECT 4.000 52.040 696.000 54.040 ;
        RECT 4.000 50.640 695.600 52.040 ;
        RECT 4.000 48.640 696.000 50.640 ;
        RECT 4.400 47.240 696.000 48.640 ;
        RECT 4.000 45.240 696.000 47.240 ;
        RECT 4.400 43.840 695.600 45.240 ;
        RECT 4.000 41.840 696.000 43.840 ;
        RECT 4.400 40.440 695.600 41.840 ;
        RECT 4.000 38.440 696.000 40.440 ;
        RECT 4.000 37.040 695.600 38.440 ;
        RECT 4.000 35.040 696.000 37.040 ;
        RECT 4.400 33.640 696.000 35.040 ;
        RECT 4.000 31.640 696.000 33.640 ;
        RECT 4.400 30.240 695.600 31.640 ;
        RECT 4.000 28.240 696.000 30.240 ;
        RECT 4.400 26.840 695.600 28.240 ;
        RECT 4.000 24.840 696.000 26.840 ;
        RECT 4.000 23.440 695.600 24.840 ;
        RECT 4.000 21.440 696.000 23.440 ;
        RECT 4.400 20.040 696.000 21.440 ;
        RECT 4.000 18.040 696.000 20.040 ;
        RECT 4.400 16.640 695.600 18.040 ;
        RECT 4.000 14.640 696.000 16.640 ;
        RECT 4.400 13.240 695.600 14.640 ;
        RECT 4.000 7.840 696.000 13.240 ;
        RECT 4.400 6.440 695.600 7.840 ;
        RECT 4.000 4.440 696.000 6.440 ;
        RECT 4.400 3.040 695.600 4.440 ;
        RECT 4.000 1.040 696.000 3.040 ;
        RECT 4.000 0.175 695.600 1.040 ;
      LAYER met4 ;
        RECT 94.135 11.735 97.440 430.945 ;
        RECT 99.840 11.735 174.240 430.945 ;
        RECT 176.640 11.735 251.040 430.945 ;
        RECT 253.440 11.735 327.840 430.945 ;
        RECT 330.240 11.735 404.640 430.945 ;
        RECT 407.040 11.735 481.440 430.945 ;
        RECT 483.840 11.735 558.240 430.945 ;
        RECT 560.640 11.735 579.305 430.945 ;
  END
END l1dcache
END LIBRARY

