magic
tech sky130B
magscale 1 2
timestamp 1662997958
<< obsli1 >>
rect 1104 2159 118864 27761
<< obsm1 >>
rect 14 1096 119862 28144
<< metal2 >>
rect 18 29200 74 30000
rect 662 29200 718 30000
rect 1306 29200 1362 30000
rect 2594 29200 2650 30000
rect 3238 29200 3294 30000
rect 4526 29200 4582 30000
rect 5170 29200 5226 30000
rect 6458 29200 6514 30000
rect 7102 29200 7158 30000
rect 7746 29200 7802 30000
rect 9034 29200 9090 30000
rect 9678 29200 9734 30000
rect 10966 29200 11022 30000
rect 11610 29200 11666 30000
rect 12254 29200 12310 30000
rect 13542 29200 13598 30000
rect 14186 29200 14242 30000
rect 15474 29200 15530 30000
rect 16118 29200 16174 30000
rect 17406 29200 17462 30000
rect 18050 29200 18106 30000
rect 18694 29200 18750 30000
rect 19982 29200 20038 30000
rect 20626 29200 20682 30000
rect 21914 29200 21970 30000
rect 22558 29200 22614 30000
rect 23846 29200 23902 30000
rect 24490 29200 24546 30000
rect 25134 29200 25190 30000
rect 26422 29200 26478 30000
rect 27066 29200 27122 30000
rect 28354 29200 28410 30000
rect 28998 29200 29054 30000
rect 29642 29200 29698 30000
rect 30930 29200 30986 30000
rect 31574 29200 31630 30000
rect 32862 29200 32918 30000
rect 33506 29200 33562 30000
rect 34794 29200 34850 30000
rect 35438 29200 35494 30000
rect 36082 29200 36138 30000
rect 37370 29200 37426 30000
rect 38014 29200 38070 30000
rect 39302 29200 39358 30000
rect 39946 29200 40002 30000
rect 41234 29200 41290 30000
rect 41878 29200 41934 30000
rect 42522 29200 42578 30000
rect 43810 29200 43866 30000
rect 44454 29200 44510 30000
rect 45742 29200 45798 30000
rect 46386 29200 46442 30000
rect 47030 29200 47086 30000
rect 48318 29200 48374 30000
rect 48962 29200 49018 30000
rect 50250 29200 50306 30000
rect 50894 29200 50950 30000
rect 52182 29200 52238 30000
rect 52826 29200 52882 30000
rect 53470 29200 53526 30000
rect 54758 29200 54814 30000
rect 55402 29200 55458 30000
rect 56690 29200 56746 30000
rect 57334 29200 57390 30000
rect 58622 29200 58678 30000
rect 59266 29200 59322 30000
rect 59910 29200 59966 30000
rect 61198 29200 61254 30000
rect 61842 29200 61898 30000
rect 63130 29200 63186 30000
rect 63774 29200 63830 30000
rect 64418 29200 64474 30000
rect 65706 29200 65762 30000
rect 66350 29200 66406 30000
rect 67638 29200 67694 30000
rect 68282 29200 68338 30000
rect 69570 29200 69626 30000
rect 70214 29200 70270 30000
rect 70858 29200 70914 30000
rect 72146 29200 72202 30000
rect 72790 29200 72846 30000
rect 74078 29200 74134 30000
rect 74722 29200 74778 30000
rect 76010 29200 76066 30000
rect 76654 29200 76710 30000
rect 77298 29200 77354 30000
rect 78586 29200 78642 30000
rect 79230 29200 79286 30000
rect 80518 29200 80574 30000
rect 81162 29200 81218 30000
rect 82450 29200 82506 30000
rect 83094 29200 83150 30000
rect 83738 29200 83794 30000
rect 85026 29200 85082 30000
rect 85670 29200 85726 30000
rect 86958 29200 87014 30000
rect 87602 29200 87658 30000
rect 88246 29200 88302 30000
rect 89534 29200 89590 30000
rect 90178 29200 90234 30000
rect 91466 29200 91522 30000
rect 92110 29200 92166 30000
rect 93398 29200 93454 30000
rect 94042 29200 94098 30000
rect 94686 29200 94742 30000
rect 95974 29200 96030 30000
rect 96618 29200 96674 30000
rect 97906 29200 97962 30000
rect 98550 29200 98606 30000
rect 99838 29200 99894 30000
rect 100482 29200 100538 30000
rect 101126 29200 101182 30000
rect 102414 29200 102470 30000
rect 103058 29200 103114 30000
rect 104346 29200 104402 30000
rect 104990 29200 105046 30000
rect 105634 29200 105690 30000
rect 106922 29200 106978 30000
rect 107566 29200 107622 30000
rect 108854 29200 108910 30000
rect 109498 29200 109554 30000
rect 110786 29200 110842 30000
rect 111430 29200 111486 30000
rect 112074 29200 112130 30000
rect 113362 29200 113418 30000
rect 114006 29200 114062 30000
rect 115294 29200 115350 30000
rect 115938 29200 115994 30000
rect 117226 29200 117282 30000
rect 117870 29200 117926 30000
rect 118514 29200 118570 30000
rect 119802 29200 119858 30000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92754 0 92810 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 100482 0 100538 800
rect 101126 0 101182 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 104346 0 104402 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106922 0 106978 800
rect 107566 0 107622 800
rect 108854 0 108910 800
rect 109498 0 109554 800
rect 110786 0 110842 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 115294 0 115350 800
rect 115938 0 115994 800
rect 116582 0 116638 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119802 0 119858 800
<< obsm2 >>
rect 130 29144 606 29322
rect 774 29144 1250 29322
rect 1418 29144 2538 29322
rect 2706 29144 3182 29322
rect 3350 29144 4470 29322
rect 4638 29144 5114 29322
rect 5282 29144 6402 29322
rect 6570 29144 7046 29322
rect 7214 29144 7690 29322
rect 7858 29144 8978 29322
rect 9146 29144 9622 29322
rect 9790 29144 10910 29322
rect 11078 29144 11554 29322
rect 11722 29144 12198 29322
rect 12366 29144 13486 29322
rect 13654 29144 14130 29322
rect 14298 29144 15418 29322
rect 15586 29144 16062 29322
rect 16230 29144 17350 29322
rect 17518 29144 17994 29322
rect 18162 29144 18638 29322
rect 18806 29144 19926 29322
rect 20094 29144 20570 29322
rect 20738 29144 21858 29322
rect 22026 29144 22502 29322
rect 22670 29144 23790 29322
rect 23958 29144 24434 29322
rect 24602 29144 25078 29322
rect 25246 29144 26366 29322
rect 26534 29144 27010 29322
rect 27178 29144 28298 29322
rect 28466 29144 28942 29322
rect 29110 29144 29586 29322
rect 29754 29144 30874 29322
rect 31042 29144 31518 29322
rect 31686 29144 32806 29322
rect 32974 29144 33450 29322
rect 33618 29144 34738 29322
rect 34906 29144 35382 29322
rect 35550 29144 36026 29322
rect 36194 29144 37314 29322
rect 37482 29144 37958 29322
rect 38126 29144 39246 29322
rect 39414 29144 39890 29322
rect 40058 29144 41178 29322
rect 41346 29144 41822 29322
rect 41990 29144 42466 29322
rect 42634 29144 43754 29322
rect 43922 29144 44398 29322
rect 44566 29144 45686 29322
rect 45854 29144 46330 29322
rect 46498 29144 46974 29322
rect 47142 29144 48262 29322
rect 48430 29144 48906 29322
rect 49074 29144 50194 29322
rect 50362 29144 50838 29322
rect 51006 29144 52126 29322
rect 52294 29144 52770 29322
rect 52938 29144 53414 29322
rect 53582 29144 54702 29322
rect 54870 29144 55346 29322
rect 55514 29144 56634 29322
rect 56802 29144 57278 29322
rect 57446 29144 58566 29322
rect 58734 29144 59210 29322
rect 59378 29144 59854 29322
rect 60022 29144 61142 29322
rect 61310 29144 61786 29322
rect 61954 29144 63074 29322
rect 63242 29144 63718 29322
rect 63886 29144 64362 29322
rect 64530 29144 65650 29322
rect 65818 29144 66294 29322
rect 66462 29144 67582 29322
rect 67750 29144 68226 29322
rect 68394 29144 69514 29322
rect 69682 29144 70158 29322
rect 70326 29144 70802 29322
rect 70970 29144 72090 29322
rect 72258 29144 72734 29322
rect 72902 29144 74022 29322
rect 74190 29144 74666 29322
rect 74834 29144 75954 29322
rect 76122 29144 76598 29322
rect 76766 29144 77242 29322
rect 77410 29144 78530 29322
rect 78698 29144 79174 29322
rect 79342 29144 80462 29322
rect 80630 29144 81106 29322
rect 81274 29144 82394 29322
rect 82562 29144 83038 29322
rect 83206 29144 83682 29322
rect 83850 29144 84970 29322
rect 85138 29144 85614 29322
rect 85782 29144 86902 29322
rect 87070 29144 87546 29322
rect 87714 29144 88190 29322
rect 88358 29144 89478 29322
rect 89646 29144 90122 29322
rect 90290 29144 91410 29322
rect 91578 29144 92054 29322
rect 92222 29144 93342 29322
rect 93510 29144 93986 29322
rect 94154 29144 94630 29322
rect 94798 29144 95918 29322
rect 96086 29144 96562 29322
rect 96730 29144 97850 29322
rect 98018 29144 98494 29322
rect 98662 29144 99782 29322
rect 99950 29144 100426 29322
rect 100594 29144 101070 29322
rect 101238 29144 102358 29322
rect 102526 29144 103002 29322
rect 103170 29144 104290 29322
rect 104458 29144 104934 29322
rect 105102 29144 105578 29322
rect 105746 29144 106866 29322
rect 107034 29144 107510 29322
rect 107678 29144 108798 29322
rect 108966 29144 109442 29322
rect 109610 29144 110730 29322
rect 110898 29144 111374 29322
rect 111542 29144 112018 29322
rect 112186 29144 113306 29322
rect 113474 29144 113950 29322
rect 114118 29144 115238 29322
rect 115406 29144 115882 29322
rect 116050 29144 117170 29322
rect 117338 29144 117814 29322
rect 117982 29144 118458 29322
rect 118626 29144 119746 29322
rect 20 856 119856 29144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 2538 856
rect 2706 31 3182 856
rect 3350 31 4470 856
rect 4638 31 5114 856
rect 5282 31 5758 856
rect 5926 31 7046 856
rect 7214 31 7690 856
rect 7858 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 13486 856
rect 13654 31 14130 856
rect 14298 31 15418 856
rect 15586 31 16062 856
rect 16230 31 17350 856
rect 17518 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19926 856
rect 20094 31 20570 856
rect 20738 31 21858 856
rect 22026 31 22502 856
rect 22670 31 23146 856
rect 23314 31 24434 856
rect 24602 31 25078 856
rect 25246 31 26366 856
rect 26534 31 27010 856
rect 27178 31 28298 856
rect 28466 31 28942 856
rect 29110 31 29586 856
rect 29754 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36026 856
rect 36194 31 37314 856
rect 37482 31 37958 856
rect 38126 31 39246 856
rect 39414 31 39890 856
rect 40058 31 40534 856
rect 40702 31 41822 856
rect 41990 31 42466 856
rect 42634 31 43754 856
rect 43922 31 44398 856
rect 44566 31 45686 856
rect 45854 31 46330 856
rect 46498 31 46974 856
rect 47142 31 48262 856
rect 48430 31 48906 856
rect 49074 31 50194 856
rect 50362 31 50838 856
rect 51006 31 52126 856
rect 52294 31 52770 856
rect 52938 31 53414 856
rect 53582 31 54702 856
rect 54870 31 55346 856
rect 55514 31 56634 856
rect 56802 31 57278 856
rect 57446 31 57922 856
rect 58090 31 59210 856
rect 59378 31 59854 856
rect 60022 31 61142 856
rect 61310 31 61786 856
rect 61954 31 63074 856
rect 63242 31 63718 856
rect 63886 31 64362 856
rect 64530 31 65650 856
rect 65818 31 66294 856
rect 66462 31 67582 856
rect 67750 31 68226 856
rect 68394 31 69514 856
rect 69682 31 70158 856
rect 70326 31 70802 856
rect 70970 31 72090 856
rect 72258 31 72734 856
rect 72902 31 74022 856
rect 74190 31 74666 856
rect 74834 31 75310 856
rect 75478 31 76598 856
rect 76766 31 77242 856
rect 77410 31 78530 856
rect 78698 31 79174 856
rect 79342 31 80462 856
rect 80630 31 81106 856
rect 81274 31 81750 856
rect 81918 31 83038 856
rect 83206 31 83682 856
rect 83850 31 84970 856
rect 85138 31 85614 856
rect 85782 31 86902 856
rect 87070 31 87546 856
rect 87714 31 88190 856
rect 88358 31 89478 856
rect 89646 31 90122 856
rect 90290 31 91410 856
rect 91578 31 92054 856
rect 92222 31 92698 856
rect 92866 31 93986 856
rect 94154 31 94630 856
rect 94798 31 95918 856
rect 96086 31 96562 856
rect 96730 31 97850 856
rect 98018 31 98494 856
rect 98662 31 99138 856
rect 99306 31 100426 856
rect 100594 31 101070 856
rect 101238 31 102358 856
rect 102526 31 103002 856
rect 103170 31 104290 856
rect 104458 31 104934 856
rect 105102 31 105578 856
rect 105746 31 106866 856
rect 107034 31 107510 856
rect 107678 31 108798 856
rect 108966 31 109442 856
rect 109610 31 110730 856
rect 110898 31 111374 856
rect 111542 31 112018 856
rect 112186 31 113306 856
rect 113474 31 113950 856
rect 114118 31 115238 856
rect 115406 31 115882 856
rect 116050 31 116526 856
rect 116694 31 117814 856
rect 117982 31 118458 856
rect 118626 31 119746 856
<< metal3 >>
rect 119200 29248 120000 29368
rect 0 28568 800 28688
rect 0 27888 800 28008
rect 119200 27888 120000 28008
rect 119200 27208 120000 27328
rect 0 26528 800 26648
rect 119200 26528 120000 26648
rect 0 25848 800 25968
rect 119200 25168 120000 25288
rect 0 24488 800 24608
rect 119200 24488 120000 24608
rect 0 23808 800 23928
rect 0 23128 800 23248
rect 119200 23128 120000 23248
rect 119200 22448 120000 22568
rect 0 21768 800 21888
rect 0 21088 800 21208
rect 119200 21088 120000 21208
rect 119200 20408 120000 20528
rect 0 19728 800 19848
rect 119200 19728 120000 19848
rect 0 19048 800 19168
rect 0 18368 800 18488
rect 119200 18368 120000 18488
rect 119200 17688 120000 17808
rect 0 17008 800 17128
rect 0 16328 800 16448
rect 119200 16328 120000 16448
rect 119200 15648 120000 15768
rect 0 14968 800 15088
rect 0 14288 800 14408
rect 119200 14288 120000 14408
rect 119200 13608 120000 13728
rect 0 12928 800 13048
rect 119200 12928 120000 13048
rect 0 12248 800 12368
rect 0 11568 800 11688
rect 119200 11568 120000 11688
rect 119200 10888 120000 11008
rect 0 10208 800 10328
rect 0 9528 800 9648
rect 119200 9528 120000 9648
rect 119200 8848 120000 8968
rect 0 8168 800 8288
rect 119200 8168 120000 8288
rect 0 7488 800 7608
rect 119200 6808 120000 6928
rect 0 6128 800 6248
rect 119200 6128 120000 6248
rect 0 5448 800 5568
rect 0 4768 800 4888
rect 119200 4768 120000 4888
rect 119200 4088 120000 4208
rect 0 3408 800 3528
rect 0 2728 800 2848
rect 119200 2728 120000 2848
rect 119200 2048 120000 2168
rect 0 1368 800 1488
rect 119200 1368 120000 1488
rect 0 688 800 808
rect 119200 8 120000 128
<< obsm3 >>
rect 800 29168 119120 29338
rect 800 28768 119200 29168
rect 880 28488 119200 28768
rect 800 28088 119200 28488
rect 880 27808 119120 28088
rect 800 27408 119200 27808
rect 800 27128 119120 27408
rect 800 26728 119200 27128
rect 880 26448 119120 26728
rect 800 26048 119200 26448
rect 880 25768 119200 26048
rect 800 25368 119200 25768
rect 800 25088 119120 25368
rect 800 24688 119200 25088
rect 880 24408 119120 24688
rect 800 24008 119200 24408
rect 880 23728 119200 24008
rect 800 23328 119200 23728
rect 880 23048 119120 23328
rect 800 22648 119200 23048
rect 800 22368 119120 22648
rect 800 21968 119200 22368
rect 880 21688 119200 21968
rect 800 21288 119200 21688
rect 880 21008 119120 21288
rect 800 20608 119200 21008
rect 800 20328 119120 20608
rect 800 19928 119200 20328
rect 880 19648 119120 19928
rect 800 19248 119200 19648
rect 880 18968 119200 19248
rect 800 18568 119200 18968
rect 880 18288 119120 18568
rect 800 17888 119200 18288
rect 800 17608 119120 17888
rect 800 17208 119200 17608
rect 880 16928 119200 17208
rect 800 16528 119200 16928
rect 880 16248 119120 16528
rect 800 15848 119200 16248
rect 800 15568 119120 15848
rect 800 15168 119200 15568
rect 880 14888 119200 15168
rect 800 14488 119200 14888
rect 880 14208 119120 14488
rect 800 13808 119200 14208
rect 800 13528 119120 13808
rect 800 13128 119200 13528
rect 880 12848 119120 13128
rect 800 12448 119200 12848
rect 880 12168 119200 12448
rect 800 11768 119200 12168
rect 880 11488 119120 11768
rect 800 11088 119200 11488
rect 800 10808 119120 11088
rect 800 10408 119200 10808
rect 880 10128 119200 10408
rect 800 9728 119200 10128
rect 880 9448 119120 9728
rect 800 9048 119200 9448
rect 800 8768 119120 9048
rect 800 8368 119200 8768
rect 880 8088 119120 8368
rect 800 7688 119200 8088
rect 880 7408 119200 7688
rect 800 7008 119200 7408
rect 800 6728 119120 7008
rect 800 6328 119200 6728
rect 880 6048 119120 6328
rect 800 5648 119200 6048
rect 880 5368 119200 5648
rect 800 4968 119200 5368
rect 880 4688 119120 4968
rect 800 4288 119200 4688
rect 800 4008 119120 4288
rect 800 3608 119200 4008
rect 880 3328 119200 3608
rect 800 2928 119200 3328
rect 880 2648 119120 2928
rect 800 2248 119200 2648
rect 800 1968 119120 2248
rect 800 1568 119200 1968
rect 880 1288 119120 1568
rect 800 888 119200 1288
rect 880 608 119200 888
rect 800 208 119200 608
rect 800 35 119120 208
<< metal4 >>
rect 15668 2128 15988 27792
rect 30392 2128 30712 27792
rect 45116 2128 45436 27792
rect 59840 2128 60160 27792
rect 74564 2128 74884 27792
rect 89288 2128 89608 27792
rect 104012 2128 104332 27792
<< obsm4 >>
rect 70347 26283 70781 26890
<< labels >>
rlabel metal3 s 119200 8848 120000 8968 6 clk
port 1 nsew signal input
rlabel metal2 s 18694 29200 18750 30000 6 m2_dcache_wbd_ack_o
port 2 nsew signal output
rlabel metal2 s 74722 29200 74778 30000 6 m2_dcache_wbd_adr_i[0]
port 3 nsew signal input
rlabel metal2 s 6458 29200 6514 30000 6 m2_dcache_wbd_adr_i[10]
port 4 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 m2_dcache_wbd_adr_i[11]
port 5 nsew signal input
rlabel metal2 s 39302 29200 39358 30000 6 m2_dcache_wbd_adr_i[12]
port 6 nsew signal input
rlabel metal2 s 43810 29200 43866 30000 6 m2_dcache_wbd_adr_i[13]
port 7 nsew signal input
rlabel metal2 s 10966 29200 11022 30000 6 m2_dcache_wbd_adr_i[14]
port 8 nsew signal input
rlabel metal2 s 28354 29200 28410 30000 6 m2_dcache_wbd_adr_i[15]
port 9 nsew signal input
rlabel metal2 s 33506 29200 33562 30000 6 m2_dcache_wbd_adr_i[16]
port 10 nsew signal input
rlabel metal3 s 119200 16328 120000 16448 6 m2_dcache_wbd_adr_i[17]
port 11 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 m2_dcache_wbd_adr_i[18]
port 12 nsew signal input
rlabel metal2 s 66350 29200 66406 30000 6 m2_dcache_wbd_adr_i[19]
port 13 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 m2_dcache_wbd_adr_i[1]
port 14 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 m2_dcache_wbd_adr_i[20]
port 15 nsew signal input
rlabel metal3 s 119200 23128 120000 23248 6 m2_dcache_wbd_adr_i[21]
port 16 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 m2_dcache_wbd_adr_i[22]
port 17 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 m2_dcache_wbd_adr_i[23]
port 18 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 m2_dcache_wbd_adr_i[24]
port 19 nsew signal input
rlabel metal2 s 102414 29200 102470 30000 6 m2_dcache_wbd_adr_i[25]
port 20 nsew signal input
rlabel metal2 s 59266 29200 59322 30000 6 m2_dcache_wbd_adr_i[26]
port 21 nsew signal input
rlabel metal3 s 0 688 800 808 6 m2_dcache_wbd_adr_i[27]
port 22 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 m2_dcache_wbd_adr_i[28]
port 23 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 m2_dcache_wbd_adr_i[29]
port 24 nsew signal input
rlabel metal2 s 115938 29200 115994 30000 6 m2_dcache_wbd_adr_i[2]
port 25 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 m2_dcache_wbd_adr_i[30]
port 26 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 m2_dcache_wbd_adr_i[31]
port 27 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 m2_dcache_wbd_adr_i[3]
port 28 nsew signal input
rlabel metal3 s 119200 2048 120000 2168 6 m2_dcache_wbd_adr_i[4]
port 29 nsew signal input
rlabel metal2 s 34794 29200 34850 30000 6 m2_dcache_wbd_adr_i[5]
port 30 nsew signal input
rlabel metal2 s 23846 29200 23902 30000 6 m2_dcache_wbd_adr_i[6]
port 31 nsew signal input
rlabel metal3 s 119200 4088 120000 4208 6 m2_dcache_wbd_adr_i[7]
port 32 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 m2_dcache_wbd_adr_i[8]
port 33 nsew signal input
rlabel metal2 s 2594 29200 2650 30000 6 m2_dcache_wbd_adr_i[9]
port 34 nsew signal input
rlabel metal2 s 662 0 718 800 6 m2_dcache_wbd_cyc_i
port 35 nsew signal input
rlabel metal3 s 119200 21088 120000 21208 6 m2_dcache_wbd_dat_i[0]
port 36 nsew signal input
rlabel metal2 s 72790 29200 72846 30000 6 m2_dcache_wbd_dat_i[10]
port 37 nsew signal input
rlabel metal2 s 65706 29200 65762 30000 6 m2_dcache_wbd_dat_i[11]
port 38 nsew signal input
rlabel metal2 s 68282 29200 68338 30000 6 m2_dcache_wbd_dat_i[12]
port 39 nsew signal input
rlabel metal2 s 37370 29200 37426 30000 6 m2_dcache_wbd_dat_i[13]
port 40 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 m2_dcache_wbd_dat_i[14]
port 41 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 m2_dcache_wbd_dat_i[15]
port 42 nsew signal input
rlabel metal2 s 28998 29200 29054 30000 6 m2_dcache_wbd_dat_i[16]
port 43 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 m2_dcache_wbd_dat_i[17]
port 44 nsew signal input
rlabel metal2 s 53470 29200 53526 30000 6 m2_dcache_wbd_dat_i[18]
port 45 nsew signal input
rlabel metal2 s 9034 29200 9090 30000 6 m2_dcache_wbd_dat_i[19]
port 46 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 m2_dcache_wbd_dat_i[1]
port 47 nsew signal input
rlabel metal2 s 5170 29200 5226 30000 6 m2_dcache_wbd_dat_i[20]
port 48 nsew signal input
rlabel metal2 s 13542 29200 13598 30000 6 m2_dcache_wbd_dat_i[21]
port 49 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 m2_dcache_wbd_dat_i[22]
port 50 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 m2_dcache_wbd_dat_i[23]
port 51 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 m2_dcache_wbd_dat_i[24]
port 52 nsew signal input
rlabel metal2 s 15474 29200 15530 30000 6 m2_dcache_wbd_dat_i[25]
port 53 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 m2_dcache_wbd_dat_i[26]
port 54 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 m2_dcache_wbd_dat_i[27]
port 55 nsew signal input
rlabel metal2 s 78586 29200 78642 30000 6 m2_dcache_wbd_dat_i[28]
port 56 nsew signal input
rlabel metal2 s 27066 29200 27122 30000 6 m2_dcache_wbd_dat_i[29]
port 57 nsew signal input
rlabel metal2 s 70858 29200 70914 30000 6 m2_dcache_wbd_dat_i[2]
port 58 nsew signal input
rlabel metal2 s 85670 29200 85726 30000 6 m2_dcache_wbd_dat_i[30]
port 59 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 m2_dcache_wbd_dat_i[31]
port 60 nsew signal input
rlabel metal2 s 63130 29200 63186 30000 6 m2_dcache_wbd_dat_i[3]
port 61 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 m2_dcache_wbd_dat_i[4]
port 62 nsew signal input
rlabel metal2 s 16118 29200 16174 30000 6 m2_dcache_wbd_dat_i[5]
port 63 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 m2_dcache_wbd_dat_i[6]
port 64 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 m2_dcache_wbd_dat_i[7]
port 65 nsew signal input
rlabel metal2 s 106922 29200 106978 30000 6 m2_dcache_wbd_dat_i[8]
port 66 nsew signal input
rlabel metal3 s 119200 2728 120000 2848 6 m2_dcache_wbd_dat_i[9]
port 67 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 m2_dcache_wbd_dat_o[0]
port 68 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 m2_dcache_wbd_dat_o[10]
port 69 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 m2_dcache_wbd_dat_o[11]
port 70 nsew signal output
rlabel metal2 s 7746 29200 7802 30000 6 m2_dcache_wbd_dat_o[12]
port 71 nsew signal output
rlabel metal2 s 57334 29200 57390 30000 6 m2_dcache_wbd_dat_o[13]
port 72 nsew signal output
rlabel metal2 s 42522 29200 42578 30000 6 m2_dcache_wbd_dat_o[14]
port 73 nsew signal output
rlabel metal2 s 104346 29200 104402 30000 6 m2_dcache_wbd_dat_o[15]
port 74 nsew signal output
rlabel metal2 s 81162 29200 81218 30000 6 m2_dcache_wbd_dat_o[16]
port 75 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 m2_dcache_wbd_dat_o[17]
port 76 nsew signal output
rlabel metal2 s 35438 29200 35494 30000 6 m2_dcache_wbd_dat_o[18]
port 77 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 m2_dcache_wbd_dat_o[19]
port 78 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 m2_dcache_wbd_dat_o[1]
port 79 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 m2_dcache_wbd_dat_o[20]
port 80 nsew signal output
rlabel metal2 s 108854 29200 108910 30000 6 m2_dcache_wbd_dat_o[21]
port 81 nsew signal output
rlabel metal2 s 45742 29200 45798 30000 6 m2_dcache_wbd_dat_o[22]
port 82 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 m2_dcache_wbd_dat_o[23]
port 83 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 m2_dcache_wbd_dat_o[24]
port 84 nsew signal output
rlabel metal2 s 9678 29200 9734 30000 6 m2_dcache_wbd_dat_o[25]
port 85 nsew signal output
rlabel metal2 s 93398 29200 93454 30000 6 m2_dcache_wbd_dat_o[26]
port 86 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 m2_dcache_wbd_dat_o[27]
port 87 nsew signal output
rlabel metal2 s 38014 29200 38070 30000 6 m2_dcache_wbd_dat_o[28]
port 88 nsew signal output
rlabel metal2 s 82450 29200 82506 30000 6 m2_dcache_wbd_dat_o[29]
port 89 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 m2_dcache_wbd_dat_o[2]
port 90 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 m2_dcache_wbd_dat_o[30]
port 91 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 m2_dcache_wbd_dat_o[31]
port 92 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 m2_dcache_wbd_dat_o[3]
port 93 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 m2_dcache_wbd_dat_o[4]
port 94 nsew signal output
rlabel metal2 s 67638 29200 67694 30000 6 m2_dcache_wbd_dat_o[5]
port 95 nsew signal output
rlabel metal3 s 119200 25168 120000 25288 6 m2_dcache_wbd_dat_o[6]
port 96 nsew signal output
rlabel metal2 s 52826 29200 52882 30000 6 m2_dcache_wbd_dat_o[7]
port 97 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 m2_dcache_wbd_dat_o[8]
port 98 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 m2_dcache_wbd_dat_o[9]
port 99 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 m2_dcache_wbd_sel_i[0]
port 100 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 m2_dcache_wbd_sel_i[1]
port 101 nsew signal input
rlabel metal2 s 117870 29200 117926 30000 6 m2_dcache_wbd_sel_i[2]
port 102 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 m2_dcache_wbd_sel_i[3]
port 103 nsew signal input
rlabel metal3 s 119200 27888 120000 28008 6 m2_dcache_wbd_stb_i
port 104 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 m2_dcache_wbd_we_i
port 105 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 m2_others_wbd_ack_o
port 106 nsew signal output
rlabel metal2 s 48962 29200 49018 30000 6 m2_others_wbd_adr_i[0]
port 107 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 m2_others_wbd_adr_i[10]
port 108 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 m2_others_wbd_adr_i[11]
port 109 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 m2_others_wbd_adr_i[12]
port 110 nsew signal input
rlabel metal3 s 119200 14288 120000 14408 6 m2_others_wbd_adr_i[13]
port 111 nsew signal input
rlabel metal2 s 63774 29200 63830 30000 6 m2_others_wbd_adr_i[14]
port 112 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 m2_others_wbd_adr_i[15]
port 113 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 m2_others_wbd_adr_i[16]
port 114 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 m2_others_wbd_adr_i[17]
port 115 nsew signal input
rlabel metal2 s 30930 29200 30986 30000 6 m2_others_wbd_adr_i[18]
port 116 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 m2_others_wbd_adr_i[19]
port 117 nsew signal input
rlabel metal2 s 12254 29200 12310 30000 6 m2_others_wbd_adr_i[1]
port 118 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 m2_others_wbd_adr_i[20]
port 119 nsew signal input
rlabel metal2 s 36082 29200 36138 30000 6 m2_others_wbd_adr_i[21]
port 120 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 m2_others_wbd_adr_i[22]
port 121 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 m2_others_wbd_adr_i[23]
port 122 nsew signal input
rlabel metal3 s 119200 6128 120000 6248 6 m2_others_wbd_adr_i[24]
port 123 nsew signal input
rlabel metal2 s 83094 29200 83150 30000 6 m2_others_wbd_adr_i[25]
port 124 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 m2_others_wbd_adr_i[26]
port 125 nsew signal input
rlabel metal2 s 17406 29200 17462 30000 6 m2_others_wbd_adr_i[27]
port 126 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 m2_others_wbd_adr_i[28]
port 127 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 m2_others_wbd_adr_i[29]
port 128 nsew signal input
rlabel metal2 s 31574 29200 31630 30000 6 m2_others_wbd_adr_i[2]
port 129 nsew signal input
rlabel metal2 s 64418 29200 64474 30000 6 m2_others_wbd_adr_i[30]
port 130 nsew signal input
rlabel metal2 s 88246 29200 88302 30000 6 m2_others_wbd_adr_i[31]
port 131 nsew signal input
rlabel metal2 s 52182 29200 52238 30000 6 m2_others_wbd_adr_i[3]
port 132 nsew signal input
rlabel metal3 s 119200 13608 120000 13728 6 m2_others_wbd_adr_i[4]
port 133 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 m2_others_wbd_adr_i[5]
port 134 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 m2_others_wbd_adr_i[6]
port 135 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 m2_others_wbd_adr_i[7]
port 136 nsew signal input
rlabel metal2 s 91466 29200 91522 30000 6 m2_others_wbd_adr_i[8]
port 137 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 m2_others_wbd_adr_i[9]
port 138 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 m2_others_wbd_cyc_i
port 139 nsew signal input
rlabel metal2 s 118514 29200 118570 30000 6 m2_others_wbd_dat_i[0]
port 140 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 m2_others_wbd_dat_i[10]
port 141 nsew signal input
rlabel metal2 s 76010 29200 76066 30000 6 m2_others_wbd_dat_i[11]
port 142 nsew signal input
rlabel metal3 s 119200 29248 120000 29368 6 m2_others_wbd_dat_i[12]
port 143 nsew signal input
rlabel metal2 s 119802 29200 119858 30000 6 m2_others_wbd_dat_i[13]
port 144 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 m2_others_wbd_dat_i[14]
port 145 nsew signal input
rlabel metal2 s 89534 29200 89590 30000 6 m2_others_wbd_dat_i[15]
port 146 nsew signal input
rlabel metal2 s 74078 29200 74134 30000 6 m2_others_wbd_dat_i[16]
port 147 nsew signal input
rlabel metal2 s 7102 29200 7158 30000 6 m2_others_wbd_dat_i[17]
port 148 nsew signal input
rlabel metal3 s 119200 8 120000 128 6 m2_others_wbd_dat_i[18]
port 149 nsew signal input
rlabel metal2 s 76654 29200 76710 30000 6 m2_others_wbd_dat_i[19]
port 150 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 m2_others_wbd_dat_i[1]
port 151 nsew signal input
rlabel metal2 s 1306 29200 1362 30000 6 m2_others_wbd_dat_i[20]
port 152 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 m2_others_wbd_dat_i[21]
port 153 nsew signal input
rlabel metal2 s 14186 29200 14242 30000 6 m2_others_wbd_dat_i[22]
port 154 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 m2_others_wbd_dat_i[23]
port 155 nsew signal input
rlabel metal2 s 112074 29200 112130 30000 6 m2_others_wbd_dat_i[24]
port 156 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 m2_others_wbd_dat_i[25]
port 157 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 m2_others_wbd_dat_i[26]
port 158 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 m2_others_wbd_dat_i[27]
port 159 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 m2_others_wbd_dat_i[28]
port 160 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 m2_others_wbd_dat_i[29]
port 161 nsew signal input
rlabel metal2 s 101126 29200 101182 30000 6 m2_others_wbd_dat_i[2]
port 162 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 m2_others_wbd_dat_i[30]
port 163 nsew signal input
rlabel metal2 s 21914 29200 21970 30000 6 m2_others_wbd_dat_i[31]
port 164 nsew signal input
rlabel metal2 s 98550 29200 98606 30000 6 m2_others_wbd_dat_i[3]
port 165 nsew signal input
rlabel metal3 s 119200 18368 120000 18488 6 m2_others_wbd_dat_i[4]
port 166 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 m2_others_wbd_dat_i[5]
port 167 nsew signal input
rlabel metal2 s 48318 29200 48374 30000 6 m2_others_wbd_dat_i[6]
port 168 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 m2_others_wbd_dat_i[7]
port 169 nsew signal input
rlabel metal2 s 18050 29200 18106 30000 6 m2_others_wbd_dat_i[8]
port 170 nsew signal input
rlabel metal2 s 25134 29200 25190 30000 6 m2_others_wbd_dat_i[9]
port 171 nsew signal input
rlabel metal2 s 20626 29200 20682 30000 6 m2_others_wbd_dat_o[0]
port 172 nsew signal output
rlabel metal3 s 119200 1368 120000 1488 6 m2_others_wbd_dat_o[10]
port 173 nsew signal output
rlabel metal3 s 119200 4768 120000 4888 6 m2_others_wbd_dat_o[11]
port 174 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 m2_others_wbd_dat_o[12]
port 175 nsew signal output
rlabel metal2 s 55402 29200 55458 30000 6 m2_others_wbd_dat_o[13]
port 176 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 m2_others_wbd_dat_o[14]
port 177 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 m2_others_wbd_dat_o[15]
port 178 nsew signal output
rlabel metal3 s 119200 12928 120000 13048 6 m2_others_wbd_dat_o[16]
port 179 nsew signal output
rlabel metal2 s 97906 29200 97962 30000 6 m2_others_wbd_dat_o[17]
port 180 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 m2_others_wbd_dat_o[18]
port 181 nsew signal output
rlabel metal2 s 92110 29200 92166 30000 6 m2_others_wbd_dat_o[19]
port 182 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 m2_others_wbd_dat_o[1]
port 183 nsew signal output
rlabel metal2 s 56690 29200 56746 30000 6 m2_others_wbd_dat_o[20]
port 184 nsew signal output
rlabel metal3 s 119200 9528 120000 9648 6 m2_others_wbd_dat_o[21]
port 185 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 m2_others_wbd_dat_o[22]
port 186 nsew signal output
rlabel metal2 s 100482 29200 100538 30000 6 m2_others_wbd_dat_o[23]
port 187 nsew signal output
rlabel metal2 s 4526 29200 4582 30000 6 m2_others_wbd_dat_o[24]
port 188 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 m2_others_wbd_dat_o[25]
port 189 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 m2_others_wbd_dat_o[26]
port 190 nsew signal output
rlabel metal3 s 119200 20408 120000 20528 6 m2_others_wbd_dat_o[27]
port 191 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 m2_others_wbd_dat_o[28]
port 192 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 m2_others_wbd_dat_o[29]
port 193 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 m2_others_wbd_dat_o[2]
port 194 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 m2_others_wbd_dat_o[30]
port 195 nsew signal output
rlabel metal2 s 29642 29200 29698 30000 6 m2_others_wbd_dat_o[31]
port 196 nsew signal output
rlabel metal2 s 50894 29200 50950 30000 6 m2_others_wbd_dat_o[3]
port 197 nsew signal output
rlabel metal2 s 94042 29200 94098 30000 6 m2_others_wbd_dat_o[4]
port 198 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 m2_others_wbd_dat_o[5]
port 199 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 m2_others_wbd_dat_o[6]
port 200 nsew signal output
rlabel metal2 s 117226 29200 117282 30000 6 m2_others_wbd_dat_o[7]
port 201 nsew signal output
rlabel metal2 s 77298 29200 77354 30000 6 m2_others_wbd_dat_o[8]
port 202 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 m2_others_wbd_dat_o[9]
port 203 nsew signal output
rlabel metal2 s 3238 29200 3294 30000 6 m2_others_wbd_sel_i[0]
port 204 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 m2_others_wbd_sel_i[1]
port 205 nsew signal input
rlabel metal2 s 110786 29200 110842 30000 6 m2_others_wbd_sel_i[2]
port 206 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 m2_others_wbd_sel_i[3]
port 207 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 m2_others_wbd_stb_i
port 208 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 m2_others_wbd_we_i
port 209 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 m2_wbd_ack_i
port 210 nsew signal input
rlabel metal2 s 61842 29200 61898 30000 6 m2_wbd_adr_o[0]
port 211 nsew signal output
rlabel metal2 s 58622 29200 58678 30000 6 m2_wbd_adr_o[10]
port 212 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 m2_wbd_adr_o[11]
port 213 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 m2_wbd_adr_o[12]
port 214 nsew signal output
rlabel metal2 s 87602 29200 87658 30000 6 m2_wbd_adr_o[13]
port 215 nsew signal output
rlabel metal3 s 119200 24488 120000 24608 6 m2_wbd_adr_o[14]
port 216 nsew signal output
rlabel metal2 s 61198 29200 61254 30000 6 m2_wbd_adr_o[15]
port 217 nsew signal output
rlabel metal2 s 83738 29200 83794 30000 6 m2_wbd_adr_o[16]
port 218 nsew signal output
rlabel metal2 s 90178 29200 90234 30000 6 m2_wbd_adr_o[17]
port 219 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 m2_wbd_adr_o[18]
port 220 nsew signal output
rlabel metal2 s 79230 29200 79286 30000 6 m2_wbd_adr_o[19]
port 221 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 m2_wbd_adr_o[1]
port 222 nsew signal output
rlabel metal2 s 111430 29200 111486 30000 6 m2_wbd_adr_o[20]
port 223 nsew signal output
rlabel metal2 s 96618 29200 96674 30000 6 m2_wbd_adr_o[21]
port 224 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 m2_wbd_adr_o[22]
port 225 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 m2_wbd_adr_o[23]
port 226 nsew signal output
rlabel metal2 s 50250 29200 50306 30000 6 m2_wbd_adr_o[24]
port 227 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 m2_wbd_adr_o[25]
port 228 nsew signal output
rlabel metal2 s 24490 29200 24546 30000 6 m2_wbd_adr_o[26]
port 229 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 m2_wbd_adr_o[27]
port 230 nsew signal output
rlabel metal2 s 47030 29200 47086 30000 6 m2_wbd_adr_o[28]
port 231 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 m2_wbd_adr_o[29]
port 232 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 m2_wbd_adr_o[2]
port 233 nsew signal output
rlabel metal2 s 107566 29200 107622 30000 6 m2_wbd_adr_o[30]
port 234 nsew signal output
rlabel metal3 s 119200 22448 120000 22568 6 m2_wbd_adr_o[31]
port 235 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 m2_wbd_adr_o[3]
port 236 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 m2_wbd_adr_o[4]
port 237 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 m2_wbd_adr_o[5]
port 238 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 m2_wbd_adr_o[6]
port 239 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 m2_wbd_adr_o[7]
port 240 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 m2_wbd_adr_o[8]
port 241 nsew signal output
rlabel metal2 s 85026 29200 85082 30000 6 m2_wbd_adr_o[9]
port 242 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 m2_wbd_bl_o[0]
port 243 nsew signal output
rlabel metal3 s 119200 15648 120000 15768 6 m2_wbd_bl_o[1]
port 244 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 m2_wbd_bl_o[2]
port 245 nsew signal output
rlabel metal2 s 115294 29200 115350 30000 6 m2_wbd_bl_o[3]
port 246 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 m2_wbd_bl_o[4]
port 247 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 m2_wbd_bl_o[5]
port 248 nsew signal output
rlabel metal2 s 113362 29200 113418 30000 6 m2_wbd_bl_o[6]
port 249 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 m2_wbd_bl_o[7]
port 250 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 m2_wbd_bl_o[8]
port 251 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 m2_wbd_bl_o[9]
port 252 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 m2_wbd_bry_o
port 253 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 m2_wbd_cyc_o
port 254 nsew signal output
rlabel metal2 s 80518 29200 80574 30000 6 m2_wbd_dat_i[0]
port 255 nsew signal input
rlabel metal3 s 119200 11568 120000 11688 6 m2_wbd_dat_i[10]
port 256 nsew signal input
rlabel metal2 s 41878 29200 41934 30000 6 m2_wbd_dat_i[11]
port 257 nsew signal input
rlabel metal2 s 46386 29200 46442 30000 6 m2_wbd_dat_i[12]
port 258 nsew signal input
rlabel metal2 s 44454 29200 44510 30000 6 m2_wbd_dat_i[13]
port 259 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 m2_wbd_dat_i[14]
port 260 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 m2_wbd_dat_i[15]
port 261 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 m2_wbd_dat_i[16]
port 262 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 m2_wbd_dat_i[17]
port 263 nsew signal input
rlabel metal2 s 104990 29200 105046 30000 6 m2_wbd_dat_i[18]
port 264 nsew signal input
rlabel metal3 s 119200 27208 120000 27328 6 m2_wbd_dat_i[19]
port 265 nsew signal input
rlabel metal2 s 59910 29200 59966 30000 6 m2_wbd_dat_i[1]
port 266 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 m2_wbd_dat_i[20]
port 267 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 m2_wbd_dat_i[21]
port 268 nsew signal input
rlabel metal3 s 119200 26528 120000 26648 6 m2_wbd_dat_i[22]
port 269 nsew signal input
rlabel metal2 s 26422 29200 26478 30000 6 m2_wbd_dat_i[23]
port 270 nsew signal input
rlabel metal3 s 119200 6808 120000 6928 6 m2_wbd_dat_i[24]
port 271 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 m2_wbd_dat_i[25]
port 272 nsew signal input
rlabel metal2 s 18 29200 74 30000 6 m2_wbd_dat_i[26]
port 273 nsew signal input
rlabel metal2 s 114006 29200 114062 30000 6 m2_wbd_dat_i[27]
port 274 nsew signal input
rlabel metal2 s 72146 29200 72202 30000 6 m2_wbd_dat_i[28]
port 275 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 m2_wbd_dat_i[29]
port 276 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 m2_wbd_dat_i[2]
port 277 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 m2_wbd_dat_i[30]
port 278 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 m2_wbd_dat_i[31]
port 279 nsew signal input
rlabel metal2 s 19982 29200 20038 30000 6 m2_wbd_dat_i[3]
port 280 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 m2_wbd_dat_i[4]
port 281 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 m2_wbd_dat_i[5]
port 282 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 m2_wbd_dat_i[6]
port 283 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 m2_wbd_dat_i[7]
port 284 nsew signal input
rlabel metal2 s 109498 29200 109554 30000 6 m2_wbd_dat_i[8]
port 285 nsew signal input
rlabel metal3 s 119200 17688 120000 17808 6 m2_wbd_dat_i[9]
port 286 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 m2_wbd_dat_o[0]
port 287 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 m2_wbd_dat_o[10]
port 288 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 m2_wbd_dat_o[11]
port 289 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 m2_wbd_dat_o[12]
port 290 nsew signal output
rlabel metal3 s 119200 19728 120000 19848 6 m2_wbd_dat_o[13]
port 291 nsew signal output
rlabel metal2 s 105634 29200 105690 30000 6 m2_wbd_dat_o[14]
port 292 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 m2_wbd_dat_o[15]
port 293 nsew signal output
rlabel metal2 s 103058 29200 103114 30000 6 m2_wbd_dat_o[16]
port 294 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 m2_wbd_dat_o[17]
port 295 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 m2_wbd_dat_o[18]
port 296 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 m2_wbd_dat_o[19]
port 297 nsew signal output
rlabel metal2 s 18 0 74 800 6 m2_wbd_dat_o[1]
port 298 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 m2_wbd_dat_o[20]
port 299 nsew signal output
rlabel metal2 s 11610 29200 11666 30000 6 m2_wbd_dat_o[21]
port 300 nsew signal output
rlabel metal2 s 39946 29200 40002 30000 6 m2_wbd_dat_o[22]
port 301 nsew signal output
rlabel metal2 s 69570 29200 69626 30000 6 m2_wbd_dat_o[23]
port 302 nsew signal output
rlabel metal2 s 662 29200 718 30000 6 m2_wbd_dat_o[24]
port 303 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 m2_wbd_dat_o[25]
port 304 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 m2_wbd_dat_o[26]
port 305 nsew signal output
rlabel metal2 s 86958 29200 87014 30000 6 m2_wbd_dat_o[27]
port 306 nsew signal output
rlabel metal2 s 70214 29200 70270 30000 6 m2_wbd_dat_o[28]
port 307 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 m2_wbd_dat_o[29]
port 308 nsew signal output
rlabel metal2 s 99838 29200 99894 30000 6 m2_wbd_dat_o[2]
port 309 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 m2_wbd_dat_o[30]
port 310 nsew signal output
rlabel metal2 s 22558 29200 22614 30000 6 m2_wbd_dat_o[31]
port 311 nsew signal output
rlabel metal3 s 119200 10888 120000 11008 6 m2_wbd_dat_o[3]
port 312 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 m2_wbd_dat_o[4]
port 313 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 m2_wbd_dat_o[5]
port 314 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 m2_wbd_dat_o[6]
port 315 nsew signal output
rlabel metal3 s 119200 8168 120000 8288 6 m2_wbd_dat_o[7]
port 316 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 m2_wbd_dat_o[8]
port 317 nsew signal output
rlabel metal2 s 95974 29200 96030 30000 6 m2_wbd_dat_o[9]
port 318 nsew signal output
rlabel metal2 s 94686 29200 94742 30000 6 m2_wbd_sel_o[0]
port 319 nsew signal output
rlabel metal2 s 41234 29200 41290 30000 6 m2_wbd_sel_o[1]
port 320 nsew signal output
rlabel metal2 s 54758 29200 54814 30000 6 m2_wbd_sel_o[2]
port 321 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 m2_wbd_sel_o[3]
port 322 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 m2_wbd_stb_o
port 323 nsew signal output
rlabel metal2 s 32862 29200 32918 30000 6 m2_wbd_we_o
port 324 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 reset
port 325 nsew signal input
rlabel metal4 s 15668 2128 15988 27792 6 vccd1
port 326 nsew power bidirectional
rlabel metal4 s 45116 2128 45436 27792 6 vccd1
port 326 nsew power bidirectional
rlabel metal4 s 74564 2128 74884 27792 6 vccd1
port 326 nsew power bidirectional
rlabel metal4 s 104012 2128 104332 27792 6 vccd1
port 326 nsew power bidirectional
rlabel metal4 s 30392 2128 30712 27792 6 vssd1
port 327 nsew ground bidirectional
rlabel metal4 s 59840 2128 60160 27792 6 vssd1
port 327 nsew ground bidirectional
rlabel metal4 s 89288 2128 89608 27792 6 vssd1
port 327 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2182396
string GDS_FILE /root/hellochip/openlane/arbitor/runs/22_09_12_23_50/results/signoff/bus_arbiter.magic.gds
string GDS_START 149640
<< end >>

