VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1950.000 BY 1950.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1009.840 1950.000 1010.440 ;
    END
  END clk
  PIN dcache_data_chip_en_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 605.240 1950.000 605.840 ;
    END
  END dcache_data_chip_en_1
  PIN dcache_data_chip_en_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END dcache_data_chip_en_2
  PIN dcache_data_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1883.640 4.000 1884.240 ;
    END
  END dcache_data_in_1[0]
  PIN dcache_data_in_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1111.840 1950.000 1112.440 ;
    END
  END dcache_data_in_1[10]
  PIN dcache_data_in_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1946.000 721.650 1950.000 ;
    END
  END dcache_data_in_1[11]
  PIN dcache_data_in_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END dcache_data_in_1[12]
  PIN dcache_data_in_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 1946.000 618.610 1950.000 ;
    END
  END dcache_data_in_1[13]
  PIN dcache_data_in_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 1946.000 1111.270 1950.000 ;
    END
  END dcache_data_in_1[14]
  PIN dcache_data_in_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END dcache_data_in_1[15]
  PIN dcache_data_in_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 0.000 1336.670 4.000 ;
    END
  END dcache_data_in_1[16]
  PIN dcache_data_in_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END dcache_data_in_1[17]
  PIN dcache_data_in_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1946.000 235.430 1950.000 ;
    END
  END dcache_data_in_1[18]
  PIN dcache_data_in_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 1946.000 972.810 1950.000 ;
    END
  END dcache_data_in_1[19]
  PIN dcache_data_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END dcache_data_in_1[1]
  PIN dcache_data_in_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.450 1946.000 1893.730 1950.000 ;
    END
  END dcache_data_in_1[20]
  PIN dcache_data_in_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END dcache_data_in_1[21]
  PIN dcache_data_in_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 1946.000 947.050 1950.000 ;
    END
  END dcache_data_in_1[22]
  PIN dcache_data_in_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 1946.000 486.590 1950.000 ;
    END
  END dcache_data_in_1[23]
  PIN dcache_data_in_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END dcache_data_in_1[24]
  PIN dcache_data_in_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1781.640 4.000 1782.240 ;
    END
  END dcache_data_in_1[25]
  PIN dcache_data_in_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1946.000 1072.630 1950.000 ;
    END
  END dcache_data_in_1[26]
  PIN dcache_data_in_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END dcache_data_in_1[27]
  PIN dcache_data_in_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END dcache_data_in_1[28]
  PIN dcache_data_in_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END dcache_data_in_1[29]
  PIN dcache_data_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 996.240 1950.000 996.840 ;
    END
  END dcache_data_in_1[2]
  PIN dcache_data_in_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.310 0.000 1935.590 4.000 ;
    END
  END dcache_data_in_1[30]
  PIN dcache_data_in_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END dcache_data_in_1[31]
  PIN dcache_data_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END dcache_data_in_1[3]
  PIN dcache_data_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1577.640 4.000 1578.240 ;
    END
  END dcache_data_in_1[4]
  PIN dcache_data_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END dcache_data_in_1[5]
  PIN dcache_data_in_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 0.000 1233.630 4.000 ;
    END
  END dcache_data_in_1[6]
  PIN dcache_data_in_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1390.640 1950.000 1391.240 ;
    END
  END dcache_data_in_1[7]
  PIN dcache_data_in_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END dcache_data_in_1[8]
  PIN dcache_data_in_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 1946.000 554.210 1950.000 ;
    END
  END dcache_data_in_1[9]
  PIN dcache_data_in_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1220.640 1950.000 1221.240 ;
    END
  END dcache_data_in_2[0]
  PIN dcache_data_in_2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END dcache_data_in_2[10]
  PIN dcache_data_in_2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 652.840 1950.000 653.440 ;
    END
  END dcache_data_in_2[11]
  PIN dcache_data_in_2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 1946.000 1816.450 1950.000 ;
    END
  END dcache_data_in_2[12]
  PIN dcache_data_in_2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END dcache_data_in_2[13]
  PIN dcache_data_in_2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.040 4.000 1445.640 ;
    END
  END dcache_data_in_2[14]
  PIN dcache_data_in_2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 1946.000 760.290 1950.000 ;
    END
  END dcache_data_in_2[15]
  PIN dcache_data_in_2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 1946.000 1362.430 1950.000 ;
    END
  END dcache_data_in_2[16]
  PIN dcache_data_in_2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 516.840 1950.000 517.440 ;
    END
  END dcache_data_in_2[17]
  PIN dcache_data_in_2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1761.240 4.000 1761.840 ;
    END
  END dcache_data_in_2[18]
  PIN dcache_data_in_2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 153.040 1950.000 153.640 ;
    END
  END dcache_data_in_2[19]
  PIN dcache_data_in_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END dcache_data_in_2[1]
  PIN dcache_data_in_2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1618.440 1950.000 1619.040 ;
    END
  END dcache_data_in_2[20]
  PIN dcache_data_in_2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END dcache_data_in_2[21]
  PIN dcache_data_in_2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 1946.000 441.510 1950.000 ;
    END
  END dcache_data_in_2[22]
  PIN dcache_data_in_2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 476.040 1950.000 476.640 ;
    END
  END dcache_data_in_2[23]
  PIN dcache_data_in_2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1570.840 1950.000 1571.440 ;
    END
  END dcache_data_in_2[24]
  PIN dcache_data_in_2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 1946.000 683.010 1950.000 ;
    END
  END dcache_data_in_2[25]
  PIN dcache_data_in_2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END dcache_data_in_2[26]
  PIN dcache_data_in_2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END dcache_data_in_2[27]
  PIN dcache_data_in_2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 329.840 1950.000 330.440 ;
    END
  END dcache_data_in_2[28]
  PIN dcache_data_in_2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 302.640 1950.000 303.240 ;
    END
  END dcache_data_in_2[29]
  PIN dcache_data_in_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 1946.000 702.330 1950.000 ;
    END
  END dcache_data_in_2[2]
  PIN dcache_data_in_2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1118.640 4.000 1119.240 ;
    END
  END dcache_data_in_2[30]
  PIN dcache_data_in_2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 1946.000 1310.910 1950.000 ;
    END
  END dcache_data_in_2[31]
  PIN dcache_data_in_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 1946.000 1143.470 1950.000 ;
    END
  END dcache_data_in_2[3]
  PIN dcache_data_in_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1700.040 4.000 1700.640 ;
    END
  END dcache_data_in_2[4]
  PIN dcache_data_in_2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 1946.000 1452.590 1950.000 ;
    END
  END dcache_data_in_2[5]
  PIN dcache_data_in_2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END dcache_data_in_2[6]
  PIN dcache_data_in_2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1502.840 4.000 1503.440 ;
    END
  END dcache_data_in_2[7]
  PIN dcache_data_in_2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 1946.000 1033.990 1950.000 ;
    END
  END dcache_data_in_2[8]
  PIN dcache_data_in_2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END dcache_data_in_2[9]
  PIN dcache_data_index_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END dcache_data_index_1[0]
  PIN dcache_data_index_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1754.440 1950.000 1755.040 ;
    END
  END dcache_data_index_1[1]
  PIN dcache_data_index_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.690 0.000 1867.970 4.000 ;
    END
  END dcache_data_index_1[2]
  PIN dcache_data_index_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END dcache_data_index_1[3]
  PIN dcache_data_index_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END dcache_data_index_1[4]
  PIN dcache_data_index_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1904.040 1950.000 1904.640 ;
    END
  END dcache_data_index_1[5]
  PIN dcache_data_index_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 1946.000 805.370 1950.000 ;
    END
  END dcache_data_index_1[6]
  PIN dcache_data_index_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 1946.000 241.870 1950.000 ;
    END
  END dcache_data_index_1[7]
  PIN dcache_data_index_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1946.000 747.410 1950.000 ;
    END
  END dcache_data_index_2[0]
  PIN dcache_data_index_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END dcache_data_index_2[1]
  PIN dcache_data_index_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 584.840 1950.000 585.440 ;
    END
  END dcache_data_index_2[2]
  PIN dcache_data_index_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END dcache_data_index_2[3]
  PIN dcache_data_index_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 1946.000 1545.970 1950.000 ;
    END
  END dcache_data_index_2[4]
  PIN dcache_data_index_2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END dcache_data_index_2[5]
  PIN dcache_data_index_2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 1946.000 357.790 1950.000 ;
    END
  END dcache_data_index_2[6]
  PIN dcache_data_index_2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1424.640 1950.000 1425.240 ;
    END
  END dcache_data_index_2[7]
  PIN dcache_data_out_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 1946.000 663.690 1950.000 ;
    END
  END dcache_data_out_1[0]
  PIN dcache_data_out_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 1946.000 985.690 1950.000 ;
    END
  END dcache_data_out_1[10]
  PIN dcache_data_out_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1557.240 4.000 1557.840 ;
    END
  END dcache_data_out_1[11]
  PIN dcache_data_out_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 0.000 1642.570 4.000 ;
    END
  END dcache_data_out_1[12]
  PIN dcache_data_out_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1679.640 4.000 1680.240 ;
    END
  END dcache_data_out_1[13]
  PIN dcache_data_out_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 0.000 1091.950 4.000 ;
    END
  END dcache_data_out_1[14]
  PIN dcache_data_out_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END dcache_data_out_1[15]
  PIN dcache_data_out_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1557.240 1950.000 1557.840 ;
    END
  END dcache_data_out_1[16]
  PIN dcache_data_out_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END dcache_data_out_1[17]
  PIN dcache_data_out_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END dcache_data_out_1[18]
  PIN dcache_data_out_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 1946.000 196.790 1950.000 ;
    END
  END dcache_data_out_1[19]
  PIN dcache_data_out_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END dcache_data_out_1[1]
  PIN dcache_data_out_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1598.040 1950.000 1598.640 ;
    END
  END dcache_data_out_1[20]
  PIN dcache_data_out_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 768.440 1950.000 769.040 ;
    END
  END dcache_data_out_1[21]
  PIN dcache_data_out_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END dcache_data_out_1[22]
  PIN dcache_data_out_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 0.000 1436.490 4.000 ;
    END
  END dcache_data_out_1[23]
  PIN dcache_data_out_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 0.000 1661.890 4.000 ;
    END
  END dcache_data_out_1[24]
  PIN dcache_data_out_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END dcache_data_out_1[25]
  PIN dcache_data_out_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 829.640 1950.000 830.240 ;
    END
  END dcache_data_out_1[26]
  PIN dcache_data_out_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END dcache_data_out_1[27]
  PIN dcache_data_out_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 1946.000 1558.850 1950.000 ;
    END
  END dcache_data_out_1[28]
  PIN dcache_data_out_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 1946.000 1104.830 1950.000 ;
    END
  END dcache_data_out_1[29]
  PIN dcache_data_out_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1645.640 1950.000 1646.240 ;
    END
  END dcache_data_out_1[2]
  PIN dcache_data_out_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END dcache_data_out_1[30]
  PIN dcache_data_out_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 673.240 1950.000 673.840 ;
    END
  END dcache_data_out_1[31]
  PIN dcache_data_out_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1946.000 0.370 1950.000 ;
    END
  END dcache_data_out_1[3]
  PIN dcache_data_out_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1740.840 1950.000 1741.440 ;
    END
  END dcache_data_out_1[4]
  PIN dcache_data_out_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END dcache_data_out_1[5]
  PIN dcache_data_out_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END dcache_data_out_1[6]
  PIN dcache_data_out_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END dcache_data_out_1[7]
  PIN dcache_data_out_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.750 0.000 1942.030 4.000 ;
    END
  END dcache_data_out_1[8]
  PIN dcache_data_out_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END dcache_data_out_1[9]
  PIN dcache_data_out_2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END dcache_data_out_2[0]
  PIN dcache_data_out_2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 384.240 1950.000 384.840 ;
    END
  END dcache_data_out_2[10]
  PIN dcache_data_out_2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END dcache_data_out_2[11]
  PIN dcache_data_out_2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1659.240 1950.000 1659.840 ;
    END
  END dcache_data_out_2[12]
  PIN dcache_data_out_2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1315.840 1950.000 1316.440 ;
    END
  END dcache_data_out_2[13]
  PIN dcache_data_out_2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 1946.000 325.590 1950.000 ;
    END
  END dcache_data_out_2[14]
  PIN dcache_data_out_2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 1946.000 402.870 1950.000 ;
    END
  END dcache_data_out_2[15]
  PIN dcache_data_out_2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 537.240 1950.000 537.840 ;
    END
  END dcache_data_out_2[16]
  PIN dcache_data_out_2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END dcache_data_out_2[17]
  PIN dcache_data_out_2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1166.240 1950.000 1166.840 ;
    END
  END dcache_data_out_2[18]
  PIN dcache_data_out_2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 1946.000 1214.310 1950.000 ;
    END
  END dcache_data_out_2[19]
  PIN dcache_data_out_2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END dcache_data_out_2[1]
  PIN dcache_data_out_2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 1946.000 499.470 1950.000 ;
    END
  END dcache_data_out_2[20]
  PIN dcache_data_out_2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.370 1946.000 1848.650 1950.000 ;
    END
  END dcache_data_out_2[21]
  PIN dcache_data_out_2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 1946.000 1085.510 1950.000 ;
    END
  END dcache_data_out_2[22]
  PIN dcache_data_out_2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END dcache_data_out_2[23]
  PIN dcache_data_out_2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 1946.000 1835.770 1950.000 ;
    END
  END dcache_data_out_2[24]
  PIN dcache_data_out_2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END dcache_data_out_2[25]
  PIN dcache_data_out_2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END dcache_data_out_2[26]
  PIN dcache_data_out_2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 445.440 1950.000 446.040 ;
    END
  END dcache_data_out_2[27]
  PIN dcache_data_out_2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END dcache_data_out_2[28]
  PIN dcache_data_out_2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END dcache_data_out_2[29]
  PIN dcache_data_out_2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 125.840 1950.000 126.440 ;
    END
  END dcache_data_out_2[2]
  PIN dcache_data_out_2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 1946.000 493.030 1950.000 ;
    END
  END dcache_data_out_2[30]
  PIN dcache_data_out_2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 1946.000 45.450 1950.000 ;
    END
  END dcache_data_out_2[31]
  PIN dcache_data_out_2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END dcache_data_out_2[3]
  PIN dcache_data_out_2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END dcache_data_out_2[4]
  PIN dcache_data_out_2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END dcache_data_out_2[5]
  PIN dcache_data_out_2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 1946.000 377.110 1950.000 ;
    END
  END dcache_data_out_2[6]
  PIN dcache_data_out_2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1727.240 1950.000 1727.840 ;
    END
  END dcache_data_out_2[7]
  PIN dcache_data_out_2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END dcache_data_out_2[8]
  PIN dcache_data_out_2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1788.440 4.000 1789.040 ;
    END
  END dcache_data_out_2[9]
  PIN dcache_data_write_en_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1336.240 1950.000 1336.840 ;
    END
  END dcache_data_write_en_1
  PIN dcache_data_write_en_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1946.000 364.230 1950.000 ;
    END
  END dcache_data_write_en_2
  PIN dcache_tag_chip_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 0.000 1713.410 4.000 ;
    END
  END dcache_tag_chip_en
  PIN dcache_tag_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 234.640 1950.000 235.240 ;
    END
  END dcache_tag_data_in[0]
  PIN dcache_tag_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 1946.000 132.390 1950.000 ;
    END
  END dcache_tag_data_in[10]
  PIN dcache_tag_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 0.000 1797.130 4.000 ;
    END
  END dcache_tag_data_in[11]
  PIN dcache_tag_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 618.840 1950.000 619.440 ;
    END
  END dcache_tag_data_in[12]
  PIN dcache_tag_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 0.000 1462.250 4.000 ;
    END
  END dcache_tag_data_in[13]
  PIN dcache_tag_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 1946.000 753.850 1950.000 ;
    END
  END dcache_tag_data_in[14]
  PIN dcache_tag_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1125.440 4.000 1126.040 ;
    END
  END dcache_tag_data_in[15]
  PIN dcache_tag_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END dcache_tag_data_in[16]
  PIN dcache_tag_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1159.440 1950.000 1160.040 ;
    END
  END dcache_tag_data_in[17]
  PIN dcache_tag_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1247.840 1950.000 1248.440 ;
    END
  END dcache_tag_data_in[18]
  PIN dcache_tag_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 1946.000 547.770 1950.000 ;
    END
  END dcache_tag_data_in[19]
  PIN dcache_tag_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END dcache_tag_data_in[1]
  PIN dcache_tag_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1946.000 528.450 1950.000 ;
    END
  END dcache_tag_data_in[20]
  PIN dcache_tag_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.870 0.000 1929.150 4.000 ;
    END
  END dcache_tag_data_in[21]
  PIN dcache_tag_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1530.040 1950.000 1530.640 ;
    END
  END dcache_tag_data_in[22]
  PIN dcache_tag_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 1946.000 1603.930 1950.000 ;
    END
  END dcache_tag_data_in[23]
  PIN dcache_tag_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1740.840 4.000 1741.440 ;
    END
  END dcache_tag_data_in[24]
  PIN dcache_tag_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 51.040 1950.000 51.640 ;
    END
  END dcache_tag_data_in[25]
  PIN dcache_tag_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END dcache_tag_data_in[26]
  PIN dcache_tag_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 0.000 1674.770 4.000 ;
    END
  END dcache_tag_data_in[27]
  PIN dcache_tag_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1241.040 1950.000 1241.640 ;
    END
  END dcache_tag_data_in[28]
  PIN dcache_tag_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END dcache_tag_data_in[29]
  PIN dcache_tag_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1693.240 4.000 1693.840 ;
    END
  END dcache_tag_data_in[2]
  PIN dcache_tag_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1604.840 1950.000 1605.440 ;
    END
  END dcache_tag_data_in[30]
  PIN dcache_tag_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 1946.000 876.210 1950.000 ;
    END
  END dcache_tag_data_in[31]
  PIN dcache_tag_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END dcache_tag_data_in[3]
  PIN dcache_tag_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END dcache_tag_data_in[4]
  PIN dcache_tag_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END dcache_tag_data_in[5]
  PIN dcache_tag_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.240 4.000 1234.840 ;
    END
  END dcache_tag_data_in[6]
  PIN dcache_tag_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.040 4.000 1207.640 ;
    END
  END dcache_tag_data_in[7]
  PIN dcache_tag_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 1946.000 1265.830 1950.000 ;
    END
  END dcache_tag_data_in[8]
  PIN dcache_tag_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1720.440 4.000 1721.040 ;
    END
  END dcache_tag_data_in[9]
  PIN dcache_tag_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 1946.000 586.410 1950.000 ;
    END
  END dcache_tag_index[0]
  PIN dcache_tag_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END dcache_tag_index[1]
  PIN dcache_tag_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1693.240 1950.000 1693.840 ;
    END
  END dcache_tag_index[2]
  PIN dcache_tag_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1611.640 1950.000 1612.240 ;
    END
  END dcache_tag_index[3]
  PIN dcache_tag_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1734.040 4.000 1734.640 ;
    END
  END dcache_tag_index[4]
  PIN dcache_tag_index[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1706.840 4.000 1707.440 ;
    END
  END dcache_tag_index[5]
  PIN dcache_tag_index[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END dcache_tag_index[6]
  PIN dcache_tag_index[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END dcache_tag_index[7]
  PIN dcache_tag_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END dcache_tag_out[0]
  PIN dcache_tag_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END dcache_tag_out[10]
  PIN dcache_tag_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 1946.000 676.570 1950.000 ;
    END
  END dcache_tag_out[11]
  PIN dcache_tag_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 391.040 1950.000 391.640 ;
    END
  END dcache_tag_out[12]
  PIN dcache_tag_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 1946.000 1381.750 1950.000 ;
    END
  END dcache_tag_out[13]
  PIN dcache_tag_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 1946.000 1649.010 1950.000 ;
    END
  END dcache_tag_out[14]
  PIN dcache_tag_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 30.640 1950.000 31.240 ;
    END
  END dcache_tag_out[15]
  PIN dcache_tag_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 1946.000 998.570 1950.000 ;
    END
  END dcache_tag_out[16]
  PIN dcache_tag_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 1946.000 254.750 1950.000 ;
    END
  END dcache_tag_out[17]
  PIN dcache_tag_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1492.640 4.000 1493.240 ;
    END
  END dcache_tag_out[18]
  PIN dcache_tag_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1336.240 4.000 1336.840 ;
    END
  END dcache_tag_out[19]
  PIN dcache_tag_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1910.840 4.000 1911.440 ;
    END
  END dcache_tag_out[1]
  PIN dcache_tag_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 1946.000 306.270 1950.000 ;
    END
  END dcache_tag_out[20]
  PIN dcache_tag_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 0.000 1603.930 4.000 ;
    END
  END dcache_tag_out[21]
  PIN dcache_tag_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END dcache_tag_out[22]
  PIN dcache_tag_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END dcache_tag_out[23]
  PIN dcache_tag_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 510.040 1950.000 510.640 ;
    END
  END dcache_tag_out[24]
  PIN dcache_tag_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1946.000 119.510 1950.000 ;
    END
  END dcache_tag_out[25]
  PIN dcache_tag_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END dcache_tag_out[26]
  PIN dcache_tag_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 1946.000 338.470 1950.000 ;
    END
  END dcache_tag_out[27]
  PIN dcache_tag_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END dcache_tag_out[28]
  PIN dcache_tag_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 1946.000 1175.670 1950.000 ;
    END
  END dcache_tag_out[29]
  PIN dcache_tag_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 0.000 1304.470 4.000 ;
    END
  END dcache_tag_out[2]
  PIN dcache_tag_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1455.240 1950.000 1455.840 ;
    END
  END dcache_tag_out[30]
  PIN dcache_tag_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 0.000 1513.770 4.000 ;
    END
  END dcache_tag_out[31]
  PIN dcache_tag_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END dcache_tag_out[3]
  PIN dcache_tag_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.610 0.000 1822.890 4.000 ;
    END
  END dcache_tag_out[4]
  PIN dcache_tag_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 295.840 1950.000 296.440 ;
    END
  END dcache_tag_out[5]
  PIN dcache_tag_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END dcache_tag_out[6]
  PIN dcache_tag_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END dcache_tag_out[7]
  PIN dcache_tag_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 1946.000 1439.710 1950.000 ;
    END
  END dcache_tag_out[8]
  PIN dcache_tag_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 1946.000 1059.750 1950.000 ;
    END
  END dcache_tag_out[9]
  PIN dcache_tag_write_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1829.240 1950.000 1829.840 ;
    END
  END dcache_tag_write_en
  PIN dcache_write_data_mask_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END dcache_write_data_mask_1[0]
  PIN dcache_write_data_mask_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 1946.000 728.090 1950.000 ;
    END
  END dcache_write_data_mask_1[1]
  PIN dcache_write_data_mask_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END dcache_write_data_mask_1[2]
  PIN dcache_write_data_mask_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1377.040 1950.000 1377.640 ;
    END
  END dcache_write_data_mask_1[3]
  PIN dcache_write_data_mask_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END dcache_write_data_mask_2[0]
  PIN dcache_write_data_mask_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1713.640 4.000 1714.240 ;
    END
  END dcache_write_data_mask_2[1]
  PIN dcache_write_data_mask_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.730 0.000 1810.010 4.000 ;
    END
  END dcache_write_data_mask_2[2]
  PIN dcache_write_data_mask_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END dcache_write_data_mask_2[3]
  PIN dcache_write_tag_mask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1536.840 1950.000 1537.440 ;
    END
  END dcache_write_tag_mask[0]
  PIN dcache_write_tag_mask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END dcache_write_tag_mask[1]
  PIN dcache_write_tag_mask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 1946.000 274.070 1950.000 ;
    END
  END dcache_write_tag_mask[2]
  PIN dcache_write_tag_mask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1071.040 1950.000 1071.640 ;
    END
  END dcache_write_tag_mask[3]
  PIN dram_addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END dram_addr0[0]
  PIN dram_addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 1946.000 1726.290 1950.000 ;
    END
  END dram_addr0[1]
  PIN dram_addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 411.440 1950.000 412.040 ;
    END
  END dram_addr0[2]
  PIN dram_addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 1946.000 1413.950 1950.000 ;
    END
  END dram_addr0[3]
  PIN dram_addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 1946.000 740.970 1950.000 ;
    END
  END dram_addr0[4]
  PIN dram_addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END dram_addr0[5]
  PIN dram_addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END dram_addr0[6]
  PIN dram_addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1186.640 1950.000 1187.240 ;
    END
  END dram_addr0[7]
  PIN dram_clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 1946.000 1571.730 1950.000 ;
    END
  END dram_clk0
  PIN dram_csb0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END dram_csb0
  PIN dram_din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 1946.000 1500.890 1950.000 ;
    END
  END dram_din0[0]
  PIN dram_din0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 0.000 1539.530 4.000 ;
    END
  END dram_din0[10]
  PIN dram_din0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 404.640 1950.000 405.240 ;
    END
  END dram_din0[11]
  PIN dram_din0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1397.440 4.000 1398.040 ;
    END
  END dram_din0[12]
  PIN dram_din0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1883.640 1950.000 1884.240 ;
    END
  END dram_din0[13]
  PIN dram_din0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 816.040 1950.000 816.640 ;
    END
  END dram_din0[14]
  PIN dram_din0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END dram_din0[15]
  PIN dram_din0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END dram_din0[16]
  PIN dram_din0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1890.440 1950.000 1891.040 ;
    END
  END dram_din0[17]
  PIN dram_din0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1431.440 1950.000 1432.040 ;
    END
  END dram_din0[18]
  PIN dram_din0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END dram_din0[19]
  PIN dram_din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END dram_din0[1]
  PIN dram_din0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 962.240 1950.000 962.840 ;
    END
  END dram_din0[20]
  PIN dram_din0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 1946.000 934.170 1950.000 ;
    END
  END dram_din0[21]
  PIN dram_din0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1917.640 4.000 1918.240 ;
    END
  END dram_din0[22]
  PIN dram_din0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END dram_din0[23]
  PIN dram_din0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END dram_din0[24]
  PIN dram_din0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END dram_din0[25]
  PIN dram_din0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END dram_din0[26]
  PIN dram_din0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END dram_din0[27]
  PIN dram_din0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1946.000 480.150 1950.000 ;
    END
  END dram_din0[28]
  PIN dram_din0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 0.000 1401.070 4.000 ;
    END
  END dram_din0[29]
  PIN dram_din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 646.040 1950.000 646.640 ;
    END
  END dram_din0[2]
  PIN dram_din0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 0.000 1855.090 4.000 ;
    END
  END dram_din0[30]
  PIN dram_din0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 105.440 1950.000 106.040 ;
    END
  END dram_din0[31]
  PIN dram_din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END dram_din0[3]
  PIN dram_din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END dram_din0[4]
  PIN dram_din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END dram_din0[5]
  PIN dram_din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1288.640 4.000 1289.240 ;
    END
  END dram_din0[6]
  PIN dram_din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 0.000 1948.470 4.000 ;
    END
  END dram_din0[7]
  PIN dram_din0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 1946.000 1668.330 1950.000 ;
    END
  END dram_din0[8]
  PIN dram_din0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 680.040 1950.000 680.640 ;
    END
  END dram_din0[9]
  PIN dram_dout0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 1946.000 959.930 1950.000 ;
    END
  END dram_dout0[0]
  PIN dram_dout0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 496.440 1950.000 497.040 ;
    END
  END dram_dout0[10]
  PIN dram_dout0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 1946.000 1520.210 1950.000 ;
    END
  END dram_dout0[11]
  PIN dram_dout0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1370.240 1950.000 1370.840 ;
    END
  END dram_dout0[12]
  PIN dram_dout0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1281.840 4.000 1282.440 ;
    END
  END dram_dout0[13]
  PIN dram_dout0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 1946.000 1304.470 1950.000 ;
    END
  END dram_dout0[14]
  PIN dram_dout0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1220.640 4.000 1221.240 ;
    END
  END dram_dout0[15]
  PIN dram_dout0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 119.040 1950.000 119.640 ;
    END
  END dram_dout0[16]
  PIN dram_dout0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.040 4.000 1241.640 ;
    END
  END dram_dout0[17]
  PIN dram_dout0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END dram_dout0[18]
  PIN dram_dout0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 788.840 1950.000 789.440 ;
    END
  END dram_dout0[19]
  PIN dram_dout0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 890.840 1950.000 891.440 ;
    END
  END dram_dout0[1]
  PIN dram_dout0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END dram_dout0[20]
  PIN dram_dout0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END dram_dout0[21]
  PIN dram_dout0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END dram_dout0[22]
  PIN dram_dout0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END dram_dout0[23]
  PIN dram_dout0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END dram_dout0[24]
  PIN dram_dout0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 1946.000 190.350 1950.000 ;
    END
  END dram_dout0[25]
  PIN dram_dout0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END dram_dout0[26]
  PIN dram_dout0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 98.640 1950.000 99.240 ;
    END
  END dram_dout0[27]
  PIN dram_dout0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1946.000 460.830 1950.000 ;
    END
  END dram_dout0[28]
  PIN dram_dout0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 1946.000 798.930 1950.000 ;
    END
  END dram_dout0[29]
  PIN dram_dout0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1652.440 1950.000 1653.040 ;
    END
  END dram_dout0[2]
  PIN dram_dout0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 1946.000 261.190 1950.000 ;
    END
  END dram_dout0[30]
  PIN dram_dout0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END dram_dout0[31]
  PIN dram_dout0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1207.040 1950.000 1207.640 ;
    END
  END dram_dout0[3]
  PIN dram_dout0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END dram_dout0[4]
  PIN dram_dout0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 1946.000 1855.090 1950.000 ;
    END
  END dram_dout0[5]
  PIN dram_dout0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 1946.000 966.370 1950.000 ;
    END
  END dram_dout0[6]
  PIN dram_dout0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END dram_dout0[7]
  PIN dram_dout0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 248.240 1950.000 248.840 ;
    END
  END dram_dout0[8]
  PIN dram_dout0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END dram_dout0[9]
  PIN dram_web0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1516.440 1950.000 1517.040 ;
    END
  END dram_web0
  PIN dram_wmask0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 1946.000 1330.230 1950.000 ;
    END
  END dram_wmask0[0]
  PIN dram_wmask0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 0.000 1407.510 4.000 ;
    END
  END dram_wmask0[1]
  PIN dram_wmask0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 1946.000 351.350 1950.000 ;
    END
  END dram_wmask0[2]
  PIN dram_wmask0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 0.000 1649.010 4.000 ;
    END
  END dram_wmask0[3]
  PIN icache_data_chip_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END icache_data_chip_en
  PIN icache_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1268.240 1950.000 1268.840 ;
    END
  END icache_data_in[0]
  PIN icache_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1946.000 32.570 1950.000 ;
    END
  END icache_data_in[10]
  PIN icache_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 1946.000 644.370 1950.000 ;
    END
  END icache_data_in[11]
  PIN icache_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 1946.000 927.730 1950.000 ;
    END
  END icache_data_in[12]
  PIN icache_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END icache_data_in[13]
  PIN icache_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.570 0.000 1719.850 4.000 ;
    END
  END icache_data_in[14]
  PIN icache_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 1946.000 1066.190 1950.000 ;
    END
  END icache_data_in[15]
  PIN icache_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.970 0.000 1784.250 4.000 ;
    END
  END icache_data_in[16]
  PIN icache_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1836.040 4.000 1836.640 ;
    END
  END icache_data_in[17]
  PIN icache_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.970 1946.000 1784.250 1950.000 ;
    END
  END icache_data_in[18]
  PIN icache_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END icache_data_in[19]
  PIN icache_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END icache_data_in[1]
  PIN icache_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END icache_data_in[20]
  PIN icache_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 1946.000 1130.590 1950.000 ;
    END
  END icache_data_in[21]
  PIN icache_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END icache_data_in[22]
  PIN icache_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END icache_data_in[23]
  PIN icache_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 323.040 1950.000 323.640 ;
    END
  END icache_data_in[24]
  PIN icache_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 1946.000 1117.710 1950.000 ;
    END
  END icache_data_in[25]
  PIN icache_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 809.240 1950.000 809.840 ;
    END
  END icache_data_in[26]
  PIN icache_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END icache_data_in[27]
  PIN icache_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 503.240 1950.000 503.840 ;
    END
  END icache_data_in[28]
  PIN icache_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.690 1946.000 1867.970 1950.000 ;
    END
  END icache_data_in[29]
  PIN icache_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1808.840 1950.000 1809.440 ;
    END
  END icache_data_in[2]
  PIN icache_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 214.240 1950.000 214.840 ;
    END
  END icache_data_in[30]
  PIN icache_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END icache_data_in[31]
  PIN icache_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END icache_data_in[3]
  PIN icache_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1856.440 4.000 1857.040 ;
    END
  END icache_data_in[4]
  PIN icache_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 1946.000 1674.770 1950.000 ;
    END
  END icache_data_in[5]
  PIN icache_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 904.440 1950.000 905.040 ;
    END
  END icache_data_in[6]
  PIN icache_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END icache_data_in[7]
  PIN icache_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 924.840 1950.000 925.440 ;
    END
  END icache_data_in[8]
  PIN icache_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.840 4.000 1180.440 ;
    END
  END icache_data_in[9]
  PIN icache_data_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 1946.000 811.810 1950.000 ;
    END
  END icache_data_index[0]
  PIN icache_data_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1666.040 1950.000 1666.640 ;
    END
  END icache_data_index[1]
  PIN icache_data_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 0.000 1681.210 4.000 ;
    END
  END icache_data_index[2]
  PIN icache_data_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.040 4.000 1479.640 ;
    END
  END icache_data_index[3]
  PIN icache_data_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.240 4.000 1268.840 ;
    END
  END icache_data_index[4]
  PIN icache_data_index[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.650 1946.000 1925.930 1950.000 ;
    END
  END icache_data_index[5]
  PIN icache_data_index[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END icache_data_index[6]
  PIN icache_data_index[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 0.000 1362.430 4.000 ;
    END
  END icache_data_index[7]
  PIN icache_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END icache_data_out[0]
  PIN icache_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1679.640 1950.000 1680.240 ;
    END
  END icache_data_out[10]
  PIN icache_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END icache_data_out[11]
  PIN icache_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1946.000 55.110 1950.000 ;
    END
  END icache_data_out[12]
  PIN icache_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 734.440 1950.000 735.040 ;
    END
  END icache_data_out[13]
  PIN icache_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1584.440 4.000 1585.040 ;
    END
  END icache_data_out[14]
  PIN icache_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 1946.000 177.470 1950.000 ;
    END
  END icache_data_out[15]
  PIN icache_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END icache_data_out[16]
  PIN icache_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 275.440 1950.000 276.040 ;
    END
  END icache_data_out[17]
  PIN icache_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END icache_data_out[18]
  PIN icache_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 282.240 1950.000 282.840 ;
    END
  END icache_data_out[19]
  PIN icache_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1946.000 428.630 1950.000 ;
    END
  END icache_data_out[1]
  PIN icache_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 1946.000 1797.130 1950.000 ;
    END
  END icache_data_out[20]
  PIN icache_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 1946.000 1375.310 1950.000 ;
    END
  END icache_data_out[21]
  PIN icache_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1173.040 1950.000 1173.640 ;
    END
  END icache_data_out[22]
  PIN icache_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 57.840 1950.000 58.440 ;
    END
  END icache_data_out[23]
  PIN icache_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1645.640 4.000 1646.240 ;
    END
  END icache_data_out[24]
  PIN icache_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.840 4.000 1452.440 ;
    END
  END icache_data_out[25]
  PIN icache_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END icache_data_out[26]
  PIN icache_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END icache_data_out[27]
  PIN icache_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.840 4.000 1214.440 ;
    END
  END icache_data_out[28]
  PIN icache_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END icache_data_out[29]
  PIN icache_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END icache_data_out[2]
  PIN icache_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1946.000 560.650 1950.000 ;
    END
  END icache_data_out[30]
  PIN icache_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 836.440 1950.000 837.040 ;
    END
  END icache_data_out[31]
  PIN icache_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END icache_data_out[3]
  PIN icache_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 1946.000 1343.110 1950.000 ;
    END
  END icache_data_out[4]
  PIN icache_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 1946.000 1597.490 1950.000 ;
    END
  END icache_data_out[5]
  PIN icache_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END icache_data_out[6]
  PIN icache_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1774.840 4.000 1775.440 ;
    END
  END icache_data_out[7]
  PIN icache_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END icache_data_out[8]
  PIN icache_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 1946.000 396.430 1950.000 ;
    END
  END icache_data_out[9]
  PIN icache_data_write_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1295.440 4.000 1296.040 ;
    END
  END icache_data_write_en
  PIN icache_tag_chip_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END icache_tag_chip_en
  PIN icache_tag_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END icache_tag_data_in[0]
  PIN icache_tag_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 1946.000 786.050 1950.000 ;
    END
  END icache_tag_data_in[10]
  PIN icache_tag_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.570 0.000 1880.850 4.000 ;
    END
  END icache_tag_data_in[11]
  PIN icache_tag_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1084.640 1950.000 1085.240 ;
    END
  END icache_tag_data_in[12]
  PIN icache_tag_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END icache_tag_data_in[13]
  PIN icache_tag_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END icache_tag_data_in[14]
  PIN icache_tag_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END icache_tag_data_in[15]
  PIN icache_tag_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1523.240 1950.000 1523.840 ;
    END
  END icache_tag_data_in[16]
  PIN icache_tag_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1761.240 1950.000 1761.840 ;
    END
  END icache_tag_data_in[17]
  PIN icache_tag_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1584.440 1950.000 1585.040 ;
    END
  END icache_tag_data_in[18]
  PIN icache_tag_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END icache_tag_data_in[19]
  PIN icache_tag_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 0.000 1481.570 4.000 ;
    END
  END icache_tag_data_in[1]
  PIN icache_tag_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END icache_tag_data_in[20]
  PIN icache_tag_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END icache_tag_data_in[21]
  PIN icache_tag_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END icache_tag_data_in[22]
  PIN icache_tag_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 1946.000 26.130 1950.000 ;
    END
  END icache_tag_data_in[23]
  PIN icache_tag_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END icache_tag_data_in[24]
  PIN icache_tag_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1550.440 1950.000 1551.040 ;
    END
  END icache_tag_data_in[25]
  PIN icache_tag_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 1946.000 992.130 1950.000 ;
    END
  END icache_tag_data_in[26]
  PIN icache_tag_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 0.000 1500.890 4.000 ;
    END
  END icache_tag_data_in[27]
  PIN icache_tag_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1193.440 1950.000 1194.040 ;
    END
  END icache_tag_data_in[28]
  PIN icache_tag_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1598.040 4.000 1598.640 ;
    END
  END icache_tag_data_in[29]
  PIN icache_tag_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END icache_tag_data_in[2]
  PIN icache_tag_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1411.040 1950.000 1411.640 ;
    END
  END icache_tag_data_in[30]
  PIN icache_tag_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END icache_tag_data_in[31]
  PIN icache_tag_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 1946.000 1745.610 1950.000 ;
    END
  END icache_tag_data_in[3]
  PIN icache_tag_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END icache_tag_data_in[4]
  PIN icache_tag_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 659.640 1950.000 660.240 ;
    END
  END icache_tag_data_in[5]
  PIN icache_tag_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 200.640 1950.000 201.240 ;
    END
  END icache_tag_data_in[6]
  PIN icache_tag_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 1946.000 1842.210 1950.000 ;
    END
  END icache_tag_data_in[7]
  PIN icache_tag_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 17.040 1950.000 17.640 ;
    END
  END icache_tag_data_in[8]
  PIN icache_tag_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END icache_tag_data_in[9]
  PIN icache_tag_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1863.240 1950.000 1863.840 ;
    END
  END icache_tag_index[0]
  PIN icache_tag_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1564.040 1950.000 1564.640 ;
    END
  END icache_tag_index[1]
  PIN icache_tag_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 0.000 1700.530 4.000 ;
    END
  END icache_tag_index[2]
  PIN icache_tag_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 911.240 1950.000 911.840 ;
    END
  END icache_tag_index[3]
  PIN icache_tag_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1946.000 1040.430 1950.000 ;
    END
  END icache_tag_index[4]
  PIN icache_tag_index[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 0.000 1887.290 4.000 ;
    END
  END icache_tag_index[5]
  PIN icache_tag_index[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1917.640 1950.000 1918.240 ;
    END
  END icache_tag_index[6]
  PIN icache_tag_index[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1064.240 1950.000 1064.840 ;
    END
  END icache_tag_index[7]
  PIN icache_tag_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END icache_tag_out[0]
  PIN icache_tag_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END icache_tag_out[10]
  PIN icache_tag_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END icache_tag_out[11]
  PIN icache_tag_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END icache_tag_out[12]
  PIN icache_tag_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 1946.000 1278.710 1950.000 ;
    END
  END icache_tag_out[13]
  PIN icache_tag_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 1946.000 505.910 1950.000 ;
    END
  END icache_tag_out[14]
  PIN icache_tag_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1931.240 1950.000 1931.840 ;
    END
  END icache_tag_out[15]
  PIN icache_tag_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 948.640 1950.000 949.240 ;
    END
  END icache_tag_out[16]
  PIN icache_tag_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 1946.000 1475.130 1950.000 ;
    END
  END icache_tag_out[17]
  PIN icache_tag_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.970 1946.000 1945.250 1950.000 ;
    END
  END icache_tag_out[18]
  PIN icache_tag_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 1946.000 605.730 1950.000 ;
    END
  END icache_tag_out[19]
  PIN icache_tag_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END icache_tag_out[1]
  PIN icache_tag_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1125.440 1950.000 1126.040 ;
    END
  END icache_tag_out[20]
  PIN icache_tag_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 0.000 1745.610 4.000 ;
    END
  END icache_tag_out[21]
  PIN icache_tag_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END icache_tag_out[22]
  PIN icache_tag_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 1946.000 1758.490 1950.000 ;
    END
  END icache_tag_out[23]
  PIN icache_tag_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1849.640 4.000 1850.240 ;
    END
  END icache_tag_out[24]
  PIN icache_tag_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 1946.000 222.550 1950.000 ;
    END
  END icache_tag_out[25]
  PIN icache_tag_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END icache_tag_out[26]
  PIN icache_tag_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END icache_tag_out[27]
  PIN icache_tag_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 1946.000 1732.730 1950.000 ;
    END
  END icache_tag_out[28]
  PIN icache_tag_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 1946.000 1694.090 1950.000 ;
    END
  END icache_tag_out[29]
  PIN icache_tag_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END icache_tag_out[2]
  PIN icache_tag_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 1946.000 1507.330 1950.000 ;
    END
  END icache_tag_out[30]
  PIN icache_tag_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END icache_tag_out[31]
  PIN icache_tag_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1179.840 1950.000 1180.440 ;
    END
  END icache_tag_out[3]
  PIN icache_tag_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.530 1946.000 1938.810 1950.000 ;
    END
  END icache_tag_out[4]
  PIN icache_tag_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 462.440 1950.000 463.040 ;
    END
  END icache_tag_out[5]
  PIN icache_tag_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 4.000 ;
    END
  END icache_tag_out[6]
  PIN icache_tag_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 0.000 1835.770 4.000 ;
    END
  END icache_tag_out[7]
  PIN icache_tag_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 863.640 1950.000 864.240 ;
    END
  END icache_tag_out[8]
  PIN icache_tag_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 1946.000 1001.790 1950.000 ;
    END
  END icache_tag_out[9]
  PIN icache_tag_write_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 0.000 1610.370 4.000 ;
    END
  END icache_tag_write_en
  PIN icache_write_data_mask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 469.240 1950.000 469.840 ;
    END
  END icache_write_data_mask[0]
  PIN icache_write_data_mask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 1946.000 1539.530 1950.000 ;
    END
  END icache_write_data_mask[1]
  PIN icache_write_data_mask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1876.840 4.000 1877.440 ;
    END
  END icache_write_data_mask[2]
  PIN icache_write_data_mask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1502.840 1950.000 1503.440 ;
    END
  END icache_write_data_mask[3]
  PIN icache_write_tag_mask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 1946.000 1426.830 1950.000 ;
    END
  END icache_write_tag_mask[0]
  PIN icache_write_tag_mask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END icache_write_tag_mask[1]
  PIN icache_write_tag_mask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END icache_write_tag_mask[2]
  PIN icache_write_tag_mask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END icache_write_tag_mask[3]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 1946.000 1336.670 1950.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 1946.000 1713.410 1950.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 0.000 1922.710 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 0.000 1771.370 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 714.040 1950.000 714.640 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 975.840 1950.000 976.440 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1618.440 4.000 1619.040 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 1946.000 773.170 1950.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1829.240 4.000 1829.840 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 1946.000 792.490 1950.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 1946.000 1401.070 1950.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 85.040 1950.000 85.640 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 0.000 1668.330 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 748.040 1950.000 748.640 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 0.000 1558.850 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 0.000 1565.290 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1016.640 1950.000 1017.240 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 1946.000 467.270 1950.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1946.000 299.830 1950.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 897.640 1950.000 898.240 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 1946.000 1014.670 1950.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1946.000 67.990 1950.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1946.000 145.270 1950.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.840 4.000 1350.440 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 132.640 1950.000 133.240 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1543.640 1950.000 1544.240 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.240 4.000 1370.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 700.440 1950.000 701.040 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 4.000 1200.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.130 1946.000 1552.410 1950.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 0.000 1545.970 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 1946.000 1565.290 1950.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 377.440 1950.000 378.040 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1343.040 1950.000 1343.640 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 918.040 1950.000 918.640 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 1946.000 1948.470 1950.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1938.040 1950.000 1938.640 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 1946.000 1317.350 1950.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1530.040 4.000 1530.640 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 625.640 1950.000 626.240 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 1946.000 518.790 1950.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.550 0.000 1909.830 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1638.840 1950.000 1639.440 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1329.440 4.000 1330.040 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1904.040 4.000 1904.640 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 564.440 1950.000 565.040 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 139.440 1950.000 140.040 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 0.000 1488.010 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1822.440 1950.000 1823.040 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 316.240 1950.000 316.840 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 1946.000 1323.790 1950.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1417.840 1950.000 1418.440 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 268.640 1950.000 269.240 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 1946.000 1874.410 1950.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 1946.000 1687.650 1950.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.770 1946.000 1591.050 1950.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 571.240 1950.000 571.840 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 1946.000 1349.550 1950.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1652.440 4.000 1653.040 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1424.640 4.000 1425.240 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1788.440 1950.000 1789.040 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1499.440 4.000 1500.040 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 557.640 1950.000 558.240 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1946.000 6.810 1950.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 1946.000 106.630 1950.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1946.000 48.670 1950.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 1946.000 895.530 1950.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.040 4.000 1309.640 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.770 0.000 1591.050 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 1946.000 921.290 1950.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1822.440 4.000 1823.040 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1003.040 1950.000 1003.640 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 1946.000 1887.290 1950.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 1946.000 1027.550 1950.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 1946.000 1481.570 1950.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1713.640 1950.000 1714.240 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1747.640 1950.000 1748.240 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.210 1946.000 1919.490 1950.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 1946.000 844.010 1950.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 1946.000 389.990 1950.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 438.640 1950.000 439.240 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 64.640 1950.000 65.240 ;
    END
  END io_out[9]
  PIN iram_addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 0.000 1533.090 4.000 ;
    END
  END iram_addr0[0]
  PIN iram_addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1802.040 4.000 1802.640 ;
    END
  END iram_addr0[1]
  PIN iram_addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 1946.000 447.950 1950.000 ;
    END
  END iram_addr0[2]
  PIN iram_addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END iram_addr0[3]
  PIN iram_addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1281.840 1950.000 1282.440 ;
    END
  END iram_addr0[4]
  PIN iram_addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END iram_addr0[5]
  PIN iram_addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 0.000 1726.290 4.000 ;
    END
  END iram_addr0[6]
  PIN iram_addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1863.240 4.000 1863.840 ;
    END
  END iram_addr0[7]
  PIN iram_clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1802.040 1950.000 1802.640 ;
    END
  END iram_clk0
  PIN iram_csb0_A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1946.000 100.190 1950.000 ;
    END
  END iram_csb0_A
  PIN iram_csb0_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END iram_csb0_B
  PIN iram_din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END iram_din0[0]
  PIN iram_din0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1275.040 1950.000 1275.640 ;
    END
  END iram_din0[10]
  PIN iram_din0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END iram_din0[11]
  PIN iram_din0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 1946.000 1526.650 1950.000 ;
    END
  END iram_din0[12]
  PIN iram_din0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END iram_din0[13]
  PIN iram_din0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 1946.000 422.190 1950.000 ;
    END
  END iram_din0[14]
  PIN iram_din0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END iram_din0[15]
  PIN iram_din0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END iram_din0[16]
  PIN iram_din0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1754.440 4.000 1755.040 ;
    END
  END iram_din0[17]
  PIN iram_din0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END iram_din0[18]
  PIN iram_din0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.290 1946.000 1803.570 1950.000 ;
    END
  END iram_din0[19]
  PIN iram_din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 1946.000 541.330 1950.000 ;
    END
  END iram_din0[1]
  PIN iram_din0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END iram_din0[20]
  PIN iram_din0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END iram_din0[21]
  PIN iram_din0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 1946.000 1771.370 1950.000 ;
    END
  END iram_din0[22]
  PIN iram_din0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1611.640 4.000 1612.240 ;
    END
  END iram_din0[23]
  PIN iram_din0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END iram_din0[24]
  PIN iram_din0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1523.240 4.000 1523.840 ;
    END
  END iram_din0[25]
  PIN iram_din0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 187.040 1950.000 187.640 ;
    END
  END iram_din0[26]
  PIN iram_din0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END iram_din0[27]
  PIN iram_din0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 0.000 1829.330 4.000 ;
    END
  END iram_din0[28]
  PIN iram_din0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 1946.000 1355.990 1950.000 ;
    END
  END iram_din0[29]
  PIN iram_din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END iram_din0[2]
  PIN iram_din0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END iram_din0[30]
  PIN iram_din0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 357.040 1950.000 357.640 ;
    END
  END iram_din0[31]
  PIN iram_din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END iram_din0[3]
  PIN iram_din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END iram_din0[4]
  PIN iram_din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 370.640 1950.000 371.240 ;
    END
  END iram_din0[5]
  PIN iram_din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 1946.000 1584.610 1950.000 ;
    END
  END iram_din0[6]
  PIN iram_din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 1946.000 1188.550 1950.000 ;
    END
  END iram_din0[7]
  PIN iram_din0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 1946.000 567.090 1950.000 ;
    END
  END iram_din0[8]
  PIN iram_din0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1686.440 1950.000 1687.040 ;
    END
  END iram_din0[9]
  PIN iram_dout0_A[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END iram_dout0_A[0]
  PIN iram_dout0_A[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 1946.000 1207.870 1950.000 ;
    END
  END iram_dout0_A[10]
  PIN iram_dout0_A[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1322.640 1950.000 1323.240 ;
    END
  END iram_dout0_A[11]
  PIN iram_dout0_A[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 0.000 1597.490 4.000 ;
    END
  END iram_dout0_A[12]
  PIN iram_dout0_A[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 931.640 1950.000 932.240 ;
    END
  END iram_dout0_A[13]
  PIN iram_dout0_A[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END iram_dout0_A[14]
  PIN iram_dout0_A[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 720.840 1950.000 721.440 ;
    END
  END iram_dout0_A[15]
  PIN iram_dout0_A[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 1946.000 831.130 1950.000 ;
    END
  END iram_dout0_A[16]
  PIN iram_dout0_A[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 1946.000 625.050 1950.000 ;
    END
  END iram_dout0_A[17]
  PIN iram_dout0_A[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 632.440 1950.000 633.040 ;
    END
  END iram_dout0_A[18]
  PIN iram_dout0_A[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 1946.000 695.890 1950.000 ;
    END
  END iram_dout0_A[19]
  PIN iram_dout0_A[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 1946.000 818.250 1950.000 ;
    END
  END iram_dout0_A[1]
  PIN iram_dout0_A[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 146.240 1950.000 146.840 ;
    END
  END iram_dout0_A[20]
  PIN iram_dout0_A[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END iram_dout0_A[21]
  PIN iram_dout0_A[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1897.240 1950.000 1897.840 ;
    END
  END iram_dout0_A[22]
  PIN iram_dout0_A[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 591.640 1950.000 592.240 ;
    END
  END iram_dout0_A[23]
  PIN iram_dout0_A[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 1946.000 953.490 1950.000 ;
    END
  END iram_dout0_A[24]
  PIN iram_dout0_A[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 1946.000 1156.350 1950.000 ;
    END
  END iram_dout0_A[25]
  PIN iram_dout0_A[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1468.840 1950.000 1469.440 ;
    END
  END iram_dout0_A[26]
  PIN iram_dout0_A[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END iram_dout0_A[27]
  PIN iram_dout0_A[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 1946.000 708.770 1950.000 ;
    END
  END iram_dout0_A[28]
  PIN iram_dout0_A[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END iram_dout0_A[29]
  PIN iram_dout0_A[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END iram_dout0_A[2]
  PIN iram_dout0_A[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 363.840 1950.000 364.440 ;
    END
  END iram_dout0_A[30]
  PIN iram_dout0_A[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1570.840 4.000 1571.440 ;
    END
  END iram_dout0_A[31]
  PIN iram_dout0_A[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1057.440 1950.000 1058.040 ;
    END
  END iram_dout0_A[3]
  PIN iram_dout0_A[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 1946.000 1201.430 1950.000 ;
    END
  END iram_dout0_A[4]
  PIN iram_dout0_A[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END iram_dout0_A[5]
  PIN iram_dout0_A[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1023.440 1950.000 1024.040 ;
    END
  END iram_dout0_A[6]
  PIN iram_dout0_A[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1700.040 1950.000 1700.640 ;
    END
  END iram_dout0_A[7]
  PIN iram_dout0_A[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END iram_dout0_A[8]
  PIN iram_dout0_A[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 1946.000 138.830 1950.000 ;
    END
  END iram_dout0_A[9]
  PIN iram_dout0_B[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1849.640 1950.000 1850.240 ;
    END
  END iram_dout0_B[0]
  PIN iram_dout0_B[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END iram_dout0_B[10]
  PIN iram_dout0_B[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 1946.000 863.330 1950.000 ;
    END
  END iram_dout0_B[11]
  PIN iram_dout0_B[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END iram_dout0_B[12]
  PIN iram_dout0_B[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 1946.000 473.710 1950.000 ;
    END
  END iram_dout0_B[13]
  PIN iram_dout0_B[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 0.000 1520.210 4.000 ;
    END
  END iram_dout0_B[14]
  PIN iram_dout0_B[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 1946.000 1533.090 1950.000 ;
    END
  END iram_dout0_B[15]
  PIN iram_dout0_B[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 955.440 1950.000 956.040 ;
    END
  END iram_dout0_B[16]
  PIN iram_dout0_B[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 707.240 1950.000 707.840 ;
    END
  END iram_dout0_B[17]
  PIN iram_dout0_B[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END iram_dout0_B[18]
  PIN iram_dout0_B[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END iram_dout0_B[19]
  PIN iram_dout0_B[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END iram_dout0_B[1]
  PIN iram_dout0_B[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 523.640 1950.000 524.240 ;
    END
  END iram_dout0_B[20]
  PIN iram_dout0_B[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 1946.000 1752.050 1950.000 ;
    END
  END iram_dout0_B[21]
  PIN iram_dout0_B[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1105.040 1950.000 1105.640 ;
    END
  END iram_dout0_B[22]
  PIN iram_dout0_B[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1781.640 1950.000 1782.240 ;
    END
  END iram_dout0_B[23]
  PIN iram_dout0_B[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 1946.000 1706.970 1950.000 ;
    END
  END iram_dout0_B[24]
  PIN iram_dout0_B[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END iram_dout0_B[25]
  PIN iram_dout0_B[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 482.840 1950.000 483.440 ;
    END
  END iram_dout0_B[26]
  PIN iram_dout0_B[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 0.000 1616.810 4.000 ;
    END
  END iram_dout0_B[27]
  PIN iram_dout0_B[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1632.040 4.000 1632.640 ;
    END
  END iram_dout0_B[28]
  PIN iram_dout0_B[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 166.640 1950.000 167.240 ;
    END
  END iram_dout0_B[29]
  PIN iram_dout0_B[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 0.000 1381.750 4.000 ;
    END
  END iram_dout0_B[2]
  PIN iram_dout0_B[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END iram_dout0_B[30]
  PIN iram_dout0_B[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1870.040 1950.000 1870.640 ;
    END
  END iram_dout0_B[31]
  PIN iram_dout0_B[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END iram_dout0_B[3]
  PIN iram_dout0_B[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 0.000 1687.650 4.000 ;
    END
  END iram_dout0_B[4]
  PIN iram_dout0_B[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 1946.000 183.910 1950.000 ;
    END
  END iram_dout0_B[5]
  PIN iram_dout0_B[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END iram_dout0_B[6]
  PIN iram_dout0_B[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END iram_dout0_B[7]
  PIN iram_dout0_B[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 1946.000 151.710 1950.000 ;
    END
  END iram_dout0_B[8]
  PIN iram_dout0_B[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END iram_dout0_B[9]
  PIN iram_web0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 1946.000 1285.150 1950.000 ;
    END
  END iram_web0
  PIN iram_wmask0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1591.240 4.000 1591.840 ;
    END
  END iram_wmask0[0]
  PIN iram_wmask0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END iram_wmask0[1]
  PIN iram_wmask0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 530.440 1950.000 531.040 ;
    END
  END iram_wmask0[2]
  PIN iram_wmask0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.110 0.000 1903.390 4.000 ;
    END
  END iram_wmask0[3]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 1946.000 979.250 1950.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 1946.000 1610.370 1950.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 1946.000 534.890 1950.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1475.640 1950.000 1476.240 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.170 0.000 1655.450 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 1946.000 1777.810 1950.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.410 1946.000 1629.690 1950.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 1946.000 670.130 1950.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 180.240 1950.000 180.840 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1897.240 4.000 1897.840 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 1946.000 1240.070 1950.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1356.640 4.000 1357.240 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1037.040 1950.000 1037.640 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 1946.000 228.990 1950.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 693.640 1950.000 694.240 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 350.240 1950.000 350.840 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1438.240 1950.000 1438.840 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 336.640 1950.000 337.240 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1200.240 1950.000 1200.840 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 754.840 1950.000 755.440 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1091.440 1950.000 1092.040 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 397.840 1950.000 398.440 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 0.000 1623.250 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1842.840 1950.000 1843.440 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 71.440 1950.000 72.040 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 1946.000 1513.770 1950.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.890 1946.000 1578.170 1950.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 343.440 1950.000 344.040 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 0.000 1842.210 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 1946.000 1149.910 1950.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 1946.000 267.630 1950.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 1946.000 286.950 1950.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1118.640 1950.000 1119.240 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 0.000 1739.170 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 666.440 1950.000 667.040 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 795.640 1950.000 796.240 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1890.440 4.000 1891.040 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1254.640 1950.000 1255.240 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 1946.000 525.230 1950.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 1946.000 1681.210 1950.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 1946.000 657.250 1950.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1946.000 80.870 1950.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 455.640 1950.000 456.240 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1604.840 4.000 1605.440 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1944.840 4.000 1945.440 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 1946.000 901.970 1950.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1302.240 1950.000 1302.840 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 255.040 1950.000 255.640 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1509.640 1950.000 1510.240 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 448.840 1950.000 449.440 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 782.040 1950.000 782.640 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 0.000 1494.450 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 1946.000 940.610 1950.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1404.240 1950.000 1404.840 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 1946.000 1091.950 1950.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 989.440 1950.000 990.040 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1132.240 1950.000 1132.840 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1462.040 1950.000 1462.640 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1946.000 689.450 1950.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.610 1946.000 1822.890 1950.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 1946.000 1053.310 1950.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 1946.000 1471.910 1950.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1349.840 1950.000 1350.440 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 1946.000 1272.270 1950.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.730 1946.000 1810.010 1950.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 1946.000 125.950 1950.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 1946.000 248.310 1950.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 1946.000 1407.510 1950.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 1946.000 1194.990 1950.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 1946.000 1446.150 1950.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 1946.000 409.310 1950.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1186.640 4.000 1187.240 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1938.040 4.000 1938.640 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1363.440 1950.000 1364.040 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 1946.000 1220.750 1950.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1946.000 579.970 1950.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 1946.000 435.070 1950.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 1946.000 599.290 1950.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 0.000 1246.510 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 775.240 1950.000 775.840 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 982.640 1950.000 983.240 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 1946.000 631.490 1950.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 1946.000 1488.010 1950.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 0.000 1194.990 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1795.240 1950.000 1795.840 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 1946.000 1137.030 1950.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 945.240 1950.000 945.840 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 1946.000 882.650 1950.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1686.440 4.000 1687.040 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.290 0.000 1803.570 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1720.440 1950.000 1721.040 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 1946.000 1298.030 1950.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 1946.000 766.730 1950.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1870.040 4.000 1870.640 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1836.040 1950.000 1836.640 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 1946.000 715.210 1950.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1591.240 1950.000 1591.840 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 0.000 1874.410 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.240 4.000 1404.840 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 856.840 1950.000 857.440 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 0.000 1764.930 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1329.440 1950.000 1330.040 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 1946.000 1079.070 1950.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1944.840 1950.000 1945.440 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 0.000 1752.050 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 1946.000 1169.230 1950.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1050.640 1950.000 1051.240 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 261.840 1950.000 262.440 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 1946.000 216.110 1950.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 1946.000 312.710 1950.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 686.840 1950.000 687.440 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 91.840 1950.000 92.440 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 1946.000 1291.590 1950.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 1946.000 1700.530 1950.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 112.240 1950.000 112.840 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 1946.000 1494.450 1950.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1910.840 1950.000 1911.440 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1946.000 87.310 1950.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1213.840 1950.000 1214.440 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1815.640 4.000 1816.240 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 598.440 1950.000 599.040 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 850.040 1950.000 850.640 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 1946.000 592.850 1950.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.890 0.000 1578.170 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 418.240 1950.000 418.840 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 1946.000 158.150 1950.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1625.240 1950.000 1625.840 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 0.000 1526.650 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1516.440 4.000 1517.040 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1672.840 4.000 1673.440 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 0.000 1732.730 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 1946.000 1636.130 1950.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.040 4.000 1768.640 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 0.000 1423.610 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 1946.000 164.590 1950.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1363.440 4.000 1364.040 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 425.040 1950.000 425.640 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1383.840 1950.000 1384.440 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1145.840 1950.000 1146.440 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.450 0.000 1893.730 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 1946.000 203.230 1950.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 37.440 1950.000 38.040 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 0.000 1584.610 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1322.640 4.000 1323.240 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.170 1946.000 1655.450 1950.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 0.000 1310.910 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 969.040 1950.000 969.640 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 550.840 1950.000 551.440 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1288.640 1950.000 1289.240 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1139.040 1950.000 1139.640 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1946.000 612.170 1950.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 159.840 1950.000 160.440 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1625.240 4.000 1625.840 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1438.240 4.000 1438.840 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 1946.000 280.510 1950.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.990 0.000 1916.270 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 207.440 1950.000 208.040 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 1946.000 332.030 1950.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 1946.000 856.890 1950.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 10.240 1950.000 10.840 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1397.440 1950.000 1398.040 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 1946.000 383.550 1950.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1509.640 4.000 1510.240 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 612.040 1950.000 612.640 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 1946.000 837.570 1950.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 884.040 1950.000 884.640 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 1946.000 415.750 1950.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 1946.000 1861.530 1950.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1946.000 779.610 1950.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.330 1946.000 1906.610 1950.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1946.000 19.690 1950.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 0.000 1790.690 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1856.440 1950.000 1857.040 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 0.000 1420.390 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 0.000 1259.390 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1489.240 1950.000 1489.840 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 639.240 1950.000 639.840 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1924.440 1950.000 1925.040 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1946.000 61.550 1950.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 1946.000 1388.190 1950.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1309.040 1950.000 1309.640 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1672.840 1950.000 1673.440 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 23.840 1950.000 24.440 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1098.240 1950.000 1098.840 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 1946.000 93.750 1950.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 877.240 1950.000 877.840 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 802.440 1950.000 803.040 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1448.440 1950.000 1449.040 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1261.440 1950.000 1262.040 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.410 0.000 1629.690 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1946.000 824.690 1950.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 0.000 1507.330 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1734.040 1950.000 1734.640 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 1946.000 1124.150 1950.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 1946.000 869.770 1950.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 1946.000 293.390 1950.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 1946.000 1162.790 1950.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1417.840 4.000 1418.440 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 544.040 1950.000 544.640 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1152.640 1950.000 1153.240 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1768.040 1950.000 1768.640 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 1946.000 13.250 1950.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 0.000 1777.810 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 1946.000 1616.810 1950.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.770 1946.000 1913.050 1950.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1946.000 1008.230 1950.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 1946.000 1420.390 1950.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 173.440 1950.000 174.040 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 1946.000 1394.630 1950.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 78.240 1950.000 78.840 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 221.040 1950.000 221.640 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1043.840 1950.000 1044.440 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 1946.000 1661.890 1950.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 1946.000 171.030 1950.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 1946.000 74.430 1950.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.040 4.000 1666.640 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 1946.000 1459.030 1950.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 431.840 1950.000 432.440 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.040 4.000 1564.640 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 1946.000 1739.170 1950.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 1946.000 637.930 1950.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 1946.000 512.350 1950.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 1946.000 914.850 1950.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 1946.000 1021.110 1950.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 1946.000 1046.870 1950.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 1946.000 319.150 1950.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 3.440 1950.000 4.040 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 727.640 1950.000 728.240 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 1946.000 573.530 1950.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 0.000 1111.270 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 1946.000 344.910 1950.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 44.240 1950.000 44.840 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 0.000 1861.530 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 1946.000 1642.570 1950.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.890 0.000 1900.170 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 489.640 1950.000 490.240 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 1946.000 1764.930 1950.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1946.000 113.070 1950.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1815.640 1950.000 1816.240 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.370 0.000 1848.650 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 1946.000 650.810 1950.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 741.240 1950.000 741.840 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1931.240 4.000 1931.840 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 289.040 1950.000 289.640 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1706.840 1950.000 1707.440 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 1946.000 1829.330 1950.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1315.840 4.000 1316.440 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 1946.000 734.530 1950.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 1946.000 1623.250 1950.000 ;
    END
  END la_oenb[9]
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 822.840 1950.000 823.440 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1936.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1936.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1936.880 ;
    END
  END vssd1
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.840 4.000 1146.440 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1227.440 1950.000 1228.040 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1842.840 4.000 1843.440 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 0.000 1285.150 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 1946.000 1790.690 1950.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.090 1946.000 1932.370 1950.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1774.840 1950.000 1775.440 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1077.840 1950.000 1078.440 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 241.440 1950.000 242.040 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 1946.000 1098.390 1950.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 0.000 1278.710 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 0.000 1816.450 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 0.000 1220.750 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1808.840 4.000 1809.440 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1632.040 1950.000 1632.640 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 1946.000 1433.270 1950.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 1946.000 908.410 1950.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1234.240 1950.000 1234.840 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 0.000 1706.970 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 0.000 1636.130 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 227.840 1950.000 228.440 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 843.240 1950.000 843.840 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1924.440 4.000 1925.040 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.570 1946.000 1719.850 1950.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1356.640 1950.000 1357.240 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 1946.000 850.450 1950.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 1946.000 1368.870 1950.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.240 4.000 1472.840 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1496.040 1950.000 1496.640 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 1946.000 1465.470 1950.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1876.840 1950.000 1877.440 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 870.440 1950.000 871.040 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 0.000 1442.930 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 1946.000 1252.950 1950.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1946.000 39.010 1950.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1445.040 1950.000 1445.640 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 761.640 1950.000 762.240 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1030.240 1950.000 1030.840 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 1946.000 1259.390 1950.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.890 1946.000 1900.170 1950.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 193.840 1950.000 194.440 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1295.440 1950.000 1296.040 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.570 1946.000 1880.850 1950.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1946.000 1233.630 1950.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 309.440 1950.000 310.040 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 1946.000 1182.110 1950.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 0.000 1343.110 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1485.840 4.000 1486.440 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 1946.000 370.670 1950.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 1946.000 889.090 1950.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1946.000 454.390 1950.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 578.040 1950.000 578.640 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1577.640 1950.000 1578.240 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 0.000 1169.230 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 1482.440 1950.000 1483.040 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 1946.000 1246.510 1950.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 1946.000 1227.190 1950.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1795.240 4.000 1795.840 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 1946.000 209.670 1950.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.840 4.000 1639.440 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1946.000 938.440 1950.000 939.040 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1944.420 1936.725 ;
      LAYER met1 ;
        RECT 0.070 10.640 1948.490 1936.880 ;
      LAYER met2 ;
        RECT 0.650 1945.720 6.250 1946.570 ;
        RECT 7.090 1945.720 12.690 1946.570 ;
        RECT 13.530 1945.720 19.130 1946.570 ;
        RECT 19.970 1945.720 25.570 1946.570 ;
        RECT 26.410 1945.720 32.010 1946.570 ;
        RECT 32.850 1945.720 38.450 1946.570 ;
        RECT 39.290 1945.720 44.890 1946.570 ;
        RECT 45.730 1945.720 48.110 1946.570 ;
        RECT 48.950 1945.720 54.550 1946.570 ;
        RECT 55.390 1945.720 60.990 1946.570 ;
        RECT 61.830 1945.720 67.430 1946.570 ;
        RECT 68.270 1945.720 73.870 1946.570 ;
        RECT 74.710 1945.720 80.310 1946.570 ;
        RECT 81.150 1945.720 86.750 1946.570 ;
        RECT 87.590 1945.720 93.190 1946.570 ;
        RECT 94.030 1945.720 99.630 1946.570 ;
        RECT 100.470 1945.720 106.070 1946.570 ;
        RECT 106.910 1945.720 112.510 1946.570 ;
        RECT 113.350 1945.720 118.950 1946.570 ;
        RECT 119.790 1945.720 125.390 1946.570 ;
        RECT 126.230 1945.720 131.830 1946.570 ;
        RECT 132.670 1945.720 138.270 1946.570 ;
        RECT 139.110 1945.720 144.710 1946.570 ;
        RECT 145.550 1945.720 151.150 1946.570 ;
        RECT 151.990 1945.720 157.590 1946.570 ;
        RECT 158.430 1945.720 164.030 1946.570 ;
        RECT 164.870 1945.720 170.470 1946.570 ;
        RECT 171.310 1945.720 176.910 1946.570 ;
        RECT 177.750 1945.720 183.350 1946.570 ;
        RECT 184.190 1945.720 189.790 1946.570 ;
        RECT 190.630 1945.720 196.230 1946.570 ;
        RECT 197.070 1945.720 202.670 1946.570 ;
        RECT 203.510 1945.720 209.110 1946.570 ;
        RECT 209.950 1945.720 215.550 1946.570 ;
        RECT 216.390 1945.720 221.990 1946.570 ;
        RECT 222.830 1945.720 228.430 1946.570 ;
        RECT 229.270 1945.720 234.870 1946.570 ;
        RECT 235.710 1945.720 241.310 1946.570 ;
        RECT 242.150 1945.720 247.750 1946.570 ;
        RECT 248.590 1945.720 254.190 1946.570 ;
        RECT 255.030 1945.720 260.630 1946.570 ;
        RECT 261.470 1945.720 267.070 1946.570 ;
        RECT 267.910 1945.720 273.510 1946.570 ;
        RECT 274.350 1945.720 279.950 1946.570 ;
        RECT 280.790 1945.720 286.390 1946.570 ;
        RECT 287.230 1945.720 292.830 1946.570 ;
        RECT 293.670 1945.720 299.270 1946.570 ;
        RECT 300.110 1945.720 305.710 1946.570 ;
        RECT 306.550 1945.720 312.150 1946.570 ;
        RECT 312.990 1945.720 318.590 1946.570 ;
        RECT 319.430 1945.720 325.030 1946.570 ;
        RECT 325.870 1945.720 331.470 1946.570 ;
        RECT 332.310 1945.720 337.910 1946.570 ;
        RECT 338.750 1945.720 344.350 1946.570 ;
        RECT 345.190 1945.720 350.790 1946.570 ;
        RECT 351.630 1945.720 357.230 1946.570 ;
        RECT 358.070 1945.720 363.670 1946.570 ;
        RECT 364.510 1945.720 370.110 1946.570 ;
        RECT 370.950 1945.720 376.550 1946.570 ;
        RECT 377.390 1945.720 382.990 1946.570 ;
        RECT 383.830 1945.720 389.430 1946.570 ;
        RECT 390.270 1945.720 395.870 1946.570 ;
        RECT 396.710 1945.720 402.310 1946.570 ;
        RECT 403.150 1945.720 408.750 1946.570 ;
        RECT 409.590 1945.720 415.190 1946.570 ;
        RECT 416.030 1945.720 421.630 1946.570 ;
        RECT 422.470 1945.720 428.070 1946.570 ;
        RECT 428.910 1945.720 434.510 1946.570 ;
        RECT 435.350 1945.720 440.950 1946.570 ;
        RECT 441.790 1945.720 447.390 1946.570 ;
        RECT 448.230 1945.720 453.830 1946.570 ;
        RECT 454.670 1945.720 460.270 1946.570 ;
        RECT 461.110 1945.720 466.710 1946.570 ;
        RECT 467.550 1945.720 473.150 1946.570 ;
        RECT 473.990 1945.720 479.590 1946.570 ;
        RECT 480.430 1945.720 486.030 1946.570 ;
        RECT 486.870 1945.720 492.470 1946.570 ;
        RECT 493.310 1945.720 498.910 1946.570 ;
        RECT 499.750 1945.720 505.350 1946.570 ;
        RECT 506.190 1945.720 511.790 1946.570 ;
        RECT 512.630 1945.720 518.230 1946.570 ;
        RECT 519.070 1945.720 524.670 1946.570 ;
        RECT 525.510 1945.720 527.890 1946.570 ;
        RECT 528.730 1945.720 534.330 1946.570 ;
        RECT 535.170 1945.720 540.770 1946.570 ;
        RECT 541.610 1945.720 547.210 1946.570 ;
        RECT 548.050 1945.720 553.650 1946.570 ;
        RECT 554.490 1945.720 560.090 1946.570 ;
        RECT 560.930 1945.720 566.530 1946.570 ;
        RECT 567.370 1945.720 572.970 1946.570 ;
        RECT 573.810 1945.720 579.410 1946.570 ;
        RECT 580.250 1945.720 585.850 1946.570 ;
        RECT 586.690 1945.720 592.290 1946.570 ;
        RECT 593.130 1945.720 598.730 1946.570 ;
        RECT 599.570 1945.720 605.170 1946.570 ;
        RECT 606.010 1945.720 611.610 1946.570 ;
        RECT 612.450 1945.720 618.050 1946.570 ;
        RECT 618.890 1945.720 624.490 1946.570 ;
        RECT 625.330 1945.720 630.930 1946.570 ;
        RECT 631.770 1945.720 637.370 1946.570 ;
        RECT 638.210 1945.720 643.810 1946.570 ;
        RECT 644.650 1945.720 650.250 1946.570 ;
        RECT 651.090 1945.720 656.690 1946.570 ;
        RECT 657.530 1945.720 663.130 1946.570 ;
        RECT 663.970 1945.720 669.570 1946.570 ;
        RECT 670.410 1945.720 676.010 1946.570 ;
        RECT 676.850 1945.720 682.450 1946.570 ;
        RECT 683.290 1945.720 688.890 1946.570 ;
        RECT 689.730 1945.720 695.330 1946.570 ;
        RECT 696.170 1945.720 701.770 1946.570 ;
        RECT 702.610 1945.720 708.210 1946.570 ;
        RECT 709.050 1945.720 714.650 1946.570 ;
        RECT 715.490 1945.720 721.090 1946.570 ;
        RECT 721.930 1945.720 727.530 1946.570 ;
        RECT 728.370 1945.720 733.970 1946.570 ;
        RECT 734.810 1945.720 740.410 1946.570 ;
        RECT 741.250 1945.720 746.850 1946.570 ;
        RECT 747.690 1945.720 753.290 1946.570 ;
        RECT 754.130 1945.720 759.730 1946.570 ;
        RECT 760.570 1945.720 766.170 1946.570 ;
        RECT 767.010 1945.720 772.610 1946.570 ;
        RECT 773.450 1945.720 779.050 1946.570 ;
        RECT 779.890 1945.720 785.490 1946.570 ;
        RECT 786.330 1945.720 791.930 1946.570 ;
        RECT 792.770 1945.720 798.370 1946.570 ;
        RECT 799.210 1945.720 804.810 1946.570 ;
        RECT 805.650 1945.720 811.250 1946.570 ;
        RECT 812.090 1945.720 817.690 1946.570 ;
        RECT 818.530 1945.720 824.130 1946.570 ;
        RECT 824.970 1945.720 830.570 1946.570 ;
        RECT 831.410 1945.720 837.010 1946.570 ;
        RECT 837.850 1945.720 843.450 1946.570 ;
        RECT 844.290 1945.720 849.890 1946.570 ;
        RECT 850.730 1945.720 856.330 1946.570 ;
        RECT 857.170 1945.720 862.770 1946.570 ;
        RECT 863.610 1945.720 869.210 1946.570 ;
        RECT 870.050 1945.720 875.650 1946.570 ;
        RECT 876.490 1945.720 882.090 1946.570 ;
        RECT 882.930 1945.720 888.530 1946.570 ;
        RECT 889.370 1945.720 894.970 1946.570 ;
        RECT 895.810 1945.720 901.410 1946.570 ;
        RECT 902.250 1945.720 907.850 1946.570 ;
        RECT 908.690 1945.720 914.290 1946.570 ;
        RECT 915.130 1945.720 920.730 1946.570 ;
        RECT 921.570 1945.720 927.170 1946.570 ;
        RECT 928.010 1945.720 933.610 1946.570 ;
        RECT 934.450 1945.720 940.050 1946.570 ;
        RECT 940.890 1945.720 946.490 1946.570 ;
        RECT 947.330 1945.720 952.930 1946.570 ;
        RECT 953.770 1945.720 959.370 1946.570 ;
        RECT 960.210 1945.720 965.810 1946.570 ;
        RECT 966.650 1945.720 972.250 1946.570 ;
        RECT 973.090 1945.720 978.690 1946.570 ;
        RECT 979.530 1945.720 985.130 1946.570 ;
        RECT 985.970 1945.720 991.570 1946.570 ;
        RECT 992.410 1945.720 998.010 1946.570 ;
        RECT 998.850 1945.720 1001.230 1946.570 ;
        RECT 1002.070 1945.720 1007.670 1946.570 ;
        RECT 1008.510 1945.720 1014.110 1946.570 ;
        RECT 1014.950 1945.720 1020.550 1946.570 ;
        RECT 1021.390 1945.720 1026.990 1946.570 ;
        RECT 1027.830 1945.720 1033.430 1946.570 ;
        RECT 1034.270 1945.720 1039.870 1946.570 ;
        RECT 1040.710 1945.720 1046.310 1946.570 ;
        RECT 1047.150 1945.720 1052.750 1946.570 ;
        RECT 1053.590 1945.720 1059.190 1946.570 ;
        RECT 1060.030 1945.720 1065.630 1946.570 ;
        RECT 1066.470 1945.720 1072.070 1946.570 ;
        RECT 1072.910 1945.720 1078.510 1946.570 ;
        RECT 1079.350 1945.720 1084.950 1946.570 ;
        RECT 1085.790 1945.720 1091.390 1946.570 ;
        RECT 1092.230 1945.720 1097.830 1946.570 ;
        RECT 1098.670 1945.720 1104.270 1946.570 ;
        RECT 1105.110 1945.720 1110.710 1946.570 ;
        RECT 1111.550 1945.720 1117.150 1946.570 ;
        RECT 1117.990 1945.720 1123.590 1946.570 ;
        RECT 1124.430 1945.720 1130.030 1946.570 ;
        RECT 1130.870 1945.720 1136.470 1946.570 ;
        RECT 1137.310 1945.720 1142.910 1946.570 ;
        RECT 1143.750 1945.720 1149.350 1946.570 ;
        RECT 1150.190 1945.720 1155.790 1946.570 ;
        RECT 1156.630 1945.720 1162.230 1946.570 ;
        RECT 1163.070 1945.720 1168.670 1946.570 ;
        RECT 1169.510 1945.720 1175.110 1946.570 ;
        RECT 1175.950 1945.720 1181.550 1946.570 ;
        RECT 1182.390 1945.720 1187.990 1946.570 ;
        RECT 1188.830 1945.720 1194.430 1946.570 ;
        RECT 1195.270 1945.720 1200.870 1946.570 ;
        RECT 1201.710 1945.720 1207.310 1946.570 ;
        RECT 1208.150 1945.720 1213.750 1946.570 ;
        RECT 1214.590 1945.720 1220.190 1946.570 ;
        RECT 1221.030 1945.720 1226.630 1946.570 ;
        RECT 1227.470 1945.720 1233.070 1946.570 ;
        RECT 1233.910 1945.720 1239.510 1946.570 ;
        RECT 1240.350 1945.720 1245.950 1946.570 ;
        RECT 1246.790 1945.720 1252.390 1946.570 ;
        RECT 1253.230 1945.720 1258.830 1946.570 ;
        RECT 1259.670 1945.720 1265.270 1946.570 ;
        RECT 1266.110 1945.720 1271.710 1946.570 ;
        RECT 1272.550 1945.720 1278.150 1946.570 ;
        RECT 1278.990 1945.720 1284.590 1946.570 ;
        RECT 1285.430 1945.720 1291.030 1946.570 ;
        RECT 1291.870 1945.720 1297.470 1946.570 ;
        RECT 1298.310 1945.720 1303.910 1946.570 ;
        RECT 1304.750 1945.720 1310.350 1946.570 ;
        RECT 1311.190 1945.720 1316.790 1946.570 ;
        RECT 1317.630 1945.720 1323.230 1946.570 ;
        RECT 1324.070 1945.720 1329.670 1946.570 ;
        RECT 1330.510 1945.720 1336.110 1946.570 ;
        RECT 1336.950 1945.720 1342.550 1946.570 ;
        RECT 1343.390 1945.720 1348.990 1946.570 ;
        RECT 1349.830 1945.720 1355.430 1946.570 ;
        RECT 1356.270 1945.720 1361.870 1946.570 ;
        RECT 1362.710 1945.720 1368.310 1946.570 ;
        RECT 1369.150 1945.720 1374.750 1946.570 ;
        RECT 1375.590 1945.720 1381.190 1946.570 ;
        RECT 1382.030 1945.720 1387.630 1946.570 ;
        RECT 1388.470 1945.720 1394.070 1946.570 ;
        RECT 1394.910 1945.720 1400.510 1946.570 ;
        RECT 1401.350 1945.720 1406.950 1946.570 ;
        RECT 1407.790 1945.720 1413.390 1946.570 ;
        RECT 1414.230 1945.720 1419.830 1946.570 ;
        RECT 1420.670 1945.720 1426.270 1946.570 ;
        RECT 1427.110 1945.720 1432.710 1946.570 ;
        RECT 1433.550 1945.720 1439.150 1946.570 ;
        RECT 1439.990 1945.720 1445.590 1946.570 ;
        RECT 1446.430 1945.720 1452.030 1946.570 ;
        RECT 1452.870 1945.720 1458.470 1946.570 ;
        RECT 1459.310 1945.720 1464.910 1946.570 ;
        RECT 1465.750 1945.720 1471.350 1946.570 ;
        RECT 1472.190 1945.720 1474.570 1946.570 ;
        RECT 1475.410 1945.720 1481.010 1946.570 ;
        RECT 1481.850 1945.720 1487.450 1946.570 ;
        RECT 1488.290 1945.720 1493.890 1946.570 ;
        RECT 1494.730 1945.720 1500.330 1946.570 ;
        RECT 1501.170 1945.720 1506.770 1946.570 ;
        RECT 1507.610 1945.720 1513.210 1946.570 ;
        RECT 1514.050 1945.720 1519.650 1946.570 ;
        RECT 1520.490 1945.720 1526.090 1946.570 ;
        RECT 1526.930 1945.720 1532.530 1946.570 ;
        RECT 1533.370 1945.720 1538.970 1946.570 ;
        RECT 1539.810 1945.720 1545.410 1946.570 ;
        RECT 1546.250 1945.720 1551.850 1946.570 ;
        RECT 1552.690 1945.720 1558.290 1946.570 ;
        RECT 1559.130 1945.720 1564.730 1946.570 ;
        RECT 1565.570 1945.720 1571.170 1946.570 ;
        RECT 1572.010 1945.720 1577.610 1946.570 ;
        RECT 1578.450 1945.720 1584.050 1946.570 ;
        RECT 1584.890 1945.720 1590.490 1946.570 ;
        RECT 1591.330 1945.720 1596.930 1946.570 ;
        RECT 1597.770 1945.720 1603.370 1946.570 ;
        RECT 1604.210 1945.720 1609.810 1946.570 ;
        RECT 1610.650 1945.720 1616.250 1946.570 ;
        RECT 1617.090 1945.720 1622.690 1946.570 ;
        RECT 1623.530 1945.720 1629.130 1946.570 ;
        RECT 1629.970 1945.720 1635.570 1946.570 ;
        RECT 1636.410 1945.720 1642.010 1946.570 ;
        RECT 1642.850 1945.720 1648.450 1946.570 ;
        RECT 1649.290 1945.720 1654.890 1946.570 ;
        RECT 1655.730 1945.720 1661.330 1946.570 ;
        RECT 1662.170 1945.720 1667.770 1946.570 ;
        RECT 1668.610 1945.720 1674.210 1946.570 ;
        RECT 1675.050 1945.720 1680.650 1946.570 ;
        RECT 1681.490 1945.720 1687.090 1946.570 ;
        RECT 1687.930 1945.720 1693.530 1946.570 ;
        RECT 1694.370 1945.720 1699.970 1946.570 ;
        RECT 1700.810 1945.720 1706.410 1946.570 ;
        RECT 1707.250 1945.720 1712.850 1946.570 ;
        RECT 1713.690 1945.720 1719.290 1946.570 ;
        RECT 1720.130 1945.720 1725.730 1946.570 ;
        RECT 1726.570 1945.720 1732.170 1946.570 ;
        RECT 1733.010 1945.720 1738.610 1946.570 ;
        RECT 1739.450 1945.720 1745.050 1946.570 ;
        RECT 1745.890 1945.720 1751.490 1946.570 ;
        RECT 1752.330 1945.720 1757.930 1946.570 ;
        RECT 1758.770 1945.720 1764.370 1946.570 ;
        RECT 1765.210 1945.720 1770.810 1946.570 ;
        RECT 1771.650 1945.720 1777.250 1946.570 ;
        RECT 1778.090 1945.720 1783.690 1946.570 ;
        RECT 1784.530 1945.720 1790.130 1946.570 ;
        RECT 1790.970 1945.720 1796.570 1946.570 ;
        RECT 1797.410 1945.720 1803.010 1946.570 ;
        RECT 1803.850 1945.720 1809.450 1946.570 ;
        RECT 1810.290 1945.720 1815.890 1946.570 ;
        RECT 1816.730 1945.720 1822.330 1946.570 ;
        RECT 1823.170 1945.720 1828.770 1946.570 ;
        RECT 1829.610 1945.720 1835.210 1946.570 ;
        RECT 1836.050 1945.720 1841.650 1946.570 ;
        RECT 1842.490 1945.720 1848.090 1946.570 ;
        RECT 1848.930 1945.720 1854.530 1946.570 ;
        RECT 1855.370 1945.720 1860.970 1946.570 ;
        RECT 1861.810 1945.720 1867.410 1946.570 ;
        RECT 1868.250 1945.720 1873.850 1946.570 ;
        RECT 1874.690 1945.720 1880.290 1946.570 ;
        RECT 1881.130 1945.720 1886.730 1946.570 ;
        RECT 1887.570 1945.720 1893.170 1946.570 ;
        RECT 1894.010 1945.720 1899.610 1946.570 ;
        RECT 1900.450 1945.720 1906.050 1946.570 ;
        RECT 1906.890 1945.720 1912.490 1946.570 ;
        RECT 1913.330 1945.720 1918.930 1946.570 ;
        RECT 1919.770 1945.720 1925.370 1946.570 ;
        RECT 1926.210 1945.720 1931.810 1946.570 ;
        RECT 1932.650 1945.720 1938.250 1946.570 ;
        RECT 1939.090 1945.720 1944.690 1946.570 ;
        RECT 1945.530 1945.720 1947.910 1946.570 ;
        RECT 0.100 4.280 1948.460 1945.720 ;
        RECT 0.650 3.670 3.030 4.280 ;
        RECT 3.870 3.670 9.470 4.280 ;
        RECT 10.310 3.670 15.910 4.280 ;
        RECT 16.750 3.670 22.350 4.280 ;
        RECT 23.190 3.670 28.790 4.280 ;
        RECT 29.630 3.670 35.230 4.280 ;
        RECT 36.070 3.670 41.670 4.280 ;
        RECT 42.510 3.670 48.110 4.280 ;
        RECT 48.950 3.670 54.550 4.280 ;
        RECT 55.390 3.670 60.990 4.280 ;
        RECT 61.830 3.670 67.430 4.280 ;
        RECT 68.270 3.670 73.870 4.280 ;
        RECT 74.710 3.670 80.310 4.280 ;
        RECT 81.150 3.670 86.750 4.280 ;
        RECT 87.590 3.670 93.190 4.280 ;
        RECT 94.030 3.670 99.630 4.280 ;
        RECT 100.470 3.670 106.070 4.280 ;
        RECT 106.910 3.670 112.510 4.280 ;
        RECT 113.350 3.670 118.950 4.280 ;
        RECT 119.790 3.670 125.390 4.280 ;
        RECT 126.230 3.670 131.830 4.280 ;
        RECT 132.670 3.670 138.270 4.280 ;
        RECT 139.110 3.670 144.710 4.280 ;
        RECT 145.550 3.670 151.150 4.280 ;
        RECT 151.990 3.670 157.590 4.280 ;
        RECT 158.430 3.670 164.030 4.280 ;
        RECT 164.870 3.670 170.470 4.280 ;
        RECT 171.310 3.670 176.910 4.280 ;
        RECT 177.750 3.670 183.350 4.280 ;
        RECT 184.190 3.670 189.790 4.280 ;
        RECT 190.630 3.670 196.230 4.280 ;
        RECT 197.070 3.670 202.670 4.280 ;
        RECT 203.510 3.670 209.110 4.280 ;
        RECT 209.950 3.670 215.550 4.280 ;
        RECT 216.390 3.670 221.990 4.280 ;
        RECT 222.830 3.670 228.430 4.280 ;
        RECT 229.270 3.670 234.870 4.280 ;
        RECT 235.710 3.670 241.310 4.280 ;
        RECT 242.150 3.670 247.750 4.280 ;
        RECT 248.590 3.670 254.190 4.280 ;
        RECT 255.030 3.670 260.630 4.280 ;
        RECT 261.470 3.670 267.070 4.280 ;
        RECT 267.910 3.670 273.510 4.280 ;
        RECT 274.350 3.670 279.950 4.280 ;
        RECT 280.790 3.670 286.390 4.280 ;
        RECT 287.230 3.670 292.830 4.280 ;
        RECT 293.670 3.670 299.270 4.280 ;
        RECT 300.110 3.670 305.710 4.280 ;
        RECT 306.550 3.670 312.150 4.280 ;
        RECT 312.990 3.670 318.590 4.280 ;
        RECT 319.430 3.670 325.030 4.280 ;
        RECT 325.870 3.670 331.470 4.280 ;
        RECT 332.310 3.670 337.910 4.280 ;
        RECT 338.750 3.670 344.350 4.280 ;
        RECT 345.190 3.670 350.790 4.280 ;
        RECT 351.630 3.670 357.230 4.280 ;
        RECT 358.070 3.670 363.670 4.280 ;
        RECT 364.510 3.670 370.110 4.280 ;
        RECT 370.950 3.670 376.550 4.280 ;
        RECT 377.390 3.670 382.990 4.280 ;
        RECT 383.830 3.670 389.430 4.280 ;
        RECT 390.270 3.670 395.870 4.280 ;
        RECT 396.710 3.670 402.310 4.280 ;
        RECT 403.150 3.670 408.750 4.280 ;
        RECT 409.590 3.670 415.190 4.280 ;
        RECT 416.030 3.670 421.630 4.280 ;
        RECT 422.470 3.670 428.070 4.280 ;
        RECT 428.910 3.670 434.510 4.280 ;
        RECT 435.350 3.670 440.950 4.280 ;
        RECT 441.790 3.670 447.390 4.280 ;
        RECT 448.230 3.670 453.830 4.280 ;
        RECT 454.670 3.670 460.270 4.280 ;
        RECT 461.110 3.670 466.710 4.280 ;
        RECT 467.550 3.670 473.150 4.280 ;
        RECT 473.990 3.670 476.370 4.280 ;
        RECT 477.210 3.670 482.810 4.280 ;
        RECT 483.650 3.670 489.250 4.280 ;
        RECT 490.090 3.670 495.690 4.280 ;
        RECT 496.530 3.670 502.130 4.280 ;
        RECT 502.970 3.670 508.570 4.280 ;
        RECT 509.410 3.670 515.010 4.280 ;
        RECT 515.850 3.670 521.450 4.280 ;
        RECT 522.290 3.670 527.890 4.280 ;
        RECT 528.730 3.670 534.330 4.280 ;
        RECT 535.170 3.670 540.770 4.280 ;
        RECT 541.610 3.670 547.210 4.280 ;
        RECT 548.050 3.670 553.650 4.280 ;
        RECT 554.490 3.670 560.090 4.280 ;
        RECT 560.930 3.670 566.530 4.280 ;
        RECT 567.370 3.670 572.970 4.280 ;
        RECT 573.810 3.670 579.410 4.280 ;
        RECT 580.250 3.670 585.850 4.280 ;
        RECT 586.690 3.670 592.290 4.280 ;
        RECT 593.130 3.670 598.730 4.280 ;
        RECT 599.570 3.670 605.170 4.280 ;
        RECT 606.010 3.670 611.610 4.280 ;
        RECT 612.450 3.670 618.050 4.280 ;
        RECT 618.890 3.670 624.490 4.280 ;
        RECT 625.330 3.670 630.930 4.280 ;
        RECT 631.770 3.670 637.370 4.280 ;
        RECT 638.210 3.670 643.810 4.280 ;
        RECT 644.650 3.670 650.250 4.280 ;
        RECT 651.090 3.670 656.690 4.280 ;
        RECT 657.530 3.670 663.130 4.280 ;
        RECT 663.970 3.670 669.570 4.280 ;
        RECT 670.410 3.670 676.010 4.280 ;
        RECT 676.850 3.670 682.450 4.280 ;
        RECT 683.290 3.670 688.890 4.280 ;
        RECT 689.730 3.670 695.330 4.280 ;
        RECT 696.170 3.670 701.770 4.280 ;
        RECT 702.610 3.670 708.210 4.280 ;
        RECT 709.050 3.670 714.650 4.280 ;
        RECT 715.490 3.670 721.090 4.280 ;
        RECT 721.930 3.670 727.530 4.280 ;
        RECT 728.370 3.670 733.970 4.280 ;
        RECT 734.810 3.670 740.410 4.280 ;
        RECT 741.250 3.670 746.850 4.280 ;
        RECT 747.690 3.670 753.290 4.280 ;
        RECT 754.130 3.670 759.730 4.280 ;
        RECT 760.570 3.670 766.170 4.280 ;
        RECT 767.010 3.670 772.610 4.280 ;
        RECT 773.450 3.670 779.050 4.280 ;
        RECT 779.890 3.670 785.490 4.280 ;
        RECT 786.330 3.670 791.930 4.280 ;
        RECT 792.770 3.670 798.370 4.280 ;
        RECT 799.210 3.670 804.810 4.280 ;
        RECT 805.650 3.670 811.250 4.280 ;
        RECT 812.090 3.670 817.690 4.280 ;
        RECT 818.530 3.670 824.130 4.280 ;
        RECT 824.970 3.670 830.570 4.280 ;
        RECT 831.410 3.670 837.010 4.280 ;
        RECT 837.850 3.670 843.450 4.280 ;
        RECT 844.290 3.670 849.890 4.280 ;
        RECT 850.730 3.670 856.330 4.280 ;
        RECT 857.170 3.670 862.770 4.280 ;
        RECT 863.610 3.670 869.210 4.280 ;
        RECT 870.050 3.670 875.650 4.280 ;
        RECT 876.490 3.670 882.090 4.280 ;
        RECT 882.930 3.670 888.530 4.280 ;
        RECT 889.370 3.670 894.970 4.280 ;
        RECT 895.810 3.670 901.410 4.280 ;
        RECT 902.250 3.670 907.850 4.280 ;
        RECT 908.690 3.670 914.290 4.280 ;
        RECT 915.130 3.670 920.730 4.280 ;
        RECT 921.570 3.670 927.170 4.280 ;
        RECT 928.010 3.670 933.610 4.280 ;
        RECT 934.450 3.670 940.050 4.280 ;
        RECT 940.890 3.670 946.490 4.280 ;
        RECT 947.330 3.670 949.710 4.280 ;
        RECT 950.550 3.670 956.150 4.280 ;
        RECT 956.990 3.670 962.590 4.280 ;
        RECT 963.430 3.670 969.030 4.280 ;
        RECT 969.870 3.670 975.470 4.280 ;
        RECT 976.310 3.670 981.910 4.280 ;
        RECT 982.750 3.670 988.350 4.280 ;
        RECT 989.190 3.670 994.790 4.280 ;
        RECT 995.630 3.670 1001.230 4.280 ;
        RECT 1002.070 3.670 1007.670 4.280 ;
        RECT 1008.510 3.670 1014.110 4.280 ;
        RECT 1014.950 3.670 1020.550 4.280 ;
        RECT 1021.390 3.670 1026.990 4.280 ;
        RECT 1027.830 3.670 1033.430 4.280 ;
        RECT 1034.270 3.670 1039.870 4.280 ;
        RECT 1040.710 3.670 1046.310 4.280 ;
        RECT 1047.150 3.670 1052.750 4.280 ;
        RECT 1053.590 3.670 1059.190 4.280 ;
        RECT 1060.030 3.670 1065.630 4.280 ;
        RECT 1066.470 3.670 1072.070 4.280 ;
        RECT 1072.910 3.670 1078.510 4.280 ;
        RECT 1079.350 3.670 1084.950 4.280 ;
        RECT 1085.790 3.670 1091.390 4.280 ;
        RECT 1092.230 3.670 1097.830 4.280 ;
        RECT 1098.670 3.670 1104.270 4.280 ;
        RECT 1105.110 3.670 1110.710 4.280 ;
        RECT 1111.550 3.670 1117.150 4.280 ;
        RECT 1117.990 3.670 1123.590 4.280 ;
        RECT 1124.430 3.670 1130.030 4.280 ;
        RECT 1130.870 3.670 1136.470 4.280 ;
        RECT 1137.310 3.670 1142.910 4.280 ;
        RECT 1143.750 3.670 1149.350 4.280 ;
        RECT 1150.190 3.670 1155.790 4.280 ;
        RECT 1156.630 3.670 1162.230 4.280 ;
        RECT 1163.070 3.670 1168.670 4.280 ;
        RECT 1169.510 3.670 1175.110 4.280 ;
        RECT 1175.950 3.670 1181.550 4.280 ;
        RECT 1182.390 3.670 1187.990 4.280 ;
        RECT 1188.830 3.670 1194.430 4.280 ;
        RECT 1195.270 3.670 1200.870 4.280 ;
        RECT 1201.710 3.670 1207.310 4.280 ;
        RECT 1208.150 3.670 1213.750 4.280 ;
        RECT 1214.590 3.670 1220.190 4.280 ;
        RECT 1221.030 3.670 1226.630 4.280 ;
        RECT 1227.470 3.670 1233.070 4.280 ;
        RECT 1233.910 3.670 1239.510 4.280 ;
        RECT 1240.350 3.670 1245.950 4.280 ;
        RECT 1246.790 3.670 1252.390 4.280 ;
        RECT 1253.230 3.670 1258.830 4.280 ;
        RECT 1259.670 3.670 1265.270 4.280 ;
        RECT 1266.110 3.670 1271.710 4.280 ;
        RECT 1272.550 3.670 1278.150 4.280 ;
        RECT 1278.990 3.670 1284.590 4.280 ;
        RECT 1285.430 3.670 1291.030 4.280 ;
        RECT 1291.870 3.670 1297.470 4.280 ;
        RECT 1298.310 3.670 1303.910 4.280 ;
        RECT 1304.750 3.670 1310.350 4.280 ;
        RECT 1311.190 3.670 1316.790 4.280 ;
        RECT 1317.630 3.670 1323.230 4.280 ;
        RECT 1324.070 3.670 1329.670 4.280 ;
        RECT 1330.510 3.670 1336.110 4.280 ;
        RECT 1336.950 3.670 1342.550 4.280 ;
        RECT 1343.390 3.670 1348.990 4.280 ;
        RECT 1349.830 3.670 1355.430 4.280 ;
        RECT 1356.270 3.670 1361.870 4.280 ;
        RECT 1362.710 3.670 1368.310 4.280 ;
        RECT 1369.150 3.670 1374.750 4.280 ;
        RECT 1375.590 3.670 1381.190 4.280 ;
        RECT 1382.030 3.670 1387.630 4.280 ;
        RECT 1388.470 3.670 1394.070 4.280 ;
        RECT 1394.910 3.670 1400.510 4.280 ;
        RECT 1401.350 3.670 1406.950 4.280 ;
        RECT 1407.790 3.670 1413.390 4.280 ;
        RECT 1414.230 3.670 1419.830 4.280 ;
        RECT 1420.670 3.670 1423.050 4.280 ;
        RECT 1423.890 3.670 1429.490 4.280 ;
        RECT 1430.330 3.670 1435.930 4.280 ;
        RECT 1436.770 3.670 1442.370 4.280 ;
        RECT 1443.210 3.670 1448.810 4.280 ;
        RECT 1449.650 3.670 1455.250 4.280 ;
        RECT 1456.090 3.670 1461.690 4.280 ;
        RECT 1462.530 3.670 1468.130 4.280 ;
        RECT 1468.970 3.670 1474.570 4.280 ;
        RECT 1475.410 3.670 1481.010 4.280 ;
        RECT 1481.850 3.670 1487.450 4.280 ;
        RECT 1488.290 3.670 1493.890 4.280 ;
        RECT 1494.730 3.670 1500.330 4.280 ;
        RECT 1501.170 3.670 1506.770 4.280 ;
        RECT 1507.610 3.670 1513.210 4.280 ;
        RECT 1514.050 3.670 1519.650 4.280 ;
        RECT 1520.490 3.670 1526.090 4.280 ;
        RECT 1526.930 3.670 1532.530 4.280 ;
        RECT 1533.370 3.670 1538.970 4.280 ;
        RECT 1539.810 3.670 1545.410 4.280 ;
        RECT 1546.250 3.670 1551.850 4.280 ;
        RECT 1552.690 3.670 1558.290 4.280 ;
        RECT 1559.130 3.670 1564.730 4.280 ;
        RECT 1565.570 3.670 1571.170 4.280 ;
        RECT 1572.010 3.670 1577.610 4.280 ;
        RECT 1578.450 3.670 1584.050 4.280 ;
        RECT 1584.890 3.670 1590.490 4.280 ;
        RECT 1591.330 3.670 1596.930 4.280 ;
        RECT 1597.770 3.670 1603.370 4.280 ;
        RECT 1604.210 3.670 1609.810 4.280 ;
        RECT 1610.650 3.670 1616.250 4.280 ;
        RECT 1617.090 3.670 1622.690 4.280 ;
        RECT 1623.530 3.670 1629.130 4.280 ;
        RECT 1629.970 3.670 1635.570 4.280 ;
        RECT 1636.410 3.670 1642.010 4.280 ;
        RECT 1642.850 3.670 1648.450 4.280 ;
        RECT 1649.290 3.670 1654.890 4.280 ;
        RECT 1655.730 3.670 1661.330 4.280 ;
        RECT 1662.170 3.670 1667.770 4.280 ;
        RECT 1668.610 3.670 1674.210 4.280 ;
        RECT 1675.050 3.670 1680.650 4.280 ;
        RECT 1681.490 3.670 1687.090 4.280 ;
        RECT 1687.930 3.670 1693.530 4.280 ;
        RECT 1694.370 3.670 1699.970 4.280 ;
        RECT 1700.810 3.670 1706.410 4.280 ;
        RECT 1707.250 3.670 1712.850 4.280 ;
        RECT 1713.690 3.670 1719.290 4.280 ;
        RECT 1720.130 3.670 1725.730 4.280 ;
        RECT 1726.570 3.670 1732.170 4.280 ;
        RECT 1733.010 3.670 1738.610 4.280 ;
        RECT 1739.450 3.670 1745.050 4.280 ;
        RECT 1745.890 3.670 1751.490 4.280 ;
        RECT 1752.330 3.670 1757.930 4.280 ;
        RECT 1758.770 3.670 1764.370 4.280 ;
        RECT 1765.210 3.670 1770.810 4.280 ;
        RECT 1771.650 3.670 1777.250 4.280 ;
        RECT 1778.090 3.670 1783.690 4.280 ;
        RECT 1784.530 3.670 1790.130 4.280 ;
        RECT 1790.970 3.670 1796.570 4.280 ;
        RECT 1797.410 3.670 1803.010 4.280 ;
        RECT 1803.850 3.670 1809.450 4.280 ;
        RECT 1810.290 3.670 1815.890 4.280 ;
        RECT 1816.730 3.670 1822.330 4.280 ;
        RECT 1823.170 3.670 1828.770 4.280 ;
        RECT 1829.610 3.670 1835.210 4.280 ;
        RECT 1836.050 3.670 1841.650 4.280 ;
        RECT 1842.490 3.670 1848.090 4.280 ;
        RECT 1848.930 3.670 1854.530 4.280 ;
        RECT 1855.370 3.670 1860.970 4.280 ;
        RECT 1861.810 3.670 1867.410 4.280 ;
        RECT 1868.250 3.670 1873.850 4.280 ;
        RECT 1874.690 3.670 1880.290 4.280 ;
        RECT 1881.130 3.670 1886.730 4.280 ;
        RECT 1887.570 3.670 1893.170 4.280 ;
        RECT 1894.010 3.670 1899.610 4.280 ;
        RECT 1900.450 3.670 1902.830 4.280 ;
        RECT 1903.670 3.670 1909.270 4.280 ;
        RECT 1910.110 3.670 1915.710 4.280 ;
        RECT 1916.550 3.670 1922.150 4.280 ;
        RECT 1922.990 3.670 1928.590 4.280 ;
        RECT 1929.430 3.670 1935.030 4.280 ;
        RECT 1935.870 3.670 1941.470 4.280 ;
        RECT 1942.310 3.670 1947.910 4.280 ;
      LAYER met3 ;
        RECT 4.400 1944.440 1945.600 1945.305 ;
        RECT 4.000 1939.040 1946.000 1944.440 ;
        RECT 4.400 1937.640 1945.600 1939.040 ;
        RECT 4.000 1932.240 1946.000 1937.640 ;
        RECT 4.400 1930.840 1945.600 1932.240 ;
        RECT 4.000 1925.440 1946.000 1930.840 ;
        RECT 4.400 1924.040 1945.600 1925.440 ;
        RECT 4.000 1918.640 1946.000 1924.040 ;
        RECT 4.400 1917.240 1945.600 1918.640 ;
        RECT 4.000 1911.840 1946.000 1917.240 ;
        RECT 4.400 1910.440 1945.600 1911.840 ;
        RECT 4.000 1905.040 1946.000 1910.440 ;
        RECT 4.400 1903.640 1945.600 1905.040 ;
        RECT 4.000 1898.240 1946.000 1903.640 ;
        RECT 4.400 1896.840 1945.600 1898.240 ;
        RECT 4.000 1891.440 1946.000 1896.840 ;
        RECT 4.400 1890.040 1945.600 1891.440 ;
        RECT 4.000 1884.640 1946.000 1890.040 ;
        RECT 4.400 1883.240 1945.600 1884.640 ;
        RECT 4.000 1877.840 1946.000 1883.240 ;
        RECT 4.400 1876.440 1945.600 1877.840 ;
        RECT 4.000 1871.040 1946.000 1876.440 ;
        RECT 4.400 1869.640 1945.600 1871.040 ;
        RECT 4.000 1864.240 1946.000 1869.640 ;
        RECT 4.400 1862.840 1945.600 1864.240 ;
        RECT 4.000 1857.440 1946.000 1862.840 ;
        RECT 4.400 1856.040 1945.600 1857.440 ;
        RECT 4.000 1850.640 1946.000 1856.040 ;
        RECT 4.400 1849.240 1945.600 1850.640 ;
        RECT 4.000 1843.840 1946.000 1849.240 ;
        RECT 4.400 1842.440 1945.600 1843.840 ;
        RECT 4.000 1837.040 1946.000 1842.440 ;
        RECT 4.400 1835.640 1945.600 1837.040 ;
        RECT 4.000 1830.240 1946.000 1835.640 ;
        RECT 4.400 1828.840 1945.600 1830.240 ;
        RECT 4.000 1823.440 1946.000 1828.840 ;
        RECT 4.400 1822.040 1945.600 1823.440 ;
        RECT 4.000 1816.640 1946.000 1822.040 ;
        RECT 4.400 1815.240 1945.600 1816.640 ;
        RECT 4.000 1809.840 1946.000 1815.240 ;
        RECT 4.400 1808.440 1945.600 1809.840 ;
        RECT 4.000 1803.040 1946.000 1808.440 ;
        RECT 4.400 1801.640 1945.600 1803.040 ;
        RECT 4.000 1796.240 1946.000 1801.640 ;
        RECT 4.400 1794.840 1945.600 1796.240 ;
        RECT 4.000 1789.440 1946.000 1794.840 ;
        RECT 4.400 1788.040 1945.600 1789.440 ;
        RECT 4.000 1782.640 1946.000 1788.040 ;
        RECT 4.400 1781.240 1945.600 1782.640 ;
        RECT 4.000 1775.840 1946.000 1781.240 ;
        RECT 4.400 1774.440 1945.600 1775.840 ;
        RECT 4.000 1769.040 1946.000 1774.440 ;
        RECT 4.400 1767.640 1945.600 1769.040 ;
        RECT 4.000 1762.240 1946.000 1767.640 ;
        RECT 4.400 1760.840 1945.600 1762.240 ;
        RECT 4.000 1755.440 1946.000 1760.840 ;
        RECT 4.400 1754.040 1945.600 1755.440 ;
        RECT 4.000 1748.640 1946.000 1754.040 ;
        RECT 4.400 1747.240 1945.600 1748.640 ;
        RECT 4.000 1741.840 1946.000 1747.240 ;
        RECT 4.400 1740.440 1945.600 1741.840 ;
        RECT 4.000 1735.040 1946.000 1740.440 ;
        RECT 4.400 1733.640 1945.600 1735.040 ;
        RECT 4.000 1728.240 1946.000 1733.640 ;
        RECT 4.400 1726.840 1945.600 1728.240 ;
        RECT 4.000 1721.440 1946.000 1726.840 ;
        RECT 4.400 1720.040 1945.600 1721.440 ;
        RECT 4.000 1714.640 1946.000 1720.040 ;
        RECT 4.400 1713.240 1945.600 1714.640 ;
        RECT 4.000 1707.840 1946.000 1713.240 ;
        RECT 4.400 1706.440 1945.600 1707.840 ;
        RECT 4.000 1701.040 1946.000 1706.440 ;
        RECT 4.400 1699.640 1945.600 1701.040 ;
        RECT 4.000 1694.240 1946.000 1699.640 ;
        RECT 4.400 1692.840 1945.600 1694.240 ;
        RECT 4.000 1687.440 1946.000 1692.840 ;
        RECT 4.400 1686.040 1945.600 1687.440 ;
        RECT 4.000 1680.640 1946.000 1686.040 ;
        RECT 4.400 1679.240 1945.600 1680.640 ;
        RECT 4.000 1673.840 1946.000 1679.240 ;
        RECT 4.400 1672.440 1945.600 1673.840 ;
        RECT 4.000 1667.040 1946.000 1672.440 ;
        RECT 4.400 1665.640 1945.600 1667.040 ;
        RECT 4.000 1660.240 1946.000 1665.640 ;
        RECT 4.400 1658.840 1945.600 1660.240 ;
        RECT 4.000 1653.440 1946.000 1658.840 ;
        RECT 4.400 1652.040 1945.600 1653.440 ;
        RECT 4.000 1646.640 1946.000 1652.040 ;
        RECT 4.400 1645.240 1945.600 1646.640 ;
        RECT 4.000 1639.840 1946.000 1645.240 ;
        RECT 4.400 1638.440 1945.600 1639.840 ;
        RECT 4.000 1633.040 1946.000 1638.440 ;
        RECT 4.400 1631.640 1945.600 1633.040 ;
        RECT 4.000 1626.240 1946.000 1631.640 ;
        RECT 4.400 1624.840 1945.600 1626.240 ;
        RECT 4.000 1619.440 1946.000 1624.840 ;
        RECT 4.400 1618.040 1945.600 1619.440 ;
        RECT 4.000 1612.640 1946.000 1618.040 ;
        RECT 4.400 1611.240 1945.600 1612.640 ;
        RECT 4.000 1605.840 1946.000 1611.240 ;
        RECT 4.400 1604.440 1945.600 1605.840 ;
        RECT 4.000 1599.040 1946.000 1604.440 ;
        RECT 4.400 1597.640 1945.600 1599.040 ;
        RECT 4.000 1592.240 1946.000 1597.640 ;
        RECT 4.400 1590.840 1945.600 1592.240 ;
        RECT 4.000 1585.440 1946.000 1590.840 ;
        RECT 4.400 1584.040 1945.600 1585.440 ;
        RECT 4.000 1578.640 1946.000 1584.040 ;
        RECT 4.400 1577.240 1945.600 1578.640 ;
        RECT 4.000 1571.840 1946.000 1577.240 ;
        RECT 4.400 1570.440 1945.600 1571.840 ;
        RECT 4.000 1565.040 1946.000 1570.440 ;
        RECT 4.400 1563.640 1945.600 1565.040 ;
        RECT 4.000 1558.240 1946.000 1563.640 ;
        RECT 4.400 1556.840 1945.600 1558.240 ;
        RECT 4.000 1551.440 1946.000 1556.840 ;
        RECT 4.400 1550.040 1945.600 1551.440 ;
        RECT 4.000 1544.640 1946.000 1550.040 ;
        RECT 4.400 1543.240 1945.600 1544.640 ;
        RECT 4.000 1537.840 1946.000 1543.240 ;
        RECT 4.400 1536.440 1945.600 1537.840 ;
        RECT 4.000 1531.040 1946.000 1536.440 ;
        RECT 4.400 1529.640 1945.600 1531.040 ;
        RECT 4.000 1524.240 1946.000 1529.640 ;
        RECT 4.400 1522.840 1945.600 1524.240 ;
        RECT 4.000 1517.440 1946.000 1522.840 ;
        RECT 4.400 1516.040 1945.600 1517.440 ;
        RECT 4.000 1510.640 1946.000 1516.040 ;
        RECT 4.400 1509.240 1945.600 1510.640 ;
        RECT 4.000 1503.840 1946.000 1509.240 ;
        RECT 4.400 1502.440 1945.600 1503.840 ;
        RECT 4.000 1500.440 1946.000 1502.440 ;
        RECT 4.400 1499.040 1946.000 1500.440 ;
        RECT 4.000 1497.040 1946.000 1499.040 ;
        RECT 4.000 1495.640 1945.600 1497.040 ;
        RECT 4.000 1493.640 1946.000 1495.640 ;
        RECT 4.400 1492.240 1946.000 1493.640 ;
        RECT 4.000 1490.240 1946.000 1492.240 ;
        RECT 4.000 1488.840 1945.600 1490.240 ;
        RECT 4.000 1486.840 1946.000 1488.840 ;
        RECT 4.400 1485.440 1946.000 1486.840 ;
        RECT 4.000 1483.440 1946.000 1485.440 ;
        RECT 4.000 1482.040 1945.600 1483.440 ;
        RECT 4.000 1480.040 1946.000 1482.040 ;
        RECT 4.400 1478.640 1946.000 1480.040 ;
        RECT 4.000 1476.640 1946.000 1478.640 ;
        RECT 4.000 1475.240 1945.600 1476.640 ;
        RECT 4.000 1473.240 1946.000 1475.240 ;
        RECT 4.400 1471.840 1946.000 1473.240 ;
        RECT 4.000 1469.840 1946.000 1471.840 ;
        RECT 4.000 1468.440 1945.600 1469.840 ;
        RECT 4.000 1466.440 1946.000 1468.440 ;
        RECT 4.400 1465.040 1946.000 1466.440 ;
        RECT 4.000 1463.040 1946.000 1465.040 ;
        RECT 4.000 1461.640 1945.600 1463.040 ;
        RECT 4.000 1459.640 1946.000 1461.640 ;
        RECT 4.400 1458.240 1946.000 1459.640 ;
        RECT 4.000 1456.240 1946.000 1458.240 ;
        RECT 4.000 1454.840 1945.600 1456.240 ;
        RECT 4.000 1452.840 1946.000 1454.840 ;
        RECT 4.400 1451.440 1946.000 1452.840 ;
        RECT 4.000 1449.440 1946.000 1451.440 ;
        RECT 4.000 1448.040 1945.600 1449.440 ;
        RECT 4.000 1446.040 1946.000 1448.040 ;
        RECT 4.400 1444.640 1945.600 1446.040 ;
        RECT 4.000 1439.240 1946.000 1444.640 ;
        RECT 4.400 1437.840 1945.600 1439.240 ;
        RECT 4.000 1432.440 1946.000 1437.840 ;
        RECT 4.400 1431.040 1945.600 1432.440 ;
        RECT 4.000 1425.640 1946.000 1431.040 ;
        RECT 4.400 1424.240 1945.600 1425.640 ;
        RECT 4.000 1418.840 1946.000 1424.240 ;
        RECT 4.400 1417.440 1945.600 1418.840 ;
        RECT 4.000 1412.040 1946.000 1417.440 ;
        RECT 4.400 1410.640 1945.600 1412.040 ;
        RECT 4.000 1405.240 1946.000 1410.640 ;
        RECT 4.400 1403.840 1945.600 1405.240 ;
        RECT 4.000 1398.440 1946.000 1403.840 ;
        RECT 4.400 1397.040 1945.600 1398.440 ;
        RECT 4.000 1391.640 1946.000 1397.040 ;
        RECT 4.400 1390.240 1945.600 1391.640 ;
        RECT 4.000 1384.840 1946.000 1390.240 ;
        RECT 4.400 1383.440 1945.600 1384.840 ;
        RECT 4.000 1378.040 1946.000 1383.440 ;
        RECT 4.400 1376.640 1945.600 1378.040 ;
        RECT 4.000 1371.240 1946.000 1376.640 ;
        RECT 4.400 1369.840 1945.600 1371.240 ;
        RECT 4.000 1364.440 1946.000 1369.840 ;
        RECT 4.400 1363.040 1945.600 1364.440 ;
        RECT 4.000 1357.640 1946.000 1363.040 ;
        RECT 4.400 1356.240 1945.600 1357.640 ;
        RECT 4.000 1350.840 1946.000 1356.240 ;
        RECT 4.400 1349.440 1945.600 1350.840 ;
        RECT 4.000 1344.040 1946.000 1349.440 ;
        RECT 4.400 1342.640 1945.600 1344.040 ;
        RECT 4.000 1337.240 1946.000 1342.640 ;
        RECT 4.400 1335.840 1945.600 1337.240 ;
        RECT 4.000 1330.440 1946.000 1335.840 ;
        RECT 4.400 1329.040 1945.600 1330.440 ;
        RECT 4.000 1323.640 1946.000 1329.040 ;
        RECT 4.400 1322.240 1945.600 1323.640 ;
        RECT 4.000 1316.840 1946.000 1322.240 ;
        RECT 4.400 1315.440 1945.600 1316.840 ;
        RECT 4.000 1310.040 1946.000 1315.440 ;
        RECT 4.400 1308.640 1945.600 1310.040 ;
        RECT 4.000 1303.240 1946.000 1308.640 ;
        RECT 4.400 1301.840 1945.600 1303.240 ;
        RECT 4.000 1296.440 1946.000 1301.840 ;
        RECT 4.400 1295.040 1945.600 1296.440 ;
        RECT 4.000 1289.640 1946.000 1295.040 ;
        RECT 4.400 1288.240 1945.600 1289.640 ;
        RECT 4.000 1282.840 1946.000 1288.240 ;
        RECT 4.400 1281.440 1945.600 1282.840 ;
        RECT 4.000 1276.040 1946.000 1281.440 ;
        RECT 4.400 1274.640 1945.600 1276.040 ;
        RECT 4.000 1269.240 1946.000 1274.640 ;
        RECT 4.400 1267.840 1945.600 1269.240 ;
        RECT 4.000 1262.440 1946.000 1267.840 ;
        RECT 4.400 1261.040 1945.600 1262.440 ;
        RECT 4.000 1255.640 1946.000 1261.040 ;
        RECT 4.400 1254.240 1945.600 1255.640 ;
        RECT 4.000 1248.840 1946.000 1254.240 ;
        RECT 4.400 1247.440 1945.600 1248.840 ;
        RECT 4.000 1242.040 1946.000 1247.440 ;
        RECT 4.400 1240.640 1945.600 1242.040 ;
        RECT 4.000 1235.240 1946.000 1240.640 ;
        RECT 4.400 1233.840 1945.600 1235.240 ;
        RECT 4.000 1228.440 1946.000 1233.840 ;
        RECT 4.400 1227.040 1945.600 1228.440 ;
        RECT 4.000 1221.640 1946.000 1227.040 ;
        RECT 4.400 1220.240 1945.600 1221.640 ;
        RECT 4.000 1214.840 1946.000 1220.240 ;
        RECT 4.400 1213.440 1945.600 1214.840 ;
        RECT 4.000 1208.040 1946.000 1213.440 ;
        RECT 4.400 1206.640 1945.600 1208.040 ;
        RECT 4.000 1201.240 1946.000 1206.640 ;
        RECT 4.400 1199.840 1945.600 1201.240 ;
        RECT 4.000 1194.440 1946.000 1199.840 ;
        RECT 4.400 1193.040 1945.600 1194.440 ;
        RECT 4.000 1187.640 1946.000 1193.040 ;
        RECT 4.400 1186.240 1945.600 1187.640 ;
        RECT 4.000 1180.840 1946.000 1186.240 ;
        RECT 4.400 1179.440 1945.600 1180.840 ;
        RECT 4.000 1174.040 1946.000 1179.440 ;
        RECT 4.400 1172.640 1945.600 1174.040 ;
        RECT 4.000 1167.240 1946.000 1172.640 ;
        RECT 4.400 1165.840 1945.600 1167.240 ;
        RECT 4.000 1160.440 1946.000 1165.840 ;
        RECT 4.400 1159.040 1945.600 1160.440 ;
        RECT 4.000 1153.640 1946.000 1159.040 ;
        RECT 4.400 1152.240 1945.600 1153.640 ;
        RECT 4.000 1146.840 1946.000 1152.240 ;
        RECT 4.400 1145.440 1945.600 1146.840 ;
        RECT 4.000 1140.040 1946.000 1145.440 ;
        RECT 4.400 1138.640 1945.600 1140.040 ;
        RECT 4.000 1133.240 1946.000 1138.640 ;
        RECT 4.400 1131.840 1945.600 1133.240 ;
        RECT 4.000 1126.440 1946.000 1131.840 ;
        RECT 4.400 1125.040 1945.600 1126.440 ;
        RECT 4.000 1119.640 1946.000 1125.040 ;
        RECT 4.400 1118.240 1945.600 1119.640 ;
        RECT 4.000 1112.840 1946.000 1118.240 ;
        RECT 4.400 1111.440 1945.600 1112.840 ;
        RECT 4.000 1106.040 1946.000 1111.440 ;
        RECT 4.400 1104.640 1945.600 1106.040 ;
        RECT 4.000 1099.240 1946.000 1104.640 ;
        RECT 4.400 1097.840 1945.600 1099.240 ;
        RECT 4.000 1092.440 1946.000 1097.840 ;
        RECT 4.400 1091.040 1945.600 1092.440 ;
        RECT 4.000 1085.640 1946.000 1091.040 ;
        RECT 4.400 1084.240 1945.600 1085.640 ;
        RECT 4.000 1078.840 1946.000 1084.240 ;
        RECT 4.400 1077.440 1945.600 1078.840 ;
        RECT 4.000 1072.040 1946.000 1077.440 ;
        RECT 4.400 1070.640 1945.600 1072.040 ;
        RECT 4.000 1065.240 1946.000 1070.640 ;
        RECT 4.400 1063.840 1945.600 1065.240 ;
        RECT 4.000 1058.440 1946.000 1063.840 ;
        RECT 4.400 1057.040 1945.600 1058.440 ;
        RECT 4.000 1051.640 1946.000 1057.040 ;
        RECT 4.400 1050.240 1945.600 1051.640 ;
        RECT 4.000 1044.840 1946.000 1050.240 ;
        RECT 4.400 1043.440 1945.600 1044.840 ;
        RECT 4.000 1038.040 1946.000 1043.440 ;
        RECT 4.400 1036.640 1945.600 1038.040 ;
        RECT 4.000 1031.240 1946.000 1036.640 ;
        RECT 4.400 1029.840 1945.600 1031.240 ;
        RECT 4.000 1024.440 1946.000 1029.840 ;
        RECT 4.400 1023.040 1945.600 1024.440 ;
        RECT 4.000 1017.640 1946.000 1023.040 ;
        RECT 4.400 1016.240 1945.600 1017.640 ;
        RECT 4.000 1010.840 1946.000 1016.240 ;
        RECT 4.400 1009.440 1945.600 1010.840 ;
        RECT 4.000 1004.040 1946.000 1009.440 ;
        RECT 4.400 1002.640 1945.600 1004.040 ;
        RECT 4.000 1000.640 1946.000 1002.640 ;
        RECT 4.400 999.240 1946.000 1000.640 ;
        RECT 4.000 997.240 1946.000 999.240 ;
        RECT 4.000 995.840 1945.600 997.240 ;
        RECT 4.000 993.840 1946.000 995.840 ;
        RECT 4.400 992.440 1946.000 993.840 ;
        RECT 4.000 990.440 1946.000 992.440 ;
        RECT 4.000 989.040 1945.600 990.440 ;
        RECT 4.000 987.040 1946.000 989.040 ;
        RECT 4.400 985.640 1946.000 987.040 ;
        RECT 4.000 983.640 1946.000 985.640 ;
        RECT 4.000 982.240 1945.600 983.640 ;
        RECT 4.000 980.240 1946.000 982.240 ;
        RECT 4.400 978.840 1946.000 980.240 ;
        RECT 4.000 976.840 1946.000 978.840 ;
        RECT 4.000 975.440 1945.600 976.840 ;
        RECT 4.000 973.440 1946.000 975.440 ;
        RECT 4.400 972.040 1946.000 973.440 ;
        RECT 4.000 970.040 1946.000 972.040 ;
        RECT 4.000 968.640 1945.600 970.040 ;
        RECT 4.000 966.640 1946.000 968.640 ;
        RECT 4.400 965.240 1946.000 966.640 ;
        RECT 4.000 963.240 1946.000 965.240 ;
        RECT 4.000 961.840 1945.600 963.240 ;
        RECT 4.000 959.840 1946.000 961.840 ;
        RECT 4.400 958.440 1946.000 959.840 ;
        RECT 4.000 956.440 1946.000 958.440 ;
        RECT 4.000 955.040 1945.600 956.440 ;
        RECT 4.000 953.040 1946.000 955.040 ;
        RECT 4.400 951.640 1946.000 953.040 ;
        RECT 4.000 949.640 1946.000 951.640 ;
        RECT 4.000 948.240 1945.600 949.640 ;
        RECT 4.000 946.240 1946.000 948.240 ;
        RECT 4.400 944.840 1945.600 946.240 ;
        RECT 4.000 939.440 1946.000 944.840 ;
        RECT 4.400 938.040 1945.600 939.440 ;
        RECT 4.000 932.640 1946.000 938.040 ;
        RECT 4.400 931.240 1945.600 932.640 ;
        RECT 4.000 925.840 1946.000 931.240 ;
        RECT 4.400 924.440 1945.600 925.840 ;
        RECT 4.000 919.040 1946.000 924.440 ;
        RECT 4.400 917.640 1945.600 919.040 ;
        RECT 4.000 912.240 1946.000 917.640 ;
        RECT 4.400 910.840 1945.600 912.240 ;
        RECT 4.000 905.440 1946.000 910.840 ;
        RECT 4.400 904.040 1945.600 905.440 ;
        RECT 4.000 898.640 1946.000 904.040 ;
        RECT 4.400 897.240 1945.600 898.640 ;
        RECT 4.000 891.840 1946.000 897.240 ;
        RECT 4.400 890.440 1945.600 891.840 ;
        RECT 4.000 885.040 1946.000 890.440 ;
        RECT 4.400 883.640 1945.600 885.040 ;
        RECT 4.000 878.240 1946.000 883.640 ;
        RECT 4.400 876.840 1945.600 878.240 ;
        RECT 4.000 871.440 1946.000 876.840 ;
        RECT 4.400 870.040 1945.600 871.440 ;
        RECT 4.000 864.640 1946.000 870.040 ;
        RECT 4.400 863.240 1945.600 864.640 ;
        RECT 4.000 857.840 1946.000 863.240 ;
        RECT 4.400 856.440 1945.600 857.840 ;
        RECT 4.000 851.040 1946.000 856.440 ;
        RECT 4.400 849.640 1945.600 851.040 ;
        RECT 4.000 844.240 1946.000 849.640 ;
        RECT 4.400 842.840 1945.600 844.240 ;
        RECT 4.000 837.440 1946.000 842.840 ;
        RECT 4.400 836.040 1945.600 837.440 ;
        RECT 4.000 830.640 1946.000 836.040 ;
        RECT 4.400 829.240 1945.600 830.640 ;
        RECT 4.000 823.840 1946.000 829.240 ;
        RECT 4.400 822.440 1945.600 823.840 ;
        RECT 4.000 817.040 1946.000 822.440 ;
        RECT 4.400 815.640 1945.600 817.040 ;
        RECT 4.000 810.240 1946.000 815.640 ;
        RECT 4.400 808.840 1945.600 810.240 ;
        RECT 4.000 803.440 1946.000 808.840 ;
        RECT 4.400 802.040 1945.600 803.440 ;
        RECT 4.000 796.640 1946.000 802.040 ;
        RECT 4.400 795.240 1945.600 796.640 ;
        RECT 4.000 789.840 1946.000 795.240 ;
        RECT 4.400 788.440 1945.600 789.840 ;
        RECT 4.000 783.040 1946.000 788.440 ;
        RECT 4.400 781.640 1945.600 783.040 ;
        RECT 4.000 776.240 1946.000 781.640 ;
        RECT 4.400 774.840 1945.600 776.240 ;
        RECT 4.000 769.440 1946.000 774.840 ;
        RECT 4.400 768.040 1945.600 769.440 ;
        RECT 4.000 762.640 1946.000 768.040 ;
        RECT 4.400 761.240 1945.600 762.640 ;
        RECT 4.000 755.840 1946.000 761.240 ;
        RECT 4.400 754.440 1945.600 755.840 ;
        RECT 4.000 749.040 1946.000 754.440 ;
        RECT 4.400 747.640 1945.600 749.040 ;
        RECT 4.000 742.240 1946.000 747.640 ;
        RECT 4.400 740.840 1945.600 742.240 ;
        RECT 4.000 735.440 1946.000 740.840 ;
        RECT 4.400 734.040 1945.600 735.440 ;
        RECT 4.000 728.640 1946.000 734.040 ;
        RECT 4.400 727.240 1945.600 728.640 ;
        RECT 4.000 721.840 1946.000 727.240 ;
        RECT 4.400 720.440 1945.600 721.840 ;
        RECT 4.000 715.040 1946.000 720.440 ;
        RECT 4.400 713.640 1945.600 715.040 ;
        RECT 4.000 708.240 1946.000 713.640 ;
        RECT 4.400 706.840 1945.600 708.240 ;
        RECT 4.000 701.440 1946.000 706.840 ;
        RECT 4.400 700.040 1945.600 701.440 ;
        RECT 4.000 694.640 1946.000 700.040 ;
        RECT 4.400 693.240 1945.600 694.640 ;
        RECT 4.000 687.840 1946.000 693.240 ;
        RECT 4.400 686.440 1945.600 687.840 ;
        RECT 4.000 681.040 1946.000 686.440 ;
        RECT 4.400 679.640 1945.600 681.040 ;
        RECT 4.000 674.240 1946.000 679.640 ;
        RECT 4.400 672.840 1945.600 674.240 ;
        RECT 4.000 667.440 1946.000 672.840 ;
        RECT 4.400 666.040 1945.600 667.440 ;
        RECT 4.000 660.640 1946.000 666.040 ;
        RECT 4.400 659.240 1945.600 660.640 ;
        RECT 4.000 653.840 1946.000 659.240 ;
        RECT 4.400 652.440 1945.600 653.840 ;
        RECT 4.000 647.040 1946.000 652.440 ;
        RECT 4.400 645.640 1945.600 647.040 ;
        RECT 4.000 640.240 1946.000 645.640 ;
        RECT 4.400 638.840 1945.600 640.240 ;
        RECT 4.000 633.440 1946.000 638.840 ;
        RECT 4.400 632.040 1945.600 633.440 ;
        RECT 4.000 626.640 1946.000 632.040 ;
        RECT 4.400 625.240 1945.600 626.640 ;
        RECT 4.000 619.840 1946.000 625.240 ;
        RECT 4.400 618.440 1945.600 619.840 ;
        RECT 4.000 613.040 1946.000 618.440 ;
        RECT 4.400 611.640 1945.600 613.040 ;
        RECT 4.000 606.240 1946.000 611.640 ;
        RECT 4.400 604.840 1945.600 606.240 ;
        RECT 4.000 599.440 1946.000 604.840 ;
        RECT 4.400 598.040 1945.600 599.440 ;
        RECT 4.000 592.640 1946.000 598.040 ;
        RECT 4.400 591.240 1945.600 592.640 ;
        RECT 4.000 585.840 1946.000 591.240 ;
        RECT 4.400 584.440 1945.600 585.840 ;
        RECT 4.000 579.040 1946.000 584.440 ;
        RECT 4.400 577.640 1945.600 579.040 ;
        RECT 4.000 572.240 1946.000 577.640 ;
        RECT 4.400 570.840 1945.600 572.240 ;
        RECT 4.000 565.440 1946.000 570.840 ;
        RECT 4.400 564.040 1945.600 565.440 ;
        RECT 4.000 558.640 1946.000 564.040 ;
        RECT 4.400 557.240 1945.600 558.640 ;
        RECT 4.000 551.840 1946.000 557.240 ;
        RECT 4.400 550.440 1945.600 551.840 ;
        RECT 4.000 545.040 1946.000 550.440 ;
        RECT 4.400 543.640 1945.600 545.040 ;
        RECT 4.000 538.240 1946.000 543.640 ;
        RECT 4.400 536.840 1945.600 538.240 ;
        RECT 4.000 531.440 1946.000 536.840 ;
        RECT 4.400 530.040 1945.600 531.440 ;
        RECT 4.000 524.640 1946.000 530.040 ;
        RECT 4.400 523.240 1945.600 524.640 ;
        RECT 4.000 517.840 1946.000 523.240 ;
        RECT 4.400 516.440 1945.600 517.840 ;
        RECT 4.000 511.040 1946.000 516.440 ;
        RECT 4.400 509.640 1945.600 511.040 ;
        RECT 4.000 504.240 1946.000 509.640 ;
        RECT 4.400 502.840 1945.600 504.240 ;
        RECT 4.000 500.840 1946.000 502.840 ;
        RECT 4.400 499.440 1946.000 500.840 ;
        RECT 4.000 497.440 1946.000 499.440 ;
        RECT 4.000 496.040 1945.600 497.440 ;
        RECT 4.000 494.040 1946.000 496.040 ;
        RECT 4.400 492.640 1946.000 494.040 ;
        RECT 4.000 490.640 1946.000 492.640 ;
        RECT 4.000 489.240 1945.600 490.640 ;
        RECT 4.000 487.240 1946.000 489.240 ;
        RECT 4.400 485.840 1946.000 487.240 ;
        RECT 4.000 483.840 1946.000 485.840 ;
        RECT 4.000 482.440 1945.600 483.840 ;
        RECT 4.000 480.440 1946.000 482.440 ;
        RECT 4.400 479.040 1946.000 480.440 ;
        RECT 4.000 477.040 1946.000 479.040 ;
        RECT 4.000 475.640 1945.600 477.040 ;
        RECT 4.000 473.640 1946.000 475.640 ;
        RECT 4.400 472.240 1946.000 473.640 ;
        RECT 4.000 470.240 1946.000 472.240 ;
        RECT 4.000 468.840 1945.600 470.240 ;
        RECT 4.000 466.840 1946.000 468.840 ;
        RECT 4.400 465.440 1946.000 466.840 ;
        RECT 4.000 463.440 1946.000 465.440 ;
        RECT 4.000 462.040 1945.600 463.440 ;
        RECT 4.000 460.040 1946.000 462.040 ;
        RECT 4.400 458.640 1946.000 460.040 ;
        RECT 4.000 456.640 1946.000 458.640 ;
        RECT 4.000 455.240 1945.600 456.640 ;
        RECT 4.000 453.240 1946.000 455.240 ;
        RECT 4.400 451.840 1946.000 453.240 ;
        RECT 4.000 449.840 1946.000 451.840 ;
        RECT 4.000 448.440 1945.600 449.840 ;
        RECT 4.000 446.440 1946.000 448.440 ;
        RECT 4.400 445.040 1945.600 446.440 ;
        RECT 4.000 439.640 1946.000 445.040 ;
        RECT 4.400 438.240 1945.600 439.640 ;
        RECT 4.000 432.840 1946.000 438.240 ;
        RECT 4.400 431.440 1945.600 432.840 ;
        RECT 4.000 426.040 1946.000 431.440 ;
        RECT 4.400 424.640 1945.600 426.040 ;
        RECT 4.000 419.240 1946.000 424.640 ;
        RECT 4.400 417.840 1945.600 419.240 ;
        RECT 4.000 412.440 1946.000 417.840 ;
        RECT 4.400 411.040 1945.600 412.440 ;
        RECT 4.000 405.640 1946.000 411.040 ;
        RECT 4.400 404.240 1945.600 405.640 ;
        RECT 4.000 398.840 1946.000 404.240 ;
        RECT 4.400 397.440 1945.600 398.840 ;
        RECT 4.000 392.040 1946.000 397.440 ;
        RECT 4.400 390.640 1945.600 392.040 ;
        RECT 4.000 385.240 1946.000 390.640 ;
        RECT 4.400 383.840 1945.600 385.240 ;
        RECT 4.000 378.440 1946.000 383.840 ;
        RECT 4.400 377.040 1945.600 378.440 ;
        RECT 4.000 371.640 1946.000 377.040 ;
        RECT 4.400 370.240 1945.600 371.640 ;
        RECT 4.000 364.840 1946.000 370.240 ;
        RECT 4.400 363.440 1945.600 364.840 ;
        RECT 4.000 358.040 1946.000 363.440 ;
        RECT 4.400 356.640 1945.600 358.040 ;
        RECT 4.000 351.240 1946.000 356.640 ;
        RECT 4.400 349.840 1945.600 351.240 ;
        RECT 4.000 344.440 1946.000 349.840 ;
        RECT 4.400 343.040 1945.600 344.440 ;
        RECT 4.000 337.640 1946.000 343.040 ;
        RECT 4.400 336.240 1945.600 337.640 ;
        RECT 4.000 330.840 1946.000 336.240 ;
        RECT 4.400 329.440 1945.600 330.840 ;
        RECT 4.000 324.040 1946.000 329.440 ;
        RECT 4.400 322.640 1945.600 324.040 ;
        RECT 4.000 317.240 1946.000 322.640 ;
        RECT 4.400 315.840 1945.600 317.240 ;
        RECT 4.000 310.440 1946.000 315.840 ;
        RECT 4.400 309.040 1945.600 310.440 ;
        RECT 4.000 303.640 1946.000 309.040 ;
        RECT 4.400 302.240 1945.600 303.640 ;
        RECT 4.000 296.840 1946.000 302.240 ;
        RECT 4.400 295.440 1945.600 296.840 ;
        RECT 4.000 290.040 1946.000 295.440 ;
        RECT 4.400 288.640 1945.600 290.040 ;
        RECT 4.000 283.240 1946.000 288.640 ;
        RECT 4.400 281.840 1945.600 283.240 ;
        RECT 4.000 276.440 1946.000 281.840 ;
        RECT 4.400 275.040 1945.600 276.440 ;
        RECT 4.000 269.640 1946.000 275.040 ;
        RECT 4.400 268.240 1945.600 269.640 ;
        RECT 4.000 262.840 1946.000 268.240 ;
        RECT 4.400 261.440 1945.600 262.840 ;
        RECT 4.000 256.040 1946.000 261.440 ;
        RECT 4.400 254.640 1945.600 256.040 ;
        RECT 4.000 249.240 1946.000 254.640 ;
        RECT 4.400 247.840 1945.600 249.240 ;
        RECT 4.000 242.440 1946.000 247.840 ;
        RECT 4.400 241.040 1945.600 242.440 ;
        RECT 4.000 235.640 1946.000 241.040 ;
        RECT 4.400 234.240 1945.600 235.640 ;
        RECT 4.000 228.840 1946.000 234.240 ;
        RECT 4.400 227.440 1945.600 228.840 ;
        RECT 4.000 222.040 1946.000 227.440 ;
        RECT 4.400 220.640 1945.600 222.040 ;
        RECT 4.000 215.240 1946.000 220.640 ;
        RECT 4.400 213.840 1945.600 215.240 ;
        RECT 4.000 208.440 1946.000 213.840 ;
        RECT 4.400 207.040 1945.600 208.440 ;
        RECT 4.000 201.640 1946.000 207.040 ;
        RECT 4.400 200.240 1945.600 201.640 ;
        RECT 4.000 194.840 1946.000 200.240 ;
        RECT 4.400 193.440 1945.600 194.840 ;
        RECT 4.000 188.040 1946.000 193.440 ;
        RECT 4.400 186.640 1945.600 188.040 ;
        RECT 4.000 181.240 1946.000 186.640 ;
        RECT 4.400 179.840 1945.600 181.240 ;
        RECT 4.000 174.440 1946.000 179.840 ;
        RECT 4.400 173.040 1945.600 174.440 ;
        RECT 4.000 167.640 1946.000 173.040 ;
        RECT 4.400 166.240 1945.600 167.640 ;
        RECT 4.000 160.840 1946.000 166.240 ;
        RECT 4.400 159.440 1945.600 160.840 ;
        RECT 4.000 154.040 1946.000 159.440 ;
        RECT 4.400 152.640 1945.600 154.040 ;
        RECT 4.000 147.240 1946.000 152.640 ;
        RECT 4.400 145.840 1945.600 147.240 ;
        RECT 4.000 140.440 1946.000 145.840 ;
        RECT 4.400 139.040 1945.600 140.440 ;
        RECT 4.000 133.640 1946.000 139.040 ;
        RECT 4.400 132.240 1945.600 133.640 ;
        RECT 4.000 126.840 1946.000 132.240 ;
        RECT 4.400 125.440 1945.600 126.840 ;
        RECT 4.000 120.040 1946.000 125.440 ;
        RECT 4.400 118.640 1945.600 120.040 ;
        RECT 4.000 113.240 1946.000 118.640 ;
        RECT 4.400 111.840 1945.600 113.240 ;
        RECT 4.000 106.440 1946.000 111.840 ;
        RECT 4.400 105.040 1945.600 106.440 ;
        RECT 4.000 99.640 1946.000 105.040 ;
        RECT 4.400 98.240 1945.600 99.640 ;
        RECT 4.000 92.840 1946.000 98.240 ;
        RECT 4.400 91.440 1945.600 92.840 ;
        RECT 4.000 86.040 1946.000 91.440 ;
        RECT 4.400 84.640 1945.600 86.040 ;
        RECT 4.000 79.240 1946.000 84.640 ;
        RECT 4.400 77.840 1945.600 79.240 ;
        RECT 4.000 72.440 1946.000 77.840 ;
        RECT 4.400 71.040 1945.600 72.440 ;
        RECT 4.000 65.640 1946.000 71.040 ;
        RECT 4.400 64.240 1945.600 65.640 ;
        RECT 4.000 58.840 1946.000 64.240 ;
        RECT 4.400 57.440 1945.600 58.840 ;
        RECT 4.000 52.040 1946.000 57.440 ;
        RECT 4.400 50.640 1945.600 52.040 ;
        RECT 4.000 45.240 1946.000 50.640 ;
        RECT 4.400 43.840 1945.600 45.240 ;
        RECT 4.000 38.440 1946.000 43.840 ;
        RECT 4.400 37.040 1945.600 38.440 ;
        RECT 4.000 31.640 1946.000 37.040 ;
        RECT 4.400 30.240 1945.600 31.640 ;
        RECT 4.000 24.840 1946.000 30.240 ;
        RECT 4.400 23.440 1945.600 24.840 ;
        RECT 4.000 18.040 1946.000 23.440 ;
        RECT 4.400 16.640 1945.600 18.040 ;
        RECT 4.000 11.240 1946.000 16.640 ;
        RECT 4.400 10.375 1945.600 11.240 ;
      LAYER met4 ;
        RECT 61.015 11.735 97.440 1935.105 ;
        RECT 99.840 11.735 174.240 1935.105 ;
        RECT 176.640 11.735 251.040 1935.105 ;
        RECT 253.440 11.735 327.840 1935.105 ;
        RECT 330.240 11.735 404.640 1935.105 ;
        RECT 407.040 11.735 481.440 1935.105 ;
        RECT 483.840 11.735 558.240 1935.105 ;
        RECT 560.640 11.735 635.040 1935.105 ;
        RECT 637.440 11.735 711.840 1935.105 ;
        RECT 714.240 11.735 788.640 1935.105 ;
        RECT 791.040 11.735 865.440 1935.105 ;
        RECT 867.840 11.735 942.240 1935.105 ;
        RECT 944.640 11.735 1019.040 1935.105 ;
        RECT 1021.440 11.735 1095.840 1935.105 ;
        RECT 1098.240 11.735 1172.640 1935.105 ;
        RECT 1175.040 11.735 1249.440 1935.105 ;
        RECT 1251.840 11.735 1326.240 1935.105 ;
        RECT 1328.640 11.735 1403.040 1935.105 ;
        RECT 1405.440 11.735 1479.840 1935.105 ;
        RECT 1482.240 11.735 1556.640 1935.105 ;
        RECT 1559.040 11.735 1633.440 1935.105 ;
        RECT 1635.840 11.735 1710.240 1935.105 ;
        RECT 1712.640 11.735 1780.825 1935.105 ;
  END
END top
END LIBRARY

