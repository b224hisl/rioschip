magic
tech sky130B
magscale 1 2
timestamp 1662987570
<< viali >>
rect 28181 13821 28215 13855
rect 28181 10013 28215 10047
rect 27997 9877 28031 9911
rect 15117 7361 15151 7395
rect 15025 7157 15059 7191
rect 7481 2397 7515 2431
rect 7297 2261 7331 2295
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 4424 27770
rect 4476 27718 4488 27770
rect 4540 27718 4552 27770
rect 4604 27718 4616 27770
rect 4668 27718 4680 27770
rect 4732 27718 11372 27770
rect 11424 27718 11436 27770
rect 11488 27718 11500 27770
rect 11552 27718 11564 27770
rect 11616 27718 11628 27770
rect 11680 27718 18320 27770
rect 18372 27718 18384 27770
rect 18436 27718 18448 27770
rect 18500 27718 18512 27770
rect 18564 27718 18576 27770
rect 18628 27718 25268 27770
rect 25320 27718 25332 27770
rect 25384 27718 25396 27770
rect 25448 27718 25460 27770
rect 25512 27718 25524 27770
rect 25576 27718 28888 27770
rect 1104 27696 28888 27718
rect 1104 27226 28888 27248
rect 1104 27174 7898 27226
rect 7950 27174 7962 27226
rect 8014 27174 8026 27226
rect 8078 27174 8090 27226
rect 8142 27174 8154 27226
rect 8206 27174 14846 27226
rect 14898 27174 14910 27226
rect 14962 27174 14974 27226
rect 15026 27174 15038 27226
rect 15090 27174 15102 27226
rect 15154 27174 21794 27226
rect 21846 27174 21858 27226
rect 21910 27174 21922 27226
rect 21974 27174 21986 27226
rect 22038 27174 22050 27226
rect 22102 27174 28888 27226
rect 1104 27152 28888 27174
rect 1104 26682 28888 26704
rect 1104 26630 4424 26682
rect 4476 26630 4488 26682
rect 4540 26630 4552 26682
rect 4604 26630 4616 26682
rect 4668 26630 4680 26682
rect 4732 26630 11372 26682
rect 11424 26630 11436 26682
rect 11488 26630 11500 26682
rect 11552 26630 11564 26682
rect 11616 26630 11628 26682
rect 11680 26630 18320 26682
rect 18372 26630 18384 26682
rect 18436 26630 18448 26682
rect 18500 26630 18512 26682
rect 18564 26630 18576 26682
rect 18628 26630 25268 26682
rect 25320 26630 25332 26682
rect 25384 26630 25396 26682
rect 25448 26630 25460 26682
rect 25512 26630 25524 26682
rect 25576 26630 28888 26682
rect 1104 26608 28888 26630
rect 1104 26138 28888 26160
rect 1104 26086 7898 26138
rect 7950 26086 7962 26138
rect 8014 26086 8026 26138
rect 8078 26086 8090 26138
rect 8142 26086 8154 26138
rect 8206 26086 14846 26138
rect 14898 26086 14910 26138
rect 14962 26086 14974 26138
rect 15026 26086 15038 26138
rect 15090 26086 15102 26138
rect 15154 26086 21794 26138
rect 21846 26086 21858 26138
rect 21910 26086 21922 26138
rect 21974 26086 21986 26138
rect 22038 26086 22050 26138
rect 22102 26086 28888 26138
rect 1104 26064 28888 26086
rect 1104 25594 28888 25616
rect 1104 25542 4424 25594
rect 4476 25542 4488 25594
rect 4540 25542 4552 25594
rect 4604 25542 4616 25594
rect 4668 25542 4680 25594
rect 4732 25542 11372 25594
rect 11424 25542 11436 25594
rect 11488 25542 11500 25594
rect 11552 25542 11564 25594
rect 11616 25542 11628 25594
rect 11680 25542 18320 25594
rect 18372 25542 18384 25594
rect 18436 25542 18448 25594
rect 18500 25542 18512 25594
rect 18564 25542 18576 25594
rect 18628 25542 25268 25594
rect 25320 25542 25332 25594
rect 25384 25542 25396 25594
rect 25448 25542 25460 25594
rect 25512 25542 25524 25594
rect 25576 25542 28888 25594
rect 1104 25520 28888 25542
rect 1104 25050 28888 25072
rect 1104 24998 7898 25050
rect 7950 24998 7962 25050
rect 8014 24998 8026 25050
rect 8078 24998 8090 25050
rect 8142 24998 8154 25050
rect 8206 24998 14846 25050
rect 14898 24998 14910 25050
rect 14962 24998 14974 25050
rect 15026 24998 15038 25050
rect 15090 24998 15102 25050
rect 15154 24998 21794 25050
rect 21846 24998 21858 25050
rect 21910 24998 21922 25050
rect 21974 24998 21986 25050
rect 22038 24998 22050 25050
rect 22102 24998 28888 25050
rect 1104 24976 28888 24998
rect 1104 24506 28888 24528
rect 1104 24454 4424 24506
rect 4476 24454 4488 24506
rect 4540 24454 4552 24506
rect 4604 24454 4616 24506
rect 4668 24454 4680 24506
rect 4732 24454 11372 24506
rect 11424 24454 11436 24506
rect 11488 24454 11500 24506
rect 11552 24454 11564 24506
rect 11616 24454 11628 24506
rect 11680 24454 18320 24506
rect 18372 24454 18384 24506
rect 18436 24454 18448 24506
rect 18500 24454 18512 24506
rect 18564 24454 18576 24506
rect 18628 24454 25268 24506
rect 25320 24454 25332 24506
rect 25384 24454 25396 24506
rect 25448 24454 25460 24506
rect 25512 24454 25524 24506
rect 25576 24454 28888 24506
rect 1104 24432 28888 24454
rect 1104 23962 28888 23984
rect 1104 23910 7898 23962
rect 7950 23910 7962 23962
rect 8014 23910 8026 23962
rect 8078 23910 8090 23962
rect 8142 23910 8154 23962
rect 8206 23910 14846 23962
rect 14898 23910 14910 23962
rect 14962 23910 14974 23962
rect 15026 23910 15038 23962
rect 15090 23910 15102 23962
rect 15154 23910 21794 23962
rect 21846 23910 21858 23962
rect 21910 23910 21922 23962
rect 21974 23910 21986 23962
rect 22038 23910 22050 23962
rect 22102 23910 28888 23962
rect 1104 23888 28888 23910
rect 1104 23418 28888 23440
rect 1104 23366 4424 23418
rect 4476 23366 4488 23418
rect 4540 23366 4552 23418
rect 4604 23366 4616 23418
rect 4668 23366 4680 23418
rect 4732 23366 11372 23418
rect 11424 23366 11436 23418
rect 11488 23366 11500 23418
rect 11552 23366 11564 23418
rect 11616 23366 11628 23418
rect 11680 23366 18320 23418
rect 18372 23366 18384 23418
rect 18436 23366 18448 23418
rect 18500 23366 18512 23418
rect 18564 23366 18576 23418
rect 18628 23366 25268 23418
rect 25320 23366 25332 23418
rect 25384 23366 25396 23418
rect 25448 23366 25460 23418
rect 25512 23366 25524 23418
rect 25576 23366 28888 23418
rect 1104 23344 28888 23366
rect 1104 22874 28888 22896
rect 1104 22822 7898 22874
rect 7950 22822 7962 22874
rect 8014 22822 8026 22874
rect 8078 22822 8090 22874
rect 8142 22822 8154 22874
rect 8206 22822 14846 22874
rect 14898 22822 14910 22874
rect 14962 22822 14974 22874
rect 15026 22822 15038 22874
rect 15090 22822 15102 22874
rect 15154 22822 21794 22874
rect 21846 22822 21858 22874
rect 21910 22822 21922 22874
rect 21974 22822 21986 22874
rect 22038 22822 22050 22874
rect 22102 22822 28888 22874
rect 1104 22800 28888 22822
rect 1104 22330 28888 22352
rect 1104 22278 4424 22330
rect 4476 22278 4488 22330
rect 4540 22278 4552 22330
rect 4604 22278 4616 22330
rect 4668 22278 4680 22330
rect 4732 22278 11372 22330
rect 11424 22278 11436 22330
rect 11488 22278 11500 22330
rect 11552 22278 11564 22330
rect 11616 22278 11628 22330
rect 11680 22278 18320 22330
rect 18372 22278 18384 22330
rect 18436 22278 18448 22330
rect 18500 22278 18512 22330
rect 18564 22278 18576 22330
rect 18628 22278 25268 22330
rect 25320 22278 25332 22330
rect 25384 22278 25396 22330
rect 25448 22278 25460 22330
rect 25512 22278 25524 22330
rect 25576 22278 28888 22330
rect 1104 22256 28888 22278
rect 1104 21786 28888 21808
rect 1104 21734 7898 21786
rect 7950 21734 7962 21786
rect 8014 21734 8026 21786
rect 8078 21734 8090 21786
rect 8142 21734 8154 21786
rect 8206 21734 14846 21786
rect 14898 21734 14910 21786
rect 14962 21734 14974 21786
rect 15026 21734 15038 21786
rect 15090 21734 15102 21786
rect 15154 21734 21794 21786
rect 21846 21734 21858 21786
rect 21910 21734 21922 21786
rect 21974 21734 21986 21786
rect 22038 21734 22050 21786
rect 22102 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 4424 21242
rect 4476 21190 4488 21242
rect 4540 21190 4552 21242
rect 4604 21190 4616 21242
rect 4668 21190 4680 21242
rect 4732 21190 11372 21242
rect 11424 21190 11436 21242
rect 11488 21190 11500 21242
rect 11552 21190 11564 21242
rect 11616 21190 11628 21242
rect 11680 21190 18320 21242
rect 18372 21190 18384 21242
rect 18436 21190 18448 21242
rect 18500 21190 18512 21242
rect 18564 21190 18576 21242
rect 18628 21190 25268 21242
rect 25320 21190 25332 21242
rect 25384 21190 25396 21242
rect 25448 21190 25460 21242
rect 25512 21190 25524 21242
rect 25576 21190 28888 21242
rect 1104 21168 28888 21190
rect 1104 20698 28888 20720
rect 1104 20646 7898 20698
rect 7950 20646 7962 20698
rect 8014 20646 8026 20698
rect 8078 20646 8090 20698
rect 8142 20646 8154 20698
rect 8206 20646 14846 20698
rect 14898 20646 14910 20698
rect 14962 20646 14974 20698
rect 15026 20646 15038 20698
rect 15090 20646 15102 20698
rect 15154 20646 21794 20698
rect 21846 20646 21858 20698
rect 21910 20646 21922 20698
rect 21974 20646 21986 20698
rect 22038 20646 22050 20698
rect 22102 20646 28888 20698
rect 1104 20624 28888 20646
rect 1104 20154 28888 20176
rect 1104 20102 4424 20154
rect 4476 20102 4488 20154
rect 4540 20102 4552 20154
rect 4604 20102 4616 20154
rect 4668 20102 4680 20154
rect 4732 20102 11372 20154
rect 11424 20102 11436 20154
rect 11488 20102 11500 20154
rect 11552 20102 11564 20154
rect 11616 20102 11628 20154
rect 11680 20102 18320 20154
rect 18372 20102 18384 20154
rect 18436 20102 18448 20154
rect 18500 20102 18512 20154
rect 18564 20102 18576 20154
rect 18628 20102 25268 20154
rect 25320 20102 25332 20154
rect 25384 20102 25396 20154
rect 25448 20102 25460 20154
rect 25512 20102 25524 20154
rect 25576 20102 28888 20154
rect 1104 20080 28888 20102
rect 1104 19610 28888 19632
rect 1104 19558 7898 19610
rect 7950 19558 7962 19610
rect 8014 19558 8026 19610
rect 8078 19558 8090 19610
rect 8142 19558 8154 19610
rect 8206 19558 14846 19610
rect 14898 19558 14910 19610
rect 14962 19558 14974 19610
rect 15026 19558 15038 19610
rect 15090 19558 15102 19610
rect 15154 19558 21794 19610
rect 21846 19558 21858 19610
rect 21910 19558 21922 19610
rect 21974 19558 21986 19610
rect 22038 19558 22050 19610
rect 22102 19558 28888 19610
rect 1104 19536 28888 19558
rect 1104 19066 28888 19088
rect 1104 19014 4424 19066
rect 4476 19014 4488 19066
rect 4540 19014 4552 19066
rect 4604 19014 4616 19066
rect 4668 19014 4680 19066
rect 4732 19014 11372 19066
rect 11424 19014 11436 19066
rect 11488 19014 11500 19066
rect 11552 19014 11564 19066
rect 11616 19014 11628 19066
rect 11680 19014 18320 19066
rect 18372 19014 18384 19066
rect 18436 19014 18448 19066
rect 18500 19014 18512 19066
rect 18564 19014 18576 19066
rect 18628 19014 25268 19066
rect 25320 19014 25332 19066
rect 25384 19014 25396 19066
rect 25448 19014 25460 19066
rect 25512 19014 25524 19066
rect 25576 19014 28888 19066
rect 1104 18992 28888 19014
rect 1104 18522 28888 18544
rect 1104 18470 7898 18522
rect 7950 18470 7962 18522
rect 8014 18470 8026 18522
rect 8078 18470 8090 18522
rect 8142 18470 8154 18522
rect 8206 18470 14846 18522
rect 14898 18470 14910 18522
rect 14962 18470 14974 18522
rect 15026 18470 15038 18522
rect 15090 18470 15102 18522
rect 15154 18470 21794 18522
rect 21846 18470 21858 18522
rect 21910 18470 21922 18522
rect 21974 18470 21986 18522
rect 22038 18470 22050 18522
rect 22102 18470 28888 18522
rect 1104 18448 28888 18470
rect 1104 17978 28888 18000
rect 1104 17926 4424 17978
rect 4476 17926 4488 17978
rect 4540 17926 4552 17978
rect 4604 17926 4616 17978
rect 4668 17926 4680 17978
rect 4732 17926 11372 17978
rect 11424 17926 11436 17978
rect 11488 17926 11500 17978
rect 11552 17926 11564 17978
rect 11616 17926 11628 17978
rect 11680 17926 18320 17978
rect 18372 17926 18384 17978
rect 18436 17926 18448 17978
rect 18500 17926 18512 17978
rect 18564 17926 18576 17978
rect 18628 17926 25268 17978
rect 25320 17926 25332 17978
rect 25384 17926 25396 17978
rect 25448 17926 25460 17978
rect 25512 17926 25524 17978
rect 25576 17926 28888 17978
rect 1104 17904 28888 17926
rect 1104 17434 28888 17456
rect 1104 17382 7898 17434
rect 7950 17382 7962 17434
rect 8014 17382 8026 17434
rect 8078 17382 8090 17434
rect 8142 17382 8154 17434
rect 8206 17382 14846 17434
rect 14898 17382 14910 17434
rect 14962 17382 14974 17434
rect 15026 17382 15038 17434
rect 15090 17382 15102 17434
rect 15154 17382 21794 17434
rect 21846 17382 21858 17434
rect 21910 17382 21922 17434
rect 21974 17382 21986 17434
rect 22038 17382 22050 17434
rect 22102 17382 28888 17434
rect 1104 17360 28888 17382
rect 1104 16890 28888 16912
rect 1104 16838 4424 16890
rect 4476 16838 4488 16890
rect 4540 16838 4552 16890
rect 4604 16838 4616 16890
rect 4668 16838 4680 16890
rect 4732 16838 11372 16890
rect 11424 16838 11436 16890
rect 11488 16838 11500 16890
rect 11552 16838 11564 16890
rect 11616 16838 11628 16890
rect 11680 16838 18320 16890
rect 18372 16838 18384 16890
rect 18436 16838 18448 16890
rect 18500 16838 18512 16890
rect 18564 16838 18576 16890
rect 18628 16838 25268 16890
rect 25320 16838 25332 16890
rect 25384 16838 25396 16890
rect 25448 16838 25460 16890
rect 25512 16838 25524 16890
rect 25576 16838 28888 16890
rect 1104 16816 28888 16838
rect 1104 16346 28888 16368
rect 1104 16294 7898 16346
rect 7950 16294 7962 16346
rect 8014 16294 8026 16346
rect 8078 16294 8090 16346
rect 8142 16294 8154 16346
rect 8206 16294 14846 16346
rect 14898 16294 14910 16346
rect 14962 16294 14974 16346
rect 15026 16294 15038 16346
rect 15090 16294 15102 16346
rect 15154 16294 21794 16346
rect 21846 16294 21858 16346
rect 21910 16294 21922 16346
rect 21974 16294 21986 16346
rect 22038 16294 22050 16346
rect 22102 16294 28888 16346
rect 1104 16272 28888 16294
rect 1104 15802 28888 15824
rect 1104 15750 4424 15802
rect 4476 15750 4488 15802
rect 4540 15750 4552 15802
rect 4604 15750 4616 15802
rect 4668 15750 4680 15802
rect 4732 15750 11372 15802
rect 11424 15750 11436 15802
rect 11488 15750 11500 15802
rect 11552 15750 11564 15802
rect 11616 15750 11628 15802
rect 11680 15750 18320 15802
rect 18372 15750 18384 15802
rect 18436 15750 18448 15802
rect 18500 15750 18512 15802
rect 18564 15750 18576 15802
rect 18628 15750 25268 15802
rect 25320 15750 25332 15802
rect 25384 15750 25396 15802
rect 25448 15750 25460 15802
rect 25512 15750 25524 15802
rect 25576 15750 28888 15802
rect 1104 15728 28888 15750
rect 1104 15258 28888 15280
rect 1104 15206 7898 15258
rect 7950 15206 7962 15258
rect 8014 15206 8026 15258
rect 8078 15206 8090 15258
rect 8142 15206 8154 15258
rect 8206 15206 14846 15258
rect 14898 15206 14910 15258
rect 14962 15206 14974 15258
rect 15026 15206 15038 15258
rect 15090 15206 15102 15258
rect 15154 15206 21794 15258
rect 21846 15206 21858 15258
rect 21910 15206 21922 15258
rect 21974 15206 21986 15258
rect 22038 15206 22050 15258
rect 22102 15206 28888 15258
rect 1104 15184 28888 15206
rect 1104 14714 28888 14736
rect 1104 14662 4424 14714
rect 4476 14662 4488 14714
rect 4540 14662 4552 14714
rect 4604 14662 4616 14714
rect 4668 14662 4680 14714
rect 4732 14662 11372 14714
rect 11424 14662 11436 14714
rect 11488 14662 11500 14714
rect 11552 14662 11564 14714
rect 11616 14662 11628 14714
rect 11680 14662 18320 14714
rect 18372 14662 18384 14714
rect 18436 14662 18448 14714
rect 18500 14662 18512 14714
rect 18564 14662 18576 14714
rect 18628 14662 25268 14714
rect 25320 14662 25332 14714
rect 25384 14662 25396 14714
rect 25448 14662 25460 14714
rect 25512 14662 25524 14714
rect 25576 14662 28888 14714
rect 1104 14640 28888 14662
rect 1104 14170 28888 14192
rect 1104 14118 7898 14170
rect 7950 14118 7962 14170
rect 8014 14118 8026 14170
rect 8078 14118 8090 14170
rect 8142 14118 8154 14170
rect 8206 14118 14846 14170
rect 14898 14118 14910 14170
rect 14962 14118 14974 14170
rect 15026 14118 15038 14170
rect 15090 14118 15102 14170
rect 15154 14118 21794 14170
rect 21846 14118 21858 14170
rect 21910 14118 21922 14170
rect 21974 14118 21986 14170
rect 22038 14118 22050 14170
rect 22102 14118 28888 14170
rect 1104 14096 28888 14118
rect 28166 13852 28172 13864
rect 28127 13824 28172 13852
rect 28166 13812 28172 13824
rect 28224 13812 28230 13864
rect 1104 13626 28888 13648
rect 1104 13574 4424 13626
rect 4476 13574 4488 13626
rect 4540 13574 4552 13626
rect 4604 13574 4616 13626
rect 4668 13574 4680 13626
rect 4732 13574 11372 13626
rect 11424 13574 11436 13626
rect 11488 13574 11500 13626
rect 11552 13574 11564 13626
rect 11616 13574 11628 13626
rect 11680 13574 18320 13626
rect 18372 13574 18384 13626
rect 18436 13574 18448 13626
rect 18500 13574 18512 13626
rect 18564 13574 18576 13626
rect 18628 13574 25268 13626
rect 25320 13574 25332 13626
rect 25384 13574 25396 13626
rect 25448 13574 25460 13626
rect 25512 13574 25524 13626
rect 25576 13574 28888 13626
rect 1104 13552 28888 13574
rect 1104 13082 28888 13104
rect 1104 13030 7898 13082
rect 7950 13030 7962 13082
rect 8014 13030 8026 13082
rect 8078 13030 8090 13082
rect 8142 13030 8154 13082
rect 8206 13030 14846 13082
rect 14898 13030 14910 13082
rect 14962 13030 14974 13082
rect 15026 13030 15038 13082
rect 15090 13030 15102 13082
rect 15154 13030 21794 13082
rect 21846 13030 21858 13082
rect 21910 13030 21922 13082
rect 21974 13030 21986 13082
rect 22038 13030 22050 13082
rect 22102 13030 28888 13082
rect 1104 13008 28888 13030
rect 1104 12538 28888 12560
rect 1104 12486 4424 12538
rect 4476 12486 4488 12538
rect 4540 12486 4552 12538
rect 4604 12486 4616 12538
rect 4668 12486 4680 12538
rect 4732 12486 11372 12538
rect 11424 12486 11436 12538
rect 11488 12486 11500 12538
rect 11552 12486 11564 12538
rect 11616 12486 11628 12538
rect 11680 12486 18320 12538
rect 18372 12486 18384 12538
rect 18436 12486 18448 12538
rect 18500 12486 18512 12538
rect 18564 12486 18576 12538
rect 18628 12486 25268 12538
rect 25320 12486 25332 12538
rect 25384 12486 25396 12538
rect 25448 12486 25460 12538
rect 25512 12486 25524 12538
rect 25576 12486 28888 12538
rect 1104 12464 28888 12486
rect 1104 11994 28888 12016
rect 1104 11942 7898 11994
rect 7950 11942 7962 11994
rect 8014 11942 8026 11994
rect 8078 11942 8090 11994
rect 8142 11942 8154 11994
rect 8206 11942 14846 11994
rect 14898 11942 14910 11994
rect 14962 11942 14974 11994
rect 15026 11942 15038 11994
rect 15090 11942 15102 11994
rect 15154 11942 21794 11994
rect 21846 11942 21858 11994
rect 21910 11942 21922 11994
rect 21974 11942 21986 11994
rect 22038 11942 22050 11994
rect 22102 11942 28888 11994
rect 1104 11920 28888 11942
rect 1104 11450 28888 11472
rect 1104 11398 4424 11450
rect 4476 11398 4488 11450
rect 4540 11398 4552 11450
rect 4604 11398 4616 11450
rect 4668 11398 4680 11450
rect 4732 11398 11372 11450
rect 11424 11398 11436 11450
rect 11488 11398 11500 11450
rect 11552 11398 11564 11450
rect 11616 11398 11628 11450
rect 11680 11398 18320 11450
rect 18372 11398 18384 11450
rect 18436 11398 18448 11450
rect 18500 11398 18512 11450
rect 18564 11398 18576 11450
rect 18628 11398 25268 11450
rect 25320 11398 25332 11450
rect 25384 11398 25396 11450
rect 25448 11398 25460 11450
rect 25512 11398 25524 11450
rect 25576 11398 28888 11450
rect 1104 11376 28888 11398
rect 1104 10906 28888 10928
rect 1104 10854 7898 10906
rect 7950 10854 7962 10906
rect 8014 10854 8026 10906
rect 8078 10854 8090 10906
rect 8142 10854 8154 10906
rect 8206 10854 14846 10906
rect 14898 10854 14910 10906
rect 14962 10854 14974 10906
rect 15026 10854 15038 10906
rect 15090 10854 15102 10906
rect 15154 10854 21794 10906
rect 21846 10854 21858 10906
rect 21910 10854 21922 10906
rect 21974 10854 21986 10906
rect 22038 10854 22050 10906
rect 22102 10854 28888 10906
rect 1104 10832 28888 10854
rect 1104 10362 28888 10384
rect 1104 10310 4424 10362
rect 4476 10310 4488 10362
rect 4540 10310 4552 10362
rect 4604 10310 4616 10362
rect 4668 10310 4680 10362
rect 4732 10310 11372 10362
rect 11424 10310 11436 10362
rect 11488 10310 11500 10362
rect 11552 10310 11564 10362
rect 11616 10310 11628 10362
rect 11680 10310 18320 10362
rect 18372 10310 18384 10362
rect 18436 10310 18448 10362
rect 18500 10310 18512 10362
rect 18564 10310 18576 10362
rect 18628 10310 25268 10362
rect 25320 10310 25332 10362
rect 25384 10310 25396 10362
rect 25448 10310 25460 10362
rect 25512 10310 25524 10362
rect 25576 10310 28888 10362
rect 1104 10288 28888 10310
rect 27522 10004 27528 10056
rect 27580 10044 27586 10056
rect 28169 10047 28227 10053
rect 28169 10044 28181 10047
rect 27580 10016 28181 10044
rect 27580 10004 27586 10016
rect 28169 10013 28181 10016
rect 28215 10013 28227 10047
rect 28169 10007 28227 10013
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 27985 9911 28043 9917
rect 27985 9908 27997 9911
rect 14792 9880 27997 9908
rect 14792 9868 14798 9880
rect 27985 9877 27997 9880
rect 28031 9877 28043 9911
rect 27985 9871 28043 9877
rect 1104 9818 28888 9840
rect 1104 9766 7898 9818
rect 7950 9766 7962 9818
rect 8014 9766 8026 9818
rect 8078 9766 8090 9818
rect 8142 9766 8154 9818
rect 8206 9766 14846 9818
rect 14898 9766 14910 9818
rect 14962 9766 14974 9818
rect 15026 9766 15038 9818
rect 15090 9766 15102 9818
rect 15154 9766 21794 9818
rect 21846 9766 21858 9818
rect 21910 9766 21922 9818
rect 21974 9766 21986 9818
rect 22038 9766 22050 9818
rect 22102 9766 28888 9818
rect 1104 9744 28888 9766
rect 1104 9274 28888 9296
rect 1104 9222 4424 9274
rect 4476 9222 4488 9274
rect 4540 9222 4552 9274
rect 4604 9222 4616 9274
rect 4668 9222 4680 9274
rect 4732 9222 11372 9274
rect 11424 9222 11436 9274
rect 11488 9222 11500 9274
rect 11552 9222 11564 9274
rect 11616 9222 11628 9274
rect 11680 9222 18320 9274
rect 18372 9222 18384 9274
rect 18436 9222 18448 9274
rect 18500 9222 18512 9274
rect 18564 9222 18576 9274
rect 18628 9222 25268 9274
rect 25320 9222 25332 9274
rect 25384 9222 25396 9274
rect 25448 9222 25460 9274
rect 25512 9222 25524 9274
rect 25576 9222 28888 9274
rect 1104 9200 28888 9222
rect 1104 8730 28888 8752
rect 1104 8678 7898 8730
rect 7950 8678 7962 8730
rect 8014 8678 8026 8730
rect 8078 8678 8090 8730
rect 8142 8678 8154 8730
rect 8206 8678 14846 8730
rect 14898 8678 14910 8730
rect 14962 8678 14974 8730
rect 15026 8678 15038 8730
rect 15090 8678 15102 8730
rect 15154 8678 21794 8730
rect 21846 8678 21858 8730
rect 21910 8678 21922 8730
rect 21974 8678 21986 8730
rect 22038 8678 22050 8730
rect 22102 8678 28888 8730
rect 1104 8656 28888 8678
rect 1104 8186 28888 8208
rect 1104 8134 4424 8186
rect 4476 8134 4488 8186
rect 4540 8134 4552 8186
rect 4604 8134 4616 8186
rect 4668 8134 4680 8186
rect 4732 8134 11372 8186
rect 11424 8134 11436 8186
rect 11488 8134 11500 8186
rect 11552 8134 11564 8186
rect 11616 8134 11628 8186
rect 11680 8134 18320 8186
rect 18372 8134 18384 8186
rect 18436 8134 18448 8186
rect 18500 8134 18512 8186
rect 18564 8134 18576 8186
rect 18628 8134 25268 8186
rect 25320 8134 25332 8186
rect 25384 8134 25396 8186
rect 25448 8134 25460 8186
rect 25512 8134 25524 8186
rect 25576 8134 28888 8186
rect 1104 8112 28888 8134
rect 1104 7642 28888 7664
rect 1104 7590 7898 7642
rect 7950 7590 7962 7642
rect 8014 7590 8026 7642
rect 8078 7590 8090 7642
rect 8142 7590 8154 7642
rect 8206 7590 14846 7642
rect 14898 7590 14910 7642
rect 14962 7590 14974 7642
rect 15026 7590 15038 7642
rect 15090 7590 15102 7642
rect 15154 7590 21794 7642
rect 21846 7590 21858 7642
rect 21910 7590 21922 7642
rect 21974 7590 21986 7642
rect 22038 7590 22050 7642
rect 22102 7590 28888 7642
rect 1104 7568 28888 7590
rect 14734 7352 14740 7404
rect 14792 7392 14798 7404
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 14792 7364 15117 7392
rect 14792 7352 14798 7364
rect 15105 7361 15117 7364
rect 15151 7361 15163 7395
rect 15105 7355 15163 7361
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 15013 7191 15071 7197
rect 15013 7188 15025 7191
rect 7524 7160 15025 7188
rect 7524 7148 7530 7160
rect 15013 7157 15025 7160
rect 15059 7157 15071 7191
rect 15013 7151 15071 7157
rect 1104 7098 28888 7120
rect 1104 7046 4424 7098
rect 4476 7046 4488 7098
rect 4540 7046 4552 7098
rect 4604 7046 4616 7098
rect 4668 7046 4680 7098
rect 4732 7046 11372 7098
rect 11424 7046 11436 7098
rect 11488 7046 11500 7098
rect 11552 7046 11564 7098
rect 11616 7046 11628 7098
rect 11680 7046 18320 7098
rect 18372 7046 18384 7098
rect 18436 7046 18448 7098
rect 18500 7046 18512 7098
rect 18564 7046 18576 7098
rect 18628 7046 25268 7098
rect 25320 7046 25332 7098
rect 25384 7046 25396 7098
rect 25448 7046 25460 7098
rect 25512 7046 25524 7098
rect 25576 7046 28888 7098
rect 1104 7024 28888 7046
rect 1104 6554 28888 6576
rect 1104 6502 7898 6554
rect 7950 6502 7962 6554
rect 8014 6502 8026 6554
rect 8078 6502 8090 6554
rect 8142 6502 8154 6554
rect 8206 6502 14846 6554
rect 14898 6502 14910 6554
rect 14962 6502 14974 6554
rect 15026 6502 15038 6554
rect 15090 6502 15102 6554
rect 15154 6502 21794 6554
rect 21846 6502 21858 6554
rect 21910 6502 21922 6554
rect 21974 6502 21986 6554
rect 22038 6502 22050 6554
rect 22102 6502 28888 6554
rect 1104 6480 28888 6502
rect 1104 6010 28888 6032
rect 1104 5958 4424 6010
rect 4476 5958 4488 6010
rect 4540 5958 4552 6010
rect 4604 5958 4616 6010
rect 4668 5958 4680 6010
rect 4732 5958 11372 6010
rect 11424 5958 11436 6010
rect 11488 5958 11500 6010
rect 11552 5958 11564 6010
rect 11616 5958 11628 6010
rect 11680 5958 18320 6010
rect 18372 5958 18384 6010
rect 18436 5958 18448 6010
rect 18500 5958 18512 6010
rect 18564 5958 18576 6010
rect 18628 5958 25268 6010
rect 25320 5958 25332 6010
rect 25384 5958 25396 6010
rect 25448 5958 25460 6010
rect 25512 5958 25524 6010
rect 25576 5958 28888 6010
rect 1104 5936 28888 5958
rect 1104 5466 28888 5488
rect 1104 5414 7898 5466
rect 7950 5414 7962 5466
rect 8014 5414 8026 5466
rect 8078 5414 8090 5466
rect 8142 5414 8154 5466
rect 8206 5414 14846 5466
rect 14898 5414 14910 5466
rect 14962 5414 14974 5466
rect 15026 5414 15038 5466
rect 15090 5414 15102 5466
rect 15154 5414 21794 5466
rect 21846 5414 21858 5466
rect 21910 5414 21922 5466
rect 21974 5414 21986 5466
rect 22038 5414 22050 5466
rect 22102 5414 28888 5466
rect 1104 5392 28888 5414
rect 1104 4922 28888 4944
rect 1104 4870 4424 4922
rect 4476 4870 4488 4922
rect 4540 4870 4552 4922
rect 4604 4870 4616 4922
rect 4668 4870 4680 4922
rect 4732 4870 11372 4922
rect 11424 4870 11436 4922
rect 11488 4870 11500 4922
rect 11552 4870 11564 4922
rect 11616 4870 11628 4922
rect 11680 4870 18320 4922
rect 18372 4870 18384 4922
rect 18436 4870 18448 4922
rect 18500 4870 18512 4922
rect 18564 4870 18576 4922
rect 18628 4870 25268 4922
rect 25320 4870 25332 4922
rect 25384 4870 25396 4922
rect 25448 4870 25460 4922
rect 25512 4870 25524 4922
rect 25576 4870 28888 4922
rect 1104 4848 28888 4870
rect 1104 4378 28888 4400
rect 1104 4326 7898 4378
rect 7950 4326 7962 4378
rect 8014 4326 8026 4378
rect 8078 4326 8090 4378
rect 8142 4326 8154 4378
rect 8206 4326 14846 4378
rect 14898 4326 14910 4378
rect 14962 4326 14974 4378
rect 15026 4326 15038 4378
rect 15090 4326 15102 4378
rect 15154 4326 21794 4378
rect 21846 4326 21858 4378
rect 21910 4326 21922 4378
rect 21974 4326 21986 4378
rect 22038 4326 22050 4378
rect 22102 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 4424 3834
rect 4476 3782 4488 3834
rect 4540 3782 4552 3834
rect 4604 3782 4616 3834
rect 4668 3782 4680 3834
rect 4732 3782 11372 3834
rect 11424 3782 11436 3834
rect 11488 3782 11500 3834
rect 11552 3782 11564 3834
rect 11616 3782 11628 3834
rect 11680 3782 18320 3834
rect 18372 3782 18384 3834
rect 18436 3782 18448 3834
rect 18500 3782 18512 3834
rect 18564 3782 18576 3834
rect 18628 3782 25268 3834
rect 25320 3782 25332 3834
rect 25384 3782 25396 3834
rect 25448 3782 25460 3834
rect 25512 3782 25524 3834
rect 25576 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 7898 3290
rect 7950 3238 7962 3290
rect 8014 3238 8026 3290
rect 8078 3238 8090 3290
rect 8142 3238 8154 3290
rect 8206 3238 14846 3290
rect 14898 3238 14910 3290
rect 14962 3238 14974 3290
rect 15026 3238 15038 3290
rect 15090 3238 15102 3290
rect 15154 3238 21794 3290
rect 21846 3238 21858 3290
rect 21910 3238 21922 3290
rect 21974 3238 21986 3290
rect 22038 3238 22050 3290
rect 22102 3238 28888 3290
rect 1104 3216 28888 3238
rect 1104 2746 28888 2768
rect 1104 2694 4424 2746
rect 4476 2694 4488 2746
rect 4540 2694 4552 2746
rect 4604 2694 4616 2746
rect 4668 2694 4680 2746
rect 4732 2694 11372 2746
rect 11424 2694 11436 2746
rect 11488 2694 11500 2746
rect 11552 2694 11564 2746
rect 11616 2694 11628 2746
rect 11680 2694 18320 2746
rect 18372 2694 18384 2746
rect 18436 2694 18448 2746
rect 18500 2694 18512 2746
rect 18564 2694 18576 2746
rect 18628 2694 25268 2746
rect 25320 2694 25332 2746
rect 25384 2694 25396 2746
rect 25448 2694 25460 2746
rect 25512 2694 25524 2746
rect 25576 2694 28888 2746
rect 1104 2672 28888 2694
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 7156 2264 7297 2292
rect 7156 2252 7162 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 1104 2202 28888 2224
rect 1104 2150 7898 2202
rect 7950 2150 7962 2202
rect 8014 2150 8026 2202
rect 8078 2150 8090 2202
rect 8142 2150 8154 2202
rect 8206 2150 14846 2202
rect 14898 2150 14910 2202
rect 14962 2150 14974 2202
rect 15026 2150 15038 2202
rect 15090 2150 15102 2202
rect 15154 2150 21794 2202
rect 21846 2150 21858 2202
rect 21910 2150 21922 2202
rect 21974 2150 21986 2202
rect 22038 2150 22050 2202
rect 22102 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 4424 27718 4476 27770
rect 4488 27718 4540 27770
rect 4552 27718 4604 27770
rect 4616 27718 4668 27770
rect 4680 27718 4732 27770
rect 11372 27718 11424 27770
rect 11436 27718 11488 27770
rect 11500 27718 11552 27770
rect 11564 27718 11616 27770
rect 11628 27718 11680 27770
rect 18320 27718 18372 27770
rect 18384 27718 18436 27770
rect 18448 27718 18500 27770
rect 18512 27718 18564 27770
rect 18576 27718 18628 27770
rect 25268 27718 25320 27770
rect 25332 27718 25384 27770
rect 25396 27718 25448 27770
rect 25460 27718 25512 27770
rect 25524 27718 25576 27770
rect 7898 27174 7950 27226
rect 7962 27174 8014 27226
rect 8026 27174 8078 27226
rect 8090 27174 8142 27226
rect 8154 27174 8206 27226
rect 14846 27174 14898 27226
rect 14910 27174 14962 27226
rect 14974 27174 15026 27226
rect 15038 27174 15090 27226
rect 15102 27174 15154 27226
rect 21794 27174 21846 27226
rect 21858 27174 21910 27226
rect 21922 27174 21974 27226
rect 21986 27174 22038 27226
rect 22050 27174 22102 27226
rect 4424 26630 4476 26682
rect 4488 26630 4540 26682
rect 4552 26630 4604 26682
rect 4616 26630 4668 26682
rect 4680 26630 4732 26682
rect 11372 26630 11424 26682
rect 11436 26630 11488 26682
rect 11500 26630 11552 26682
rect 11564 26630 11616 26682
rect 11628 26630 11680 26682
rect 18320 26630 18372 26682
rect 18384 26630 18436 26682
rect 18448 26630 18500 26682
rect 18512 26630 18564 26682
rect 18576 26630 18628 26682
rect 25268 26630 25320 26682
rect 25332 26630 25384 26682
rect 25396 26630 25448 26682
rect 25460 26630 25512 26682
rect 25524 26630 25576 26682
rect 7898 26086 7950 26138
rect 7962 26086 8014 26138
rect 8026 26086 8078 26138
rect 8090 26086 8142 26138
rect 8154 26086 8206 26138
rect 14846 26086 14898 26138
rect 14910 26086 14962 26138
rect 14974 26086 15026 26138
rect 15038 26086 15090 26138
rect 15102 26086 15154 26138
rect 21794 26086 21846 26138
rect 21858 26086 21910 26138
rect 21922 26086 21974 26138
rect 21986 26086 22038 26138
rect 22050 26086 22102 26138
rect 4424 25542 4476 25594
rect 4488 25542 4540 25594
rect 4552 25542 4604 25594
rect 4616 25542 4668 25594
rect 4680 25542 4732 25594
rect 11372 25542 11424 25594
rect 11436 25542 11488 25594
rect 11500 25542 11552 25594
rect 11564 25542 11616 25594
rect 11628 25542 11680 25594
rect 18320 25542 18372 25594
rect 18384 25542 18436 25594
rect 18448 25542 18500 25594
rect 18512 25542 18564 25594
rect 18576 25542 18628 25594
rect 25268 25542 25320 25594
rect 25332 25542 25384 25594
rect 25396 25542 25448 25594
rect 25460 25542 25512 25594
rect 25524 25542 25576 25594
rect 7898 24998 7950 25050
rect 7962 24998 8014 25050
rect 8026 24998 8078 25050
rect 8090 24998 8142 25050
rect 8154 24998 8206 25050
rect 14846 24998 14898 25050
rect 14910 24998 14962 25050
rect 14974 24998 15026 25050
rect 15038 24998 15090 25050
rect 15102 24998 15154 25050
rect 21794 24998 21846 25050
rect 21858 24998 21910 25050
rect 21922 24998 21974 25050
rect 21986 24998 22038 25050
rect 22050 24998 22102 25050
rect 4424 24454 4476 24506
rect 4488 24454 4540 24506
rect 4552 24454 4604 24506
rect 4616 24454 4668 24506
rect 4680 24454 4732 24506
rect 11372 24454 11424 24506
rect 11436 24454 11488 24506
rect 11500 24454 11552 24506
rect 11564 24454 11616 24506
rect 11628 24454 11680 24506
rect 18320 24454 18372 24506
rect 18384 24454 18436 24506
rect 18448 24454 18500 24506
rect 18512 24454 18564 24506
rect 18576 24454 18628 24506
rect 25268 24454 25320 24506
rect 25332 24454 25384 24506
rect 25396 24454 25448 24506
rect 25460 24454 25512 24506
rect 25524 24454 25576 24506
rect 7898 23910 7950 23962
rect 7962 23910 8014 23962
rect 8026 23910 8078 23962
rect 8090 23910 8142 23962
rect 8154 23910 8206 23962
rect 14846 23910 14898 23962
rect 14910 23910 14962 23962
rect 14974 23910 15026 23962
rect 15038 23910 15090 23962
rect 15102 23910 15154 23962
rect 21794 23910 21846 23962
rect 21858 23910 21910 23962
rect 21922 23910 21974 23962
rect 21986 23910 22038 23962
rect 22050 23910 22102 23962
rect 4424 23366 4476 23418
rect 4488 23366 4540 23418
rect 4552 23366 4604 23418
rect 4616 23366 4668 23418
rect 4680 23366 4732 23418
rect 11372 23366 11424 23418
rect 11436 23366 11488 23418
rect 11500 23366 11552 23418
rect 11564 23366 11616 23418
rect 11628 23366 11680 23418
rect 18320 23366 18372 23418
rect 18384 23366 18436 23418
rect 18448 23366 18500 23418
rect 18512 23366 18564 23418
rect 18576 23366 18628 23418
rect 25268 23366 25320 23418
rect 25332 23366 25384 23418
rect 25396 23366 25448 23418
rect 25460 23366 25512 23418
rect 25524 23366 25576 23418
rect 7898 22822 7950 22874
rect 7962 22822 8014 22874
rect 8026 22822 8078 22874
rect 8090 22822 8142 22874
rect 8154 22822 8206 22874
rect 14846 22822 14898 22874
rect 14910 22822 14962 22874
rect 14974 22822 15026 22874
rect 15038 22822 15090 22874
rect 15102 22822 15154 22874
rect 21794 22822 21846 22874
rect 21858 22822 21910 22874
rect 21922 22822 21974 22874
rect 21986 22822 22038 22874
rect 22050 22822 22102 22874
rect 4424 22278 4476 22330
rect 4488 22278 4540 22330
rect 4552 22278 4604 22330
rect 4616 22278 4668 22330
rect 4680 22278 4732 22330
rect 11372 22278 11424 22330
rect 11436 22278 11488 22330
rect 11500 22278 11552 22330
rect 11564 22278 11616 22330
rect 11628 22278 11680 22330
rect 18320 22278 18372 22330
rect 18384 22278 18436 22330
rect 18448 22278 18500 22330
rect 18512 22278 18564 22330
rect 18576 22278 18628 22330
rect 25268 22278 25320 22330
rect 25332 22278 25384 22330
rect 25396 22278 25448 22330
rect 25460 22278 25512 22330
rect 25524 22278 25576 22330
rect 7898 21734 7950 21786
rect 7962 21734 8014 21786
rect 8026 21734 8078 21786
rect 8090 21734 8142 21786
rect 8154 21734 8206 21786
rect 14846 21734 14898 21786
rect 14910 21734 14962 21786
rect 14974 21734 15026 21786
rect 15038 21734 15090 21786
rect 15102 21734 15154 21786
rect 21794 21734 21846 21786
rect 21858 21734 21910 21786
rect 21922 21734 21974 21786
rect 21986 21734 22038 21786
rect 22050 21734 22102 21786
rect 4424 21190 4476 21242
rect 4488 21190 4540 21242
rect 4552 21190 4604 21242
rect 4616 21190 4668 21242
rect 4680 21190 4732 21242
rect 11372 21190 11424 21242
rect 11436 21190 11488 21242
rect 11500 21190 11552 21242
rect 11564 21190 11616 21242
rect 11628 21190 11680 21242
rect 18320 21190 18372 21242
rect 18384 21190 18436 21242
rect 18448 21190 18500 21242
rect 18512 21190 18564 21242
rect 18576 21190 18628 21242
rect 25268 21190 25320 21242
rect 25332 21190 25384 21242
rect 25396 21190 25448 21242
rect 25460 21190 25512 21242
rect 25524 21190 25576 21242
rect 7898 20646 7950 20698
rect 7962 20646 8014 20698
rect 8026 20646 8078 20698
rect 8090 20646 8142 20698
rect 8154 20646 8206 20698
rect 14846 20646 14898 20698
rect 14910 20646 14962 20698
rect 14974 20646 15026 20698
rect 15038 20646 15090 20698
rect 15102 20646 15154 20698
rect 21794 20646 21846 20698
rect 21858 20646 21910 20698
rect 21922 20646 21974 20698
rect 21986 20646 22038 20698
rect 22050 20646 22102 20698
rect 4424 20102 4476 20154
rect 4488 20102 4540 20154
rect 4552 20102 4604 20154
rect 4616 20102 4668 20154
rect 4680 20102 4732 20154
rect 11372 20102 11424 20154
rect 11436 20102 11488 20154
rect 11500 20102 11552 20154
rect 11564 20102 11616 20154
rect 11628 20102 11680 20154
rect 18320 20102 18372 20154
rect 18384 20102 18436 20154
rect 18448 20102 18500 20154
rect 18512 20102 18564 20154
rect 18576 20102 18628 20154
rect 25268 20102 25320 20154
rect 25332 20102 25384 20154
rect 25396 20102 25448 20154
rect 25460 20102 25512 20154
rect 25524 20102 25576 20154
rect 7898 19558 7950 19610
rect 7962 19558 8014 19610
rect 8026 19558 8078 19610
rect 8090 19558 8142 19610
rect 8154 19558 8206 19610
rect 14846 19558 14898 19610
rect 14910 19558 14962 19610
rect 14974 19558 15026 19610
rect 15038 19558 15090 19610
rect 15102 19558 15154 19610
rect 21794 19558 21846 19610
rect 21858 19558 21910 19610
rect 21922 19558 21974 19610
rect 21986 19558 22038 19610
rect 22050 19558 22102 19610
rect 4424 19014 4476 19066
rect 4488 19014 4540 19066
rect 4552 19014 4604 19066
rect 4616 19014 4668 19066
rect 4680 19014 4732 19066
rect 11372 19014 11424 19066
rect 11436 19014 11488 19066
rect 11500 19014 11552 19066
rect 11564 19014 11616 19066
rect 11628 19014 11680 19066
rect 18320 19014 18372 19066
rect 18384 19014 18436 19066
rect 18448 19014 18500 19066
rect 18512 19014 18564 19066
rect 18576 19014 18628 19066
rect 25268 19014 25320 19066
rect 25332 19014 25384 19066
rect 25396 19014 25448 19066
rect 25460 19014 25512 19066
rect 25524 19014 25576 19066
rect 7898 18470 7950 18522
rect 7962 18470 8014 18522
rect 8026 18470 8078 18522
rect 8090 18470 8142 18522
rect 8154 18470 8206 18522
rect 14846 18470 14898 18522
rect 14910 18470 14962 18522
rect 14974 18470 15026 18522
rect 15038 18470 15090 18522
rect 15102 18470 15154 18522
rect 21794 18470 21846 18522
rect 21858 18470 21910 18522
rect 21922 18470 21974 18522
rect 21986 18470 22038 18522
rect 22050 18470 22102 18522
rect 4424 17926 4476 17978
rect 4488 17926 4540 17978
rect 4552 17926 4604 17978
rect 4616 17926 4668 17978
rect 4680 17926 4732 17978
rect 11372 17926 11424 17978
rect 11436 17926 11488 17978
rect 11500 17926 11552 17978
rect 11564 17926 11616 17978
rect 11628 17926 11680 17978
rect 18320 17926 18372 17978
rect 18384 17926 18436 17978
rect 18448 17926 18500 17978
rect 18512 17926 18564 17978
rect 18576 17926 18628 17978
rect 25268 17926 25320 17978
rect 25332 17926 25384 17978
rect 25396 17926 25448 17978
rect 25460 17926 25512 17978
rect 25524 17926 25576 17978
rect 7898 17382 7950 17434
rect 7962 17382 8014 17434
rect 8026 17382 8078 17434
rect 8090 17382 8142 17434
rect 8154 17382 8206 17434
rect 14846 17382 14898 17434
rect 14910 17382 14962 17434
rect 14974 17382 15026 17434
rect 15038 17382 15090 17434
rect 15102 17382 15154 17434
rect 21794 17382 21846 17434
rect 21858 17382 21910 17434
rect 21922 17382 21974 17434
rect 21986 17382 22038 17434
rect 22050 17382 22102 17434
rect 4424 16838 4476 16890
rect 4488 16838 4540 16890
rect 4552 16838 4604 16890
rect 4616 16838 4668 16890
rect 4680 16838 4732 16890
rect 11372 16838 11424 16890
rect 11436 16838 11488 16890
rect 11500 16838 11552 16890
rect 11564 16838 11616 16890
rect 11628 16838 11680 16890
rect 18320 16838 18372 16890
rect 18384 16838 18436 16890
rect 18448 16838 18500 16890
rect 18512 16838 18564 16890
rect 18576 16838 18628 16890
rect 25268 16838 25320 16890
rect 25332 16838 25384 16890
rect 25396 16838 25448 16890
rect 25460 16838 25512 16890
rect 25524 16838 25576 16890
rect 7898 16294 7950 16346
rect 7962 16294 8014 16346
rect 8026 16294 8078 16346
rect 8090 16294 8142 16346
rect 8154 16294 8206 16346
rect 14846 16294 14898 16346
rect 14910 16294 14962 16346
rect 14974 16294 15026 16346
rect 15038 16294 15090 16346
rect 15102 16294 15154 16346
rect 21794 16294 21846 16346
rect 21858 16294 21910 16346
rect 21922 16294 21974 16346
rect 21986 16294 22038 16346
rect 22050 16294 22102 16346
rect 4424 15750 4476 15802
rect 4488 15750 4540 15802
rect 4552 15750 4604 15802
rect 4616 15750 4668 15802
rect 4680 15750 4732 15802
rect 11372 15750 11424 15802
rect 11436 15750 11488 15802
rect 11500 15750 11552 15802
rect 11564 15750 11616 15802
rect 11628 15750 11680 15802
rect 18320 15750 18372 15802
rect 18384 15750 18436 15802
rect 18448 15750 18500 15802
rect 18512 15750 18564 15802
rect 18576 15750 18628 15802
rect 25268 15750 25320 15802
rect 25332 15750 25384 15802
rect 25396 15750 25448 15802
rect 25460 15750 25512 15802
rect 25524 15750 25576 15802
rect 7898 15206 7950 15258
rect 7962 15206 8014 15258
rect 8026 15206 8078 15258
rect 8090 15206 8142 15258
rect 8154 15206 8206 15258
rect 14846 15206 14898 15258
rect 14910 15206 14962 15258
rect 14974 15206 15026 15258
rect 15038 15206 15090 15258
rect 15102 15206 15154 15258
rect 21794 15206 21846 15258
rect 21858 15206 21910 15258
rect 21922 15206 21974 15258
rect 21986 15206 22038 15258
rect 22050 15206 22102 15258
rect 4424 14662 4476 14714
rect 4488 14662 4540 14714
rect 4552 14662 4604 14714
rect 4616 14662 4668 14714
rect 4680 14662 4732 14714
rect 11372 14662 11424 14714
rect 11436 14662 11488 14714
rect 11500 14662 11552 14714
rect 11564 14662 11616 14714
rect 11628 14662 11680 14714
rect 18320 14662 18372 14714
rect 18384 14662 18436 14714
rect 18448 14662 18500 14714
rect 18512 14662 18564 14714
rect 18576 14662 18628 14714
rect 25268 14662 25320 14714
rect 25332 14662 25384 14714
rect 25396 14662 25448 14714
rect 25460 14662 25512 14714
rect 25524 14662 25576 14714
rect 7898 14118 7950 14170
rect 7962 14118 8014 14170
rect 8026 14118 8078 14170
rect 8090 14118 8142 14170
rect 8154 14118 8206 14170
rect 14846 14118 14898 14170
rect 14910 14118 14962 14170
rect 14974 14118 15026 14170
rect 15038 14118 15090 14170
rect 15102 14118 15154 14170
rect 21794 14118 21846 14170
rect 21858 14118 21910 14170
rect 21922 14118 21974 14170
rect 21986 14118 22038 14170
rect 22050 14118 22102 14170
rect 28172 13855 28224 13864
rect 28172 13821 28181 13855
rect 28181 13821 28215 13855
rect 28215 13821 28224 13855
rect 28172 13812 28224 13821
rect 4424 13574 4476 13626
rect 4488 13574 4540 13626
rect 4552 13574 4604 13626
rect 4616 13574 4668 13626
rect 4680 13574 4732 13626
rect 11372 13574 11424 13626
rect 11436 13574 11488 13626
rect 11500 13574 11552 13626
rect 11564 13574 11616 13626
rect 11628 13574 11680 13626
rect 18320 13574 18372 13626
rect 18384 13574 18436 13626
rect 18448 13574 18500 13626
rect 18512 13574 18564 13626
rect 18576 13574 18628 13626
rect 25268 13574 25320 13626
rect 25332 13574 25384 13626
rect 25396 13574 25448 13626
rect 25460 13574 25512 13626
rect 25524 13574 25576 13626
rect 7898 13030 7950 13082
rect 7962 13030 8014 13082
rect 8026 13030 8078 13082
rect 8090 13030 8142 13082
rect 8154 13030 8206 13082
rect 14846 13030 14898 13082
rect 14910 13030 14962 13082
rect 14974 13030 15026 13082
rect 15038 13030 15090 13082
rect 15102 13030 15154 13082
rect 21794 13030 21846 13082
rect 21858 13030 21910 13082
rect 21922 13030 21974 13082
rect 21986 13030 22038 13082
rect 22050 13030 22102 13082
rect 4424 12486 4476 12538
rect 4488 12486 4540 12538
rect 4552 12486 4604 12538
rect 4616 12486 4668 12538
rect 4680 12486 4732 12538
rect 11372 12486 11424 12538
rect 11436 12486 11488 12538
rect 11500 12486 11552 12538
rect 11564 12486 11616 12538
rect 11628 12486 11680 12538
rect 18320 12486 18372 12538
rect 18384 12486 18436 12538
rect 18448 12486 18500 12538
rect 18512 12486 18564 12538
rect 18576 12486 18628 12538
rect 25268 12486 25320 12538
rect 25332 12486 25384 12538
rect 25396 12486 25448 12538
rect 25460 12486 25512 12538
rect 25524 12486 25576 12538
rect 7898 11942 7950 11994
rect 7962 11942 8014 11994
rect 8026 11942 8078 11994
rect 8090 11942 8142 11994
rect 8154 11942 8206 11994
rect 14846 11942 14898 11994
rect 14910 11942 14962 11994
rect 14974 11942 15026 11994
rect 15038 11942 15090 11994
rect 15102 11942 15154 11994
rect 21794 11942 21846 11994
rect 21858 11942 21910 11994
rect 21922 11942 21974 11994
rect 21986 11942 22038 11994
rect 22050 11942 22102 11994
rect 4424 11398 4476 11450
rect 4488 11398 4540 11450
rect 4552 11398 4604 11450
rect 4616 11398 4668 11450
rect 4680 11398 4732 11450
rect 11372 11398 11424 11450
rect 11436 11398 11488 11450
rect 11500 11398 11552 11450
rect 11564 11398 11616 11450
rect 11628 11398 11680 11450
rect 18320 11398 18372 11450
rect 18384 11398 18436 11450
rect 18448 11398 18500 11450
rect 18512 11398 18564 11450
rect 18576 11398 18628 11450
rect 25268 11398 25320 11450
rect 25332 11398 25384 11450
rect 25396 11398 25448 11450
rect 25460 11398 25512 11450
rect 25524 11398 25576 11450
rect 7898 10854 7950 10906
rect 7962 10854 8014 10906
rect 8026 10854 8078 10906
rect 8090 10854 8142 10906
rect 8154 10854 8206 10906
rect 14846 10854 14898 10906
rect 14910 10854 14962 10906
rect 14974 10854 15026 10906
rect 15038 10854 15090 10906
rect 15102 10854 15154 10906
rect 21794 10854 21846 10906
rect 21858 10854 21910 10906
rect 21922 10854 21974 10906
rect 21986 10854 22038 10906
rect 22050 10854 22102 10906
rect 4424 10310 4476 10362
rect 4488 10310 4540 10362
rect 4552 10310 4604 10362
rect 4616 10310 4668 10362
rect 4680 10310 4732 10362
rect 11372 10310 11424 10362
rect 11436 10310 11488 10362
rect 11500 10310 11552 10362
rect 11564 10310 11616 10362
rect 11628 10310 11680 10362
rect 18320 10310 18372 10362
rect 18384 10310 18436 10362
rect 18448 10310 18500 10362
rect 18512 10310 18564 10362
rect 18576 10310 18628 10362
rect 25268 10310 25320 10362
rect 25332 10310 25384 10362
rect 25396 10310 25448 10362
rect 25460 10310 25512 10362
rect 25524 10310 25576 10362
rect 27528 10004 27580 10056
rect 14740 9868 14792 9920
rect 7898 9766 7950 9818
rect 7962 9766 8014 9818
rect 8026 9766 8078 9818
rect 8090 9766 8142 9818
rect 8154 9766 8206 9818
rect 14846 9766 14898 9818
rect 14910 9766 14962 9818
rect 14974 9766 15026 9818
rect 15038 9766 15090 9818
rect 15102 9766 15154 9818
rect 21794 9766 21846 9818
rect 21858 9766 21910 9818
rect 21922 9766 21974 9818
rect 21986 9766 22038 9818
rect 22050 9766 22102 9818
rect 4424 9222 4476 9274
rect 4488 9222 4540 9274
rect 4552 9222 4604 9274
rect 4616 9222 4668 9274
rect 4680 9222 4732 9274
rect 11372 9222 11424 9274
rect 11436 9222 11488 9274
rect 11500 9222 11552 9274
rect 11564 9222 11616 9274
rect 11628 9222 11680 9274
rect 18320 9222 18372 9274
rect 18384 9222 18436 9274
rect 18448 9222 18500 9274
rect 18512 9222 18564 9274
rect 18576 9222 18628 9274
rect 25268 9222 25320 9274
rect 25332 9222 25384 9274
rect 25396 9222 25448 9274
rect 25460 9222 25512 9274
rect 25524 9222 25576 9274
rect 7898 8678 7950 8730
rect 7962 8678 8014 8730
rect 8026 8678 8078 8730
rect 8090 8678 8142 8730
rect 8154 8678 8206 8730
rect 14846 8678 14898 8730
rect 14910 8678 14962 8730
rect 14974 8678 15026 8730
rect 15038 8678 15090 8730
rect 15102 8678 15154 8730
rect 21794 8678 21846 8730
rect 21858 8678 21910 8730
rect 21922 8678 21974 8730
rect 21986 8678 22038 8730
rect 22050 8678 22102 8730
rect 4424 8134 4476 8186
rect 4488 8134 4540 8186
rect 4552 8134 4604 8186
rect 4616 8134 4668 8186
rect 4680 8134 4732 8186
rect 11372 8134 11424 8186
rect 11436 8134 11488 8186
rect 11500 8134 11552 8186
rect 11564 8134 11616 8186
rect 11628 8134 11680 8186
rect 18320 8134 18372 8186
rect 18384 8134 18436 8186
rect 18448 8134 18500 8186
rect 18512 8134 18564 8186
rect 18576 8134 18628 8186
rect 25268 8134 25320 8186
rect 25332 8134 25384 8186
rect 25396 8134 25448 8186
rect 25460 8134 25512 8186
rect 25524 8134 25576 8186
rect 7898 7590 7950 7642
rect 7962 7590 8014 7642
rect 8026 7590 8078 7642
rect 8090 7590 8142 7642
rect 8154 7590 8206 7642
rect 14846 7590 14898 7642
rect 14910 7590 14962 7642
rect 14974 7590 15026 7642
rect 15038 7590 15090 7642
rect 15102 7590 15154 7642
rect 21794 7590 21846 7642
rect 21858 7590 21910 7642
rect 21922 7590 21974 7642
rect 21986 7590 22038 7642
rect 22050 7590 22102 7642
rect 14740 7352 14792 7404
rect 7472 7148 7524 7200
rect 4424 7046 4476 7098
rect 4488 7046 4540 7098
rect 4552 7046 4604 7098
rect 4616 7046 4668 7098
rect 4680 7046 4732 7098
rect 11372 7046 11424 7098
rect 11436 7046 11488 7098
rect 11500 7046 11552 7098
rect 11564 7046 11616 7098
rect 11628 7046 11680 7098
rect 18320 7046 18372 7098
rect 18384 7046 18436 7098
rect 18448 7046 18500 7098
rect 18512 7046 18564 7098
rect 18576 7046 18628 7098
rect 25268 7046 25320 7098
rect 25332 7046 25384 7098
rect 25396 7046 25448 7098
rect 25460 7046 25512 7098
rect 25524 7046 25576 7098
rect 7898 6502 7950 6554
rect 7962 6502 8014 6554
rect 8026 6502 8078 6554
rect 8090 6502 8142 6554
rect 8154 6502 8206 6554
rect 14846 6502 14898 6554
rect 14910 6502 14962 6554
rect 14974 6502 15026 6554
rect 15038 6502 15090 6554
rect 15102 6502 15154 6554
rect 21794 6502 21846 6554
rect 21858 6502 21910 6554
rect 21922 6502 21974 6554
rect 21986 6502 22038 6554
rect 22050 6502 22102 6554
rect 4424 5958 4476 6010
rect 4488 5958 4540 6010
rect 4552 5958 4604 6010
rect 4616 5958 4668 6010
rect 4680 5958 4732 6010
rect 11372 5958 11424 6010
rect 11436 5958 11488 6010
rect 11500 5958 11552 6010
rect 11564 5958 11616 6010
rect 11628 5958 11680 6010
rect 18320 5958 18372 6010
rect 18384 5958 18436 6010
rect 18448 5958 18500 6010
rect 18512 5958 18564 6010
rect 18576 5958 18628 6010
rect 25268 5958 25320 6010
rect 25332 5958 25384 6010
rect 25396 5958 25448 6010
rect 25460 5958 25512 6010
rect 25524 5958 25576 6010
rect 7898 5414 7950 5466
rect 7962 5414 8014 5466
rect 8026 5414 8078 5466
rect 8090 5414 8142 5466
rect 8154 5414 8206 5466
rect 14846 5414 14898 5466
rect 14910 5414 14962 5466
rect 14974 5414 15026 5466
rect 15038 5414 15090 5466
rect 15102 5414 15154 5466
rect 21794 5414 21846 5466
rect 21858 5414 21910 5466
rect 21922 5414 21974 5466
rect 21986 5414 22038 5466
rect 22050 5414 22102 5466
rect 4424 4870 4476 4922
rect 4488 4870 4540 4922
rect 4552 4870 4604 4922
rect 4616 4870 4668 4922
rect 4680 4870 4732 4922
rect 11372 4870 11424 4922
rect 11436 4870 11488 4922
rect 11500 4870 11552 4922
rect 11564 4870 11616 4922
rect 11628 4870 11680 4922
rect 18320 4870 18372 4922
rect 18384 4870 18436 4922
rect 18448 4870 18500 4922
rect 18512 4870 18564 4922
rect 18576 4870 18628 4922
rect 25268 4870 25320 4922
rect 25332 4870 25384 4922
rect 25396 4870 25448 4922
rect 25460 4870 25512 4922
rect 25524 4870 25576 4922
rect 7898 4326 7950 4378
rect 7962 4326 8014 4378
rect 8026 4326 8078 4378
rect 8090 4326 8142 4378
rect 8154 4326 8206 4378
rect 14846 4326 14898 4378
rect 14910 4326 14962 4378
rect 14974 4326 15026 4378
rect 15038 4326 15090 4378
rect 15102 4326 15154 4378
rect 21794 4326 21846 4378
rect 21858 4326 21910 4378
rect 21922 4326 21974 4378
rect 21986 4326 22038 4378
rect 22050 4326 22102 4378
rect 4424 3782 4476 3834
rect 4488 3782 4540 3834
rect 4552 3782 4604 3834
rect 4616 3782 4668 3834
rect 4680 3782 4732 3834
rect 11372 3782 11424 3834
rect 11436 3782 11488 3834
rect 11500 3782 11552 3834
rect 11564 3782 11616 3834
rect 11628 3782 11680 3834
rect 18320 3782 18372 3834
rect 18384 3782 18436 3834
rect 18448 3782 18500 3834
rect 18512 3782 18564 3834
rect 18576 3782 18628 3834
rect 25268 3782 25320 3834
rect 25332 3782 25384 3834
rect 25396 3782 25448 3834
rect 25460 3782 25512 3834
rect 25524 3782 25576 3834
rect 7898 3238 7950 3290
rect 7962 3238 8014 3290
rect 8026 3238 8078 3290
rect 8090 3238 8142 3290
rect 8154 3238 8206 3290
rect 14846 3238 14898 3290
rect 14910 3238 14962 3290
rect 14974 3238 15026 3290
rect 15038 3238 15090 3290
rect 15102 3238 15154 3290
rect 21794 3238 21846 3290
rect 21858 3238 21910 3290
rect 21922 3238 21974 3290
rect 21986 3238 22038 3290
rect 22050 3238 22102 3290
rect 4424 2694 4476 2746
rect 4488 2694 4540 2746
rect 4552 2694 4604 2746
rect 4616 2694 4668 2746
rect 4680 2694 4732 2746
rect 11372 2694 11424 2746
rect 11436 2694 11488 2746
rect 11500 2694 11552 2746
rect 11564 2694 11616 2746
rect 11628 2694 11680 2746
rect 18320 2694 18372 2746
rect 18384 2694 18436 2746
rect 18448 2694 18500 2746
rect 18512 2694 18564 2746
rect 18576 2694 18628 2746
rect 25268 2694 25320 2746
rect 25332 2694 25384 2746
rect 25396 2694 25448 2746
rect 25460 2694 25512 2746
rect 25524 2694 25576 2746
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 7104 2252 7156 2304
rect 7898 2150 7950 2202
rect 7962 2150 8014 2202
rect 8026 2150 8078 2202
rect 8090 2150 8142 2202
rect 8154 2150 8206 2202
rect 14846 2150 14898 2202
rect 14910 2150 14962 2202
rect 14974 2150 15026 2202
rect 15038 2150 15090 2202
rect 15102 2150 15154 2202
rect 21794 2150 21846 2202
rect 21858 2150 21910 2202
rect 21922 2150 21974 2202
rect 21986 2150 22038 2202
rect 22050 2150 22102 2202
<< metal2 >>
rect 18 29200 74 30000
rect 1306 29200 1362 30000
rect 1950 29200 2006 30000
rect 2594 29200 2650 30000
rect 3882 29200 3938 30000
rect 4526 29200 4582 30000
rect 5814 29200 5870 30000
rect 6458 29200 6514 30000
rect 7746 29200 7802 30000
rect 8390 29200 8446 30000
rect 9034 29200 9090 30000
rect 10322 29200 10378 30000
rect 10966 29200 11022 30000
rect 12254 29200 12310 30000
rect 12898 29200 12954 30000
rect 13542 29200 13598 30000
rect 14830 29200 14886 30000
rect 15474 29200 15530 30000
rect 16118 29200 16174 30000
rect 17406 29200 17462 30000
rect 18050 29200 18106 30000
rect 19338 29200 19394 30000
rect 19982 29200 20038 30000
rect 20626 29200 20682 30000
rect 21914 29200 21970 30000
rect 22558 29200 22614 30000
rect 23846 29200 23902 30000
rect 24490 29200 24546 30000
rect 25134 29200 25190 30000
rect 26422 29200 26478 30000
rect 27066 29200 27122 30000
rect 28354 29200 28410 30000
rect 28998 29200 29054 30000
rect 29642 29200 29698 30000
rect 4424 27772 4732 27781
rect 4424 27770 4430 27772
rect 4486 27770 4510 27772
rect 4566 27770 4590 27772
rect 4646 27770 4670 27772
rect 4726 27770 4732 27772
rect 4486 27718 4488 27770
rect 4668 27718 4670 27770
rect 4424 27716 4430 27718
rect 4486 27716 4510 27718
rect 4566 27716 4590 27718
rect 4646 27716 4670 27718
rect 4726 27716 4732 27718
rect 4424 27707 4732 27716
rect 11372 27772 11680 27781
rect 11372 27770 11378 27772
rect 11434 27770 11458 27772
rect 11514 27770 11538 27772
rect 11594 27770 11618 27772
rect 11674 27770 11680 27772
rect 11434 27718 11436 27770
rect 11616 27718 11618 27770
rect 11372 27716 11378 27718
rect 11434 27716 11458 27718
rect 11514 27716 11538 27718
rect 11594 27716 11618 27718
rect 11674 27716 11680 27718
rect 11372 27707 11680 27716
rect 18320 27772 18628 27781
rect 18320 27770 18326 27772
rect 18382 27770 18406 27772
rect 18462 27770 18486 27772
rect 18542 27770 18566 27772
rect 18622 27770 18628 27772
rect 18382 27718 18384 27770
rect 18564 27718 18566 27770
rect 18320 27716 18326 27718
rect 18382 27716 18406 27718
rect 18462 27716 18486 27718
rect 18542 27716 18566 27718
rect 18622 27716 18628 27718
rect 18320 27707 18628 27716
rect 25268 27772 25576 27781
rect 25268 27770 25274 27772
rect 25330 27770 25354 27772
rect 25410 27770 25434 27772
rect 25490 27770 25514 27772
rect 25570 27770 25576 27772
rect 25330 27718 25332 27770
rect 25512 27718 25514 27770
rect 25268 27716 25274 27718
rect 25330 27716 25354 27718
rect 25410 27716 25434 27718
rect 25490 27716 25514 27718
rect 25570 27716 25576 27718
rect 25268 27707 25576 27716
rect 7898 27228 8206 27237
rect 7898 27226 7904 27228
rect 7960 27226 7984 27228
rect 8040 27226 8064 27228
rect 8120 27226 8144 27228
rect 8200 27226 8206 27228
rect 7960 27174 7962 27226
rect 8142 27174 8144 27226
rect 7898 27172 7904 27174
rect 7960 27172 7984 27174
rect 8040 27172 8064 27174
rect 8120 27172 8144 27174
rect 8200 27172 8206 27174
rect 7898 27163 8206 27172
rect 14846 27228 15154 27237
rect 14846 27226 14852 27228
rect 14908 27226 14932 27228
rect 14988 27226 15012 27228
rect 15068 27226 15092 27228
rect 15148 27226 15154 27228
rect 14908 27174 14910 27226
rect 15090 27174 15092 27226
rect 14846 27172 14852 27174
rect 14908 27172 14932 27174
rect 14988 27172 15012 27174
rect 15068 27172 15092 27174
rect 15148 27172 15154 27174
rect 14846 27163 15154 27172
rect 21794 27228 22102 27237
rect 21794 27226 21800 27228
rect 21856 27226 21880 27228
rect 21936 27226 21960 27228
rect 22016 27226 22040 27228
rect 22096 27226 22102 27228
rect 21856 27174 21858 27226
rect 22038 27174 22040 27226
rect 21794 27172 21800 27174
rect 21856 27172 21880 27174
rect 21936 27172 21960 27174
rect 22016 27172 22040 27174
rect 22096 27172 22102 27174
rect 21794 27163 22102 27172
rect 4424 26684 4732 26693
rect 4424 26682 4430 26684
rect 4486 26682 4510 26684
rect 4566 26682 4590 26684
rect 4646 26682 4670 26684
rect 4726 26682 4732 26684
rect 4486 26630 4488 26682
rect 4668 26630 4670 26682
rect 4424 26628 4430 26630
rect 4486 26628 4510 26630
rect 4566 26628 4590 26630
rect 4646 26628 4670 26630
rect 4726 26628 4732 26630
rect 4424 26619 4732 26628
rect 11372 26684 11680 26693
rect 11372 26682 11378 26684
rect 11434 26682 11458 26684
rect 11514 26682 11538 26684
rect 11594 26682 11618 26684
rect 11674 26682 11680 26684
rect 11434 26630 11436 26682
rect 11616 26630 11618 26682
rect 11372 26628 11378 26630
rect 11434 26628 11458 26630
rect 11514 26628 11538 26630
rect 11594 26628 11618 26630
rect 11674 26628 11680 26630
rect 11372 26619 11680 26628
rect 18320 26684 18628 26693
rect 18320 26682 18326 26684
rect 18382 26682 18406 26684
rect 18462 26682 18486 26684
rect 18542 26682 18566 26684
rect 18622 26682 18628 26684
rect 18382 26630 18384 26682
rect 18564 26630 18566 26682
rect 18320 26628 18326 26630
rect 18382 26628 18406 26630
rect 18462 26628 18486 26630
rect 18542 26628 18566 26630
rect 18622 26628 18628 26630
rect 18320 26619 18628 26628
rect 25268 26684 25576 26693
rect 25268 26682 25274 26684
rect 25330 26682 25354 26684
rect 25410 26682 25434 26684
rect 25490 26682 25514 26684
rect 25570 26682 25576 26684
rect 25330 26630 25332 26682
rect 25512 26630 25514 26682
rect 25268 26628 25274 26630
rect 25330 26628 25354 26630
rect 25410 26628 25434 26630
rect 25490 26628 25514 26630
rect 25570 26628 25576 26630
rect 25268 26619 25576 26628
rect 7898 26140 8206 26149
rect 7898 26138 7904 26140
rect 7960 26138 7984 26140
rect 8040 26138 8064 26140
rect 8120 26138 8144 26140
rect 8200 26138 8206 26140
rect 7960 26086 7962 26138
rect 8142 26086 8144 26138
rect 7898 26084 7904 26086
rect 7960 26084 7984 26086
rect 8040 26084 8064 26086
rect 8120 26084 8144 26086
rect 8200 26084 8206 26086
rect 7898 26075 8206 26084
rect 14846 26140 15154 26149
rect 14846 26138 14852 26140
rect 14908 26138 14932 26140
rect 14988 26138 15012 26140
rect 15068 26138 15092 26140
rect 15148 26138 15154 26140
rect 14908 26086 14910 26138
rect 15090 26086 15092 26138
rect 14846 26084 14852 26086
rect 14908 26084 14932 26086
rect 14988 26084 15012 26086
rect 15068 26084 15092 26086
rect 15148 26084 15154 26086
rect 14846 26075 15154 26084
rect 21794 26140 22102 26149
rect 21794 26138 21800 26140
rect 21856 26138 21880 26140
rect 21936 26138 21960 26140
rect 22016 26138 22040 26140
rect 22096 26138 22102 26140
rect 21856 26086 21858 26138
rect 22038 26086 22040 26138
rect 21794 26084 21800 26086
rect 21856 26084 21880 26086
rect 21936 26084 21960 26086
rect 22016 26084 22040 26086
rect 22096 26084 22102 26086
rect 21794 26075 22102 26084
rect 4424 25596 4732 25605
rect 4424 25594 4430 25596
rect 4486 25594 4510 25596
rect 4566 25594 4590 25596
rect 4646 25594 4670 25596
rect 4726 25594 4732 25596
rect 4486 25542 4488 25594
rect 4668 25542 4670 25594
rect 4424 25540 4430 25542
rect 4486 25540 4510 25542
rect 4566 25540 4590 25542
rect 4646 25540 4670 25542
rect 4726 25540 4732 25542
rect 4424 25531 4732 25540
rect 11372 25596 11680 25605
rect 11372 25594 11378 25596
rect 11434 25594 11458 25596
rect 11514 25594 11538 25596
rect 11594 25594 11618 25596
rect 11674 25594 11680 25596
rect 11434 25542 11436 25594
rect 11616 25542 11618 25594
rect 11372 25540 11378 25542
rect 11434 25540 11458 25542
rect 11514 25540 11538 25542
rect 11594 25540 11618 25542
rect 11674 25540 11680 25542
rect 11372 25531 11680 25540
rect 18320 25596 18628 25605
rect 18320 25594 18326 25596
rect 18382 25594 18406 25596
rect 18462 25594 18486 25596
rect 18542 25594 18566 25596
rect 18622 25594 18628 25596
rect 18382 25542 18384 25594
rect 18564 25542 18566 25594
rect 18320 25540 18326 25542
rect 18382 25540 18406 25542
rect 18462 25540 18486 25542
rect 18542 25540 18566 25542
rect 18622 25540 18628 25542
rect 18320 25531 18628 25540
rect 25268 25596 25576 25605
rect 25268 25594 25274 25596
rect 25330 25594 25354 25596
rect 25410 25594 25434 25596
rect 25490 25594 25514 25596
rect 25570 25594 25576 25596
rect 25330 25542 25332 25594
rect 25512 25542 25514 25594
rect 25268 25540 25274 25542
rect 25330 25540 25354 25542
rect 25410 25540 25434 25542
rect 25490 25540 25514 25542
rect 25570 25540 25576 25542
rect 25268 25531 25576 25540
rect 7898 25052 8206 25061
rect 7898 25050 7904 25052
rect 7960 25050 7984 25052
rect 8040 25050 8064 25052
rect 8120 25050 8144 25052
rect 8200 25050 8206 25052
rect 7960 24998 7962 25050
rect 8142 24998 8144 25050
rect 7898 24996 7904 24998
rect 7960 24996 7984 24998
rect 8040 24996 8064 24998
rect 8120 24996 8144 24998
rect 8200 24996 8206 24998
rect 7898 24987 8206 24996
rect 14846 25052 15154 25061
rect 14846 25050 14852 25052
rect 14908 25050 14932 25052
rect 14988 25050 15012 25052
rect 15068 25050 15092 25052
rect 15148 25050 15154 25052
rect 14908 24998 14910 25050
rect 15090 24998 15092 25050
rect 14846 24996 14852 24998
rect 14908 24996 14932 24998
rect 14988 24996 15012 24998
rect 15068 24996 15092 24998
rect 15148 24996 15154 24998
rect 14846 24987 15154 24996
rect 21794 25052 22102 25061
rect 21794 25050 21800 25052
rect 21856 25050 21880 25052
rect 21936 25050 21960 25052
rect 22016 25050 22040 25052
rect 22096 25050 22102 25052
rect 21856 24998 21858 25050
rect 22038 24998 22040 25050
rect 21794 24996 21800 24998
rect 21856 24996 21880 24998
rect 21936 24996 21960 24998
rect 22016 24996 22040 24998
rect 22096 24996 22102 24998
rect 21794 24987 22102 24996
rect 4424 24508 4732 24517
rect 4424 24506 4430 24508
rect 4486 24506 4510 24508
rect 4566 24506 4590 24508
rect 4646 24506 4670 24508
rect 4726 24506 4732 24508
rect 4486 24454 4488 24506
rect 4668 24454 4670 24506
rect 4424 24452 4430 24454
rect 4486 24452 4510 24454
rect 4566 24452 4590 24454
rect 4646 24452 4670 24454
rect 4726 24452 4732 24454
rect 4424 24443 4732 24452
rect 11372 24508 11680 24517
rect 11372 24506 11378 24508
rect 11434 24506 11458 24508
rect 11514 24506 11538 24508
rect 11594 24506 11618 24508
rect 11674 24506 11680 24508
rect 11434 24454 11436 24506
rect 11616 24454 11618 24506
rect 11372 24452 11378 24454
rect 11434 24452 11458 24454
rect 11514 24452 11538 24454
rect 11594 24452 11618 24454
rect 11674 24452 11680 24454
rect 11372 24443 11680 24452
rect 18320 24508 18628 24517
rect 18320 24506 18326 24508
rect 18382 24506 18406 24508
rect 18462 24506 18486 24508
rect 18542 24506 18566 24508
rect 18622 24506 18628 24508
rect 18382 24454 18384 24506
rect 18564 24454 18566 24506
rect 18320 24452 18326 24454
rect 18382 24452 18406 24454
rect 18462 24452 18486 24454
rect 18542 24452 18566 24454
rect 18622 24452 18628 24454
rect 18320 24443 18628 24452
rect 25268 24508 25576 24517
rect 25268 24506 25274 24508
rect 25330 24506 25354 24508
rect 25410 24506 25434 24508
rect 25490 24506 25514 24508
rect 25570 24506 25576 24508
rect 25330 24454 25332 24506
rect 25512 24454 25514 24506
rect 25268 24452 25274 24454
rect 25330 24452 25354 24454
rect 25410 24452 25434 24454
rect 25490 24452 25514 24454
rect 25570 24452 25576 24454
rect 25268 24443 25576 24452
rect 7898 23964 8206 23973
rect 7898 23962 7904 23964
rect 7960 23962 7984 23964
rect 8040 23962 8064 23964
rect 8120 23962 8144 23964
rect 8200 23962 8206 23964
rect 7960 23910 7962 23962
rect 8142 23910 8144 23962
rect 7898 23908 7904 23910
rect 7960 23908 7984 23910
rect 8040 23908 8064 23910
rect 8120 23908 8144 23910
rect 8200 23908 8206 23910
rect 7898 23899 8206 23908
rect 14846 23964 15154 23973
rect 14846 23962 14852 23964
rect 14908 23962 14932 23964
rect 14988 23962 15012 23964
rect 15068 23962 15092 23964
rect 15148 23962 15154 23964
rect 14908 23910 14910 23962
rect 15090 23910 15092 23962
rect 14846 23908 14852 23910
rect 14908 23908 14932 23910
rect 14988 23908 15012 23910
rect 15068 23908 15092 23910
rect 15148 23908 15154 23910
rect 14846 23899 15154 23908
rect 21794 23964 22102 23973
rect 21794 23962 21800 23964
rect 21856 23962 21880 23964
rect 21936 23962 21960 23964
rect 22016 23962 22040 23964
rect 22096 23962 22102 23964
rect 21856 23910 21858 23962
rect 22038 23910 22040 23962
rect 21794 23908 21800 23910
rect 21856 23908 21880 23910
rect 21936 23908 21960 23910
rect 22016 23908 22040 23910
rect 22096 23908 22102 23910
rect 21794 23899 22102 23908
rect 4424 23420 4732 23429
rect 4424 23418 4430 23420
rect 4486 23418 4510 23420
rect 4566 23418 4590 23420
rect 4646 23418 4670 23420
rect 4726 23418 4732 23420
rect 4486 23366 4488 23418
rect 4668 23366 4670 23418
rect 4424 23364 4430 23366
rect 4486 23364 4510 23366
rect 4566 23364 4590 23366
rect 4646 23364 4670 23366
rect 4726 23364 4732 23366
rect 4424 23355 4732 23364
rect 11372 23420 11680 23429
rect 11372 23418 11378 23420
rect 11434 23418 11458 23420
rect 11514 23418 11538 23420
rect 11594 23418 11618 23420
rect 11674 23418 11680 23420
rect 11434 23366 11436 23418
rect 11616 23366 11618 23418
rect 11372 23364 11378 23366
rect 11434 23364 11458 23366
rect 11514 23364 11538 23366
rect 11594 23364 11618 23366
rect 11674 23364 11680 23366
rect 11372 23355 11680 23364
rect 18320 23420 18628 23429
rect 18320 23418 18326 23420
rect 18382 23418 18406 23420
rect 18462 23418 18486 23420
rect 18542 23418 18566 23420
rect 18622 23418 18628 23420
rect 18382 23366 18384 23418
rect 18564 23366 18566 23418
rect 18320 23364 18326 23366
rect 18382 23364 18406 23366
rect 18462 23364 18486 23366
rect 18542 23364 18566 23366
rect 18622 23364 18628 23366
rect 18320 23355 18628 23364
rect 25268 23420 25576 23429
rect 25268 23418 25274 23420
rect 25330 23418 25354 23420
rect 25410 23418 25434 23420
rect 25490 23418 25514 23420
rect 25570 23418 25576 23420
rect 25330 23366 25332 23418
rect 25512 23366 25514 23418
rect 25268 23364 25274 23366
rect 25330 23364 25354 23366
rect 25410 23364 25434 23366
rect 25490 23364 25514 23366
rect 25570 23364 25576 23366
rect 25268 23355 25576 23364
rect 7898 22876 8206 22885
rect 7898 22874 7904 22876
rect 7960 22874 7984 22876
rect 8040 22874 8064 22876
rect 8120 22874 8144 22876
rect 8200 22874 8206 22876
rect 7960 22822 7962 22874
rect 8142 22822 8144 22874
rect 7898 22820 7904 22822
rect 7960 22820 7984 22822
rect 8040 22820 8064 22822
rect 8120 22820 8144 22822
rect 8200 22820 8206 22822
rect 7898 22811 8206 22820
rect 14846 22876 15154 22885
rect 14846 22874 14852 22876
rect 14908 22874 14932 22876
rect 14988 22874 15012 22876
rect 15068 22874 15092 22876
rect 15148 22874 15154 22876
rect 14908 22822 14910 22874
rect 15090 22822 15092 22874
rect 14846 22820 14852 22822
rect 14908 22820 14932 22822
rect 14988 22820 15012 22822
rect 15068 22820 15092 22822
rect 15148 22820 15154 22822
rect 14846 22811 15154 22820
rect 21794 22876 22102 22885
rect 21794 22874 21800 22876
rect 21856 22874 21880 22876
rect 21936 22874 21960 22876
rect 22016 22874 22040 22876
rect 22096 22874 22102 22876
rect 21856 22822 21858 22874
rect 22038 22822 22040 22874
rect 21794 22820 21800 22822
rect 21856 22820 21880 22822
rect 21936 22820 21960 22822
rect 22016 22820 22040 22822
rect 22096 22820 22102 22822
rect 21794 22811 22102 22820
rect 4424 22332 4732 22341
rect 4424 22330 4430 22332
rect 4486 22330 4510 22332
rect 4566 22330 4590 22332
rect 4646 22330 4670 22332
rect 4726 22330 4732 22332
rect 4486 22278 4488 22330
rect 4668 22278 4670 22330
rect 4424 22276 4430 22278
rect 4486 22276 4510 22278
rect 4566 22276 4590 22278
rect 4646 22276 4670 22278
rect 4726 22276 4732 22278
rect 4424 22267 4732 22276
rect 11372 22332 11680 22341
rect 11372 22330 11378 22332
rect 11434 22330 11458 22332
rect 11514 22330 11538 22332
rect 11594 22330 11618 22332
rect 11674 22330 11680 22332
rect 11434 22278 11436 22330
rect 11616 22278 11618 22330
rect 11372 22276 11378 22278
rect 11434 22276 11458 22278
rect 11514 22276 11538 22278
rect 11594 22276 11618 22278
rect 11674 22276 11680 22278
rect 11372 22267 11680 22276
rect 18320 22332 18628 22341
rect 18320 22330 18326 22332
rect 18382 22330 18406 22332
rect 18462 22330 18486 22332
rect 18542 22330 18566 22332
rect 18622 22330 18628 22332
rect 18382 22278 18384 22330
rect 18564 22278 18566 22330
rect 18320 22276 18326 22278
rect 18382 22276 18406 22278
rect 18462 22276 18486 22278
rect 18542 22276 18566 22278
rect 18622 22276 18628 22278
rect 18320 22267 18628 22276
rect 25268 22332 25576 22341
rect 25268 22330 25274 22332
rect 25330 22330 25354 22332
rect 25410 22330 25434 22332
rect 25490 22330 25514 22332
rect 25570 22330 25576 22332
rect 25330 22278 25332 22330
rect 25512 22278 25514 22330
rect 25268 22276 25274 22278
rect 25330 22276 25354 22278
rect 25410 22276 25434 22278
rect 25490 22276 25514 22278
rect 25570 22276 25576 22278
rect 25268 22267 25576 22276
rect 7898 21788 8206 21797
rect 7898 21786 7904 21788
rect 7960 21786 7984 21788
rect 8040 21786 8064 21788
rect 8120 21786 8144 21788
rect 8200 21786 8206 21788
rect 7960 21734 7962 21786
rect 8142 21734 8144 21786
rect 7898 21732 7904 21734
rect 7960 21732 7984 21734
rect 8040 21732 8064 21734
rect 8120 21732 8144 21734
rect 8200 21732 8206 21734
rect 7898 21723 8206 21732
rect 14846 21788 15154 21797
rect 14846 21786 14852 21788
rect 14908 21786 14932 21788
rect 14988 21786 15012 21788
rect 15068 21786 15092 21788
rect 15148 21786 15154 21788
rect 14908 21734 14910 21786
rect 15090 21734 15092 21786
rect 14846 21732 14852 21734
rect 14908 21732 14932 21734
rect 14988 21732 15012 21734
rect 15068 21732 15092 21734
rect 15148 21732 15154 21734
rect 14846 21723 15154 21732
rect 21794 21788 22102 21797
rect 21794 21786 21800 21788
rect 21856 21786 21880 21788
rect 21936 21786 21960 21788
rect 22016 21786 22040 21788
rect 22096 21786 22102 21788
rect 21856 21734 21858 21786
rect 22038 21734 22040 21786
rect 21794 21732 21800 21734
rect 21856 21732 21880 21734
rect 21936 21732 21960 21734
rect 22016 21732 22040 21734
rect 22096 21732 22102 21734
rect 21794 21723 22102 21732
rect 4424 21244 4732 21253
rect 4424 21242 4430 21244
rect 4486 21242 4510 21244
rect 4566 21242 4590 21244
rect 4646 21242 4670 21244
rect 4726 21242 4732 21244
rect 4486 21190 4488 21242
rect 4668 21190 4670 21242
rect 4424 21188 4430 21190
rect 4486 21188 4510 21190
rect 4566 21188 4590 21190
rect 4646 21188 4670 21190
rect 4726 21188 4732 21190
rect 4424 21179 4732 21188
rect 11372 21244 11680 21253
rect 11372 21242 11378 21244
rect 11434 21242 11458 21244
rect 11514 21242 11538 21244
rect 11594 21242 11618 21244
rect 11674 21242 11680 21244
rect 11434 21190 11436 21242
rect 11616 21190 11618 21242
rect 11372 21188 11378 21190
rect 11434 21188 11458 21190
rect 11514 21188 11538 21190
rect 11594 21188 11618 21190
rect 11674 21188 11680 21190
rect 11372 21179 11680 21188
rect 18320 21244 18628 21253
rect 18320 21242 18326 21244
rect 18382 21242 18406 21244
rect 18462 21242 18486 21244
rect 18542 21242 18566 21244
rect 18622 21242 18628 21244
rect 18382 21190 18384 21242
rect 18564 21190 18566 21242
rect 18320 21188 18326 21190
rect 18382 21188 18406 21190
rect 18462 21188 18486 21190
rect 18542 21188 18566 21190
rect 18622 21188 18628 21190
rect 18320 21179 18628 21188
rect 25268 21244 25576 21253
rect 25268 21242 25274 21244
rect 25330 21242 25354 21244
rect 25410 21242 25434 21244
rect 25490 21242 25514 21244
rect 25570 21242 25576 21244
rect 25330 21190 25332 21242
rect 25512 21190 25514 21242
rect 25268 21188 25274 21190
rect 25330 21188 25354 21190
rect 25410 21188 25434 21190
rect 25490 21188 25514 21190
rect 25570 21188 25576 21190
rect 25268 21179 25576 21188
rect 7898 20700 8206 20709
rect 7898 20698 7904 20700
rect 7960 20698 7984 20700
rect 8040 20698 8064 20700
rect 8120 20698 8144 20700
rect 8200 20698 8206 20700
rect 7960 20646 7962 20698
rect 8142 20646 8144 20698
rect 7898 20644 7904 20646
rect 7960 20644 7984 20646
rect 8040 20644 8064 20646
rect 8120 20644 8144 20646
rect 8200 20644 8206 20646
rect 7898 20635 8206 20644
rect 14846 20700 15154 20709
rect 14846 20698 14852 20700
rect 14908 20698 14932 20700
rect 14988 20698 15012 20700
rect 15068 20698 15092 20700
rect 15148 20698 15154 20700
rect 14908 20646 14910 20698
rect 15090 20646 15092 20698
rect 14846 20644 14852 20646
rect 14908 20644 14932 20646
rect 14988 20644 15012 20646
rect 15068 20644 15092 20646
rect 15148 20644 15154 20646
rect 14846 20635 15154 20644
rect 21794 20700 22102 20709
rect 21794 20698 21800 20700
rect 21856 20698 21880 20700
rect 21936 20698 21960 20700
rect 22016 20698 22040 20700
rect 22096 20698 22102 20700
rect 21856 20646 21858 20698
rect 22038 20646 22040 20698
rect 21794 20644 21800 20646
rect 21856 20644 21880 20646
rect 21936 20644 21960 20646
rect 22016 20644 22040 20646
rect 22096 20644 22102 20646
rect 21794 20635 22102 20644
rect 4424 20156 4732 20165
rect 4424 20154 4430 20156
rect 4486 20154 4510 20156
rect 4566 20154 4590 20156
rect 4646 20154 4670 20156
rect 4726 20154 4732 20156
rect 4486 20102 4488 20154
rect 4668 20102 4670 20154
rect 4424 20100 4430 20102
rect 4486 20100 4510 20102
rect 4566 20100 4590 20102
rect 4646 20100 4670 20102
rect 4726 20100 4732 20102
rect 4424 20091 4732 20100
rect 11372 20156 11680 20165
rect 11372 20154 11378 20156
rect 11434 20154 11458 20156
rect 11514 20154 11538 20156
rect 11594 20154 11618 20156
rect 11674 20154 11680 20156
rect 11434 20102 11436 20154
rect 11616 20102 11618 20154
rect 11372 20100 11378 20102
rect 11434 20100 11458 20102
rect 11514 20100 11538 20102
rect 11594 20100 11618 20102
rect 11674 20100 11680 20102
rect 11372 20091 11680 20100
rect 18320 20156 18628 20165
rect 18320 20154 18326 20156
rect 18382 20154 18406 20156
rect 18462 20154 18486 20156
rect 18542 20154 18566 20156
rect 18622 20154 18628 20156
rect 18382 20102 18384 20154
rect 18564 20102 18566 20154
rect 18320 20100 18326 20102
rect 18382 20100 18406 20102
rect 18462 20100 18486 20102
rect 18542 20100 18566 20102
rect 18622 20100 18628 20102
rect 18320 20091 18628 20100
rect 25268 20156 25576 20165
rect 25268 20154 25274 20156
rect 25330 20154 25354 20156
rect 25410 20154 25434 20156
rect 25490 20154 25514 20156
rect 25570 20154 25576 20156
rect 25330 20102 25332 20154
rect 25512 20102 25514 20154
rect 25268 20100 25274 20102
rect 25330 20100 25354 20102
rect 25410 20100 25434 20102
rect 25490 20100 25514 20102
rect 25570 20100 25576 20102
rect 25268 20091 25576 20100
rect 7898 19612 8206 19621
rect 7898 19610 7904 19612
rect 7960 19610 7984 19612
rect 8040 19610 8064 19612
rect 8120 19610 8144 19612
rect 8200 19610 8206 19612
rect 7960 19558 7962 19610
rect 8142 19558 8144 19610
rect 7898 19556 7904 19558
rect 7960 19556 7984 19558
rect 8040 19556 8064 19558
rect 8120 19556 8144 19558
rect 8200 19556 8206 19558
rect 7898 19547 8206 19556
rect 14846 19612 15154 19621
rect 14846 19610 14852 19612
rect 14908 19610 14932 19612
rect 14988 19610 15012 19612
rect 15068 19610 15092 19612
rect 15148 19610 15154 19612
rect 14908 19558 14910 19610
rect 15090 19558 15092 19610
rect 14846 19556 14852 19558
rect 14908 19556 14932 19558
rect 14988 19556 15012 19558
rect 15068 19556 15092 19558
rect 15148 19556 15154 19558
rect 14846 19547 15154 19556
rect 21794 19612 22102 19621
rect 21794 19610 21800 19612
rect 21856 19610 21880 19612
rect 21936 19610 21960 19612
rect 22016 19610 22040 19612
rect 22096 19610 22102 19612
rect 21856 19558 21858 19610
rect 22038 19558 22040 19610
rect 21794 19556 21800 19558
rect 21856 19556 21880 19558
rect 21936 19556 21960 19558
rect 22016 19556 22040 19558
rect 22096 19556 22102 19558
rect 21794 19547 22102 19556
rect 4424 19068 4732 19077
rect 4424 19066 4430 19068
rect 4486 19066 4510 19068
rect 4566 19066 4590 19068
rect 4646 19066 4670 19068
rect 4726 19066 4732 19068
rect 4486 19014 4488 19066
rect 4668 19014 4670 19066
rect 4424 19012 4430 19014
rect 4486 19012 4510 19014
rect 4566 19012 4590 19014
rect 4646 19012 4670 19014
rect 4726 19012 4732 19014
rect 4424 19003 4732 19012
rect 11372 19068 11680 19077
rect 11372 19066 11378 19068
rect 11434 19066 11458 19068
rect 11514 19066 11538 19068
rect 11594 19066 11618 19068
rect 11674 19066 11680 19068
rect 11434 19014 11436 19066
rect 11616 19014 11618 19066
rect 11372 19012 11378 19014
rect 11434 19012 11458 19014
rect 11514 19012 11538 19014
rect 11594 19012 11618 19014
rect 11674 19012 11680 19014
rect 11372 19003 11680 19012
rect 18320 19068 18628 19077
rect 18320 19066 18326 19068
rect 18382 19066 18406 19068
rect 18462 19066 18486 19068
rect 18542 19066 18566 19068
rect 18622 19066 18628 19068
rect 18382 19014 18384 19066
rect 18564 19014 18566 19066
rect 18320 19012 18326 19014
rect 18382 19012 18406 19014
rect 18462 19012 18486 19014
rect 18542 19012 18566 19014
rect 18622 19012 18628 19014
rect 18320 19003 18628 19012
rect 25268 19068 25576 19077
rect 25268 19066 25274 19068
rect 25330 19066 25354 19068
rect 25410 19066 25434 19068
rect 25490 19066 25514 19068
rect 25570 19066 25576 19068
rect 25330 19014 25332 19066
rect 25512 19014 25514 19066
rect 25268 19012 25274 19014
rect 25330 19012 25354 19014
rect 25410 19012 25434 19014
rect 25490 19012 25514 19014
rect 25570 19012 25576 19014
rect 25268 19003 25576 19012
rect 7898 18524 8206 18533
rect 7898 18522 7904 18524
rect 7960 18522 7984 18524
rect 8040 18522 8064 18524
rect 8120 18522 8144 18524
rect 8200 18522 8206 18524
rect 7960 18470 7962 18522
rect 8142 18470 8144 18522
rect 7898 18468 7904 18470
rect 7960 18468 7984 18470
rect 8040 18468 8064 18470
rect 8120 18468 8144 18470
rect 8200 18468 8206 18470
rect 7898 18459 8206 18468
rect 14846 18524 15154 18533
rect 14846 18522 14852 18524
rect 14908 18522 14932 18524
rect 14988 18522 15012 18524
rect 15068 18522 15092 18524
rect 15148 18522 15154 18524
rect 14908 18470 14910 18522
rect 15090 18470 15092 18522
rect 14846 18468 14852 18470
rect 14908 18468 14932 18470
rect 14988 18468 15012 18470
rect 15068 18468 15092 18470
rect 15148 18468 15154 18470
rect 14846 18459 15154 18468
rect 21794 18524 22102 18533
rect 21794 18522 21800 18524
rect 21856 18522 21880 18524
rect 21936 18522 21960 18524
rect 22016 18522 22040 18524
rect 22096 18522 22102 18524
rect 21856 18470 21858 18522
rect 22038 18470 22040 18522
rect 21794 18468 21800 18470
rect 21856 18468 21880 18470
rect 21936 18468 21960 18470
rect 22016 18468 22040 18470
rect 22096 18468 22102 18470
rect 21794 18459 22102 18468
rect 4424 17980 4732 17989
rect 4424 17978 4430 17980
rect 4486 17978 4510 17980
rect 4566 17978 4590 17980
rect 4646 17978 4670 17980
rect 4726 17978 4732 17980
rect 4486 17926 4488 17978
rect 4668 17926 4670 17978
rect 4424 17924 4430 17926
rect 4486 17924 4510 17926
rect 4566 17924 4590 17926
rect 4646 17924 4670 17926
rect 4726 17924 4732 17926
rect 4424 17915 4732 17924
rect 11372 17980 11680 17989
rect 11372 17978 11378 17980
rect 11434 17978 11458 17980
rect 11514 17978 11538 17980
rect 11594 17978 11618 17980
rect 11674 17978 11680 17980
rect 11434 17926 11436 17978
rect 11616 17926 11618 17978
rect 11372 17924 11378 17926
rect 11434 17924 11458 17926
rect 11514 17924 11538 17926
rect 11594 17924 11618 17926
rect 11674 17924 11680 17926
rect 11372 17915 11680 17924
rect 18320 17980 18628 17989
rect 18320 17978 18326 17980
rect 18382 17978 18406 17980
rect 18462 17978 18486 17980
rect 18542 17978 18566 17980
rect 18622 17978 18628 17980
rect 18382 17926 18384 17978
rect 18564 17926 18566 17978
rect 18320 17924 18326 17926
rect 18382 17924 18406 17926
rect 18462 17924 18486 17926
rect 18542 17924 18566 17926
rect 18622 17924 18628 17926
rect 18320 17915 18628 17924
rect 25268 17980 25576 17989
rect 25268 17978 25274 17980
rect 25330 17978 25354 17980
rect 25410 17978 25434 17980
rect 25490 17978 25514 17980
rect 25570 17978 25576 17980
rect 25330 17926 25332 17978
rect 25512 17926 25514 17978
rect 25268 17924 25274 17926
rect 25330 17924 25354 17926
rect 25410 17924 25434 17926
rect 25490 17924 25514 17926
rect 25570 17924 25576 17926
rect 25268 17915 25576 17924
rect 7898 17436 8206 17445
rect 7898 17434 7904 17436
rect 7960 17434 7984 17436
rect 8040 17434 8064 17436
rect 8120 17434 8144 17436
rect 8200 17434 8206 17436
rect 7960 17382 7962 17434
rect 8142 17382 8144 17434
rect 7898 17380 7904 17382
rect 7960 17380 7984 17382
rect 8040 17380 8064 17382
rect 8120 17380 8144 17382
rect 8200 17380 8206 17382
rect 7898 17371 8206 17380
rect 14846 17436 15154 17445
rect 14846 17434 14852 17436
rect 14908 17434 14932 17436
rect 14988 17434 15012 17436
rect 15068 17434 15092 17436
rect 15148 17434 15154 17436
rect 14908 17382 14910 17434
rect 15090 17382 15092 17434
rect 14846 17380 14852 17382
rect 14908 17380 14932 17382
rect 14988 17380 15012 17382
rect 15068 17380 15092 17382
rect 15148 17380 15154 17382
rect 14846 17371 15154 17380
rect 21794 17436 22102 17445
rect 21794 17434 21800 17436
rect 21856 17434 21880 17436
rect 21936 17434 21960 17436
rect 22016 17434 22040 17436
rect 22096 17434 22102 17436
rect 21856 17382 21858 17434
rect 22038 17382 22040 17434
rect 21794 17380 21800 17382
rect 21856 17380 21880 17382
rect 21936 17380 21960 17382
rect 22016 17380 22040 17382
rect 22096 17380 22102 17382
rect 21794 17371 22102 17380
rect 4424 16892 4732 16901
rect 4424 16890 4430 16892
rect 4486 16890 4510 16892
rect 4566 16890 4590 16892
rect 4646 16890 4670 16892
rect 4726 16890 4732 16892
rect 4486 16838 4488 16890
rect 4668 16838 4670 16890
rect 4424 16836 4430 16838
rect 4486 16836 4510 16838
rect 4566 16836 4590 16838
rect 4646 16836 4670 16838
rect 4726 16836 4732 16838
rect 4424 16827 4732 16836
rect 11372 16892 11680 16901
rect 11372 16890 11378 16892
rect 11434 16890 11458 16892
rect 11514 16890 11538 16892
rect 11594 16890 11618 16892
rect 11674 16890 11680 16892
rect 11434 16838 11436 16890
rect 11616 16838 11618 16890
rect 11372 16836 11378 16838
rect 11434 16836 11458 16838
rect 11514 16836 11538 16838
rect 11594 16836 11618 16838
rect 11674 16836 11680 16838
rect 11372 16827 11680 16836
rect 18320 16892 18628 16901
rect 18320 16890 18326 16892
rect 18382 16890 18406 16892
rect 18462 16890 18486 16892
rect 18542 16890 18566 16892
rect 18622 16890 18628 16892
rect 18382 16838 18384 16890
rect 18564 16838 18566 16890
rect 18320 16836 18326 16838
rect 18382 16836 18406 16838
rect 18462 16836 18486 16838
rect 18542 16836 18566 16838
rect 18622 16836 18628 16838
rect 18320 16827 18628 16836
rect 25268 16892 25576 16901
rect 25268 16890 25274 16892
rect 25330 16890 25354 16892
rect 25410 16890 25434 16892
rect 25490 16890 25514 16892
rect 25570 16890 25576 16892
rect 25330 16838 25332 16890
rect 25512 16838 25514 16890
rect 25268 16836 25274 16838
rect 25330 16836 25354 16838
rect 25410 16836 25434 16838
rect 25490 16836 25514 16838
rect 25570 16836 25576 16838
rect 25268 16827 25576 16836
rect 7898 16348 8206 16357
rect 7898 16346 7904 16348
rect 7960 16346 7984 16348
rect 8040 16346 8064 16348
rect 8120 16346 8144 16348
rect 8200 16346 8206 16348
rect 7960 16294 7962 16346
rect 8142 16294 8144 16346
rect 7898 16292 7904 16294
rect 7960 16292 7984 16294
rect 8040 16292 8064 16294
rect 8120 16292 8144 16294
rect 8200 16292 8206 16294
rect 7898 16283 8206 16292
rect 14846 16348 15154 16357
rect 14846 16346 14852 16348
rect 14908 16346 14932 16348
rect 14988 16346 15012 16348
rect 15068 16346 15092 16348
rect 15148 16346 15154 16348
rect 14908 16294 14910 16346
rect 15090 16294 15092 16346
rect 14846 16292 14852 16294
rect 14908 16292 14932 16294
rect 14988 16292 15012 16294
rect 15068 16292 15092 16294
rect 15148 16292 15154 16294
rect 14846 16283 15154 16292
rect 21794 16348 22102 16357
rect 21794 16346 21800 16348
rect 21856 16346 21880 16348
rect 21936 16346 21960 16348
rect 22016 16346 22040 16348
rect 22096 16346 22102 16348
rect 21856 16294 21858 16346
rect 22038 16294 22040 16346
rect 21794 16292 21800 16294
rect 21856 16292 21880 16294
rect 21936 16292 21960 16294
rect 22016 16292 22040 16294
rect 22096 16292 22102 16294
rect 21794 16283 22102 16292
rect 4424 15804 4732 15813
rect 4424 15802 4430 15804
rect 4486 15802 4510 15804
rect 4566 15802 4590 15804
rect 4646 15802 4670 15804
rect 4726 15802 4732 15804
rect 4486 15750 4488 15802
rect 4668 15750 4670 15802
rect 4424 15748 4430 15750
rect 4486 15748 4510 15750
rect 4566 15748 4590 15750
rect 4646 15748 4670 15750
rect 4726 15748 4732 15750
rect 4424 15739 4732 15748
rect 11372 15804 11680 15813
rect 11372 15802 11378 15804
rect 11434 15802 11458 15804
rect 11514 15802 11538 15804
rect 11594 15802 11618 15804
rect 11674 15802 11680 15804
rect 11434 15750 11436 15802
rect 11616 15750 11618 15802
rect 11372 15748 11378 15750
rect 11434 15748 11458 15750
rect 11514 15748 11538 15750
rect 11594 15748 11618 15750
rect 11674 15748 11680 15750
rect 11372 15739 11680 15748
rect 18320 15804 18628 15813
rect 18320 15802 18326 15804
rect 18382 15802 18406 15804
rect 18462 15802 18486 15804
rect 18542 15802 18566 15804
rect 18622 15802 18628 15804
rect 18382 15750 18384 15802
rect 18564 15750 18566 15802
rect 18320 15748 18326 15750
rect 18382 15748 18406 15750
rect 18462 15748 18486 15750
rect 18542 15748 18566 15750
rect 18622 15748 18628 15750
rect 18320 15739 18628 15748
rect 25268 15804 25576 15813
rect 25268 15802 25274 15804
rect 25330 15802 25354 15804
rect 25410 15802 25434 15804
rect 25490 15802 25514 15804
rect 25570 15802 25576 15804
rect 25330 15750 25332 15802
rect 25512 15750 25514 15802
rect 25268 15748 25274 15750
rect 25330 15748 25354 15750
rect 25410 15748 25434 15750
rect 25490 15748 25514 15750
rect 25570 15748 25576 15750
rect 25268 15739 25576 15748
rect 7898 15260 8206 15269
rect 7898 15258 7904 15260
rect 7960 15258 7984 15260
rect 8040 15258 8064 15260
rect 8120 15258 8144 15260
rect 8200 15258 8206 15260
rect 7960 15206 7962 15258
rect 8142 15206 8144 15258
rect 7898 15204 7904 15206
rect 7960 15204 7984 15206
rect 8040 15204 8064 15206
rect 8120 15204 8144 15206
rect 8200 15204 8206 15206
rect 7898 15195 8206 15204
rect 14846 15260 15154 15269
rect 14846 15258 14852 15260
rect 14908 15258 14932 15260
rect 14988 15258 15012 15260
rect 15068 15258 15092 15260
rect 15148 15258 15154 15260
rect 14908 15206 14910 15258
rect 15090 15206 15092 15258
rect 14846 15204 14852 15206
rect 14908 15204 14932 15206
rect 14988 15204 15012 15206
rect 15068 15204 15092 15206
rect 15148 15204 15154 15206
rect 14846 15195 15154 15204
rect 21794 15260 22102 15269
rect 21794 15258 21800 15260
rect 21856 15258 21880 15260
rect 21936 15258 21960 15260
rect 22016 15258 22040 15260
rect 22096 15258 22102 15260
rect 21856 15206 21858 15258
rect 22038 15206 22040 15258
rect 21794 15204 21800 15206
rect 21856 15204 21880 15206
rect 21936 15204 21960 15206
rect 22016 15204 22040 15206
rect 22096 15204 22102 15206
rect 21794 15195 22102 15204
rect 4424 14716 4732 14725
rect 4424 14714 4430 14716
rect 4486 14714 4510 14716
rect 4566 14714 4590 14716
rect 4646 14714 4670 14716
rect 4726 14714 4732 14716
rect 4486 14662 4488 14714
rect 4668 14662 4670 14714
rect 4424 14660 4430 14662
rect 4486 14660 4510 14662
rect 4566 14660 4590 14662
rect 4646 14660 4670 14662
rect 4726 14660 4732 14662
rect 4424 14651 4732 14660
rect 11372 14716 11680 14725
rect 11372 14714 11378 14716
rect 11434 14714 11458 14716
rect 11514 14714 11538 14716
rect 11594 14714 11618 14716
rect 11674 14714 11680 14716
rect 11434 14662 11436 14714
rect 11616 14662 11618 14714
rect 11372 14660 11378 14662
rect 11434 14660 11458 14662
rect 11514 14660 11538 14662
rect 11594 14660 11618 14662
rect 11674 14660 11680 14662
rect 11372 14651 11680 14660
rect 18320 14716 18628 14725
rect 18320 14714 18326 14716
rect 18382 14714 18406 14716
rect 18462 14714 18486 14716
rect 18542 14714 18566 14716
rect 18622 14714 18628 14716
rect 18382 14662 18384 14714
rect 18564 14662 18566 14714
rect 18320 14660 18326 14662
rect 18382 14660 18406 14662
rect 18462 14660 18486 14662
rect 18542 14660 18566 14662
rect 18622 14660 18628 14662
rect 18320 14651 18628 14660
rect 25268 14716 25576 14725
rect 25268 14714 25274 14716
rect 25330 14714 25354 14716
rect 25410 14714 25434 14716
rect 25490 14714 25514 14716
rect 25570 14714 25576 14716
rect 25330 14662 25332 14714
rect 25512 14662 25514 14714
rect 25268 14660 25274 14662
rect 25330 14660 25354 14662
rect 25410 14660 25434 14662
rect 25490 14660 25514 14662
rect 25570 14660 25576 14662
rect 25268 14651 25576 14660
rect 7898 14172 8206 14181
rect 7898 14170 7904 14172
rect 7960 14170 7984 14172
rect 8040 14170 8064 14172
rect 8120 14170 8144 14172
rect 8200 14170 8206 14172
rect 7960 14118 7962 14170
rect 8142 14118 8144 14170
rect 7898 14116 7904 14118
rect 7960 14116 7984 14118
rect 8040 14116 8064 14118
rect 8120 14116 8144 14118
rect 8200 14116 8206 14118
rect 7898 14107 8206 14116
rect 14846 14172 15154 14181
rect 14846 14170 14852 14172
rect 14908 14170 14932 14172
rect 14988 14170 15012 14172
rect 15068 14170 15092 14172
rect 15148 14170 15154 14172
rect 14908 14118 14910 14170
rect 15090 14118 15092 14170
rect 14846 14116 14852 14118
rect 14908 14116 14932 14118
rect 14988 14116 15012 14118
rect 15068 14116 15092 14118
rect 15148 14116 15154 14118
rect 14846 14107 15154 14116
rect 21794 14172 22102 14181
rect 21794 14170 21800 14172
rect 21856 14170 21880 14172
rect 21936 14170 21960 14172
rect 22016 14170 22040 14172
rect 22096 14170 22102 14172
rect 21856 14118 21858 14170
rect 22038 14118 22040 14170
rect 21794 14116 21800 14118
rect 21856 14116 21880 14118
rect 21936 14116 21960 14118
rect 22016 14116 22040 14118
rect 22096 14116 22102 14118
rect 21794 14107 22102 14116
rect 28172 13864 28224 13870
rect 28172 13806 28224 13812
rect 28184 13705 28212 13806
rect 28170 13696 28226 13705
rect 4424 13628 4732 13637
rect 4424 13626 4430 13628
rect 4486 13626 4510 13628
rect 4566 13626 4590 13628
rect 4646 13626 4670 13628
rect 4726 13626 4732 13628
rect 4486 13574 4488 13626
rect 4668 13574 4670 13626
rect 4424 13572 4430 13574
rect 4486 13572 4510 13574
rect 4566 13572 4590 13574
rect 4646 13572 4670 13574
rect 4726 13572 4732 13574
rect 4424 13563 4732 13572
rect 11372 13628 11680 13637
rect 11372 13626 11378 13628
rect 11434 13626 11458 13628
rect 11514 13626 11538 13628
rect 11594 13626 11618 13628
rect 11674 13626 11680 13628
rect 11434 13574 11436 13626
rect 11616 13574 11618 13626
rect 11372 13572 11378 13574
rect 11434 13572 11458 13574
rect 11514 13572 11538 13574
rect 11594 13572 11618 13574
rect 11674 13572 11680 13574
rect 11372 13563 11680 13572
rect 18320 13628 18628 13637
rect 18320 13626 18326 13628
rect 18382 13626 18406 13628
rect 18462 13626 18486 13628
rect 18542 13626 18566 13628
rect 18622 13626 18628 13628
rect 18382 13574 18384 13626
rect 18564 13574 18566 13626
rect 18320 13572 18326 13574
rect 18382 13572 18406 13574
rect 18462 13572 18486 13574
rect 18542 13572 18566 13574
rect 18622 13572 18628 13574
rect 18320 13563 18628 13572
rect 25268 13628 25576 13637
rect 28170 13631 28226 13640
rect 25268 13626 25274 13628
rect 25330 13626 25354 13628
rect 25410 13626 25434 13628
rect 25490 13626 25514 13628
rect 25570 13626 25576 13628
rect 25330 13574 25332 13626
rect 25512 13574 25514 13626
rect 25268 13572 25274 13574
rect 25330 13572 25354 13574
rect 25410 13572 25434 13574
rect 25490 13572 25514 13574
rect 25570 13572 25576 13574
rect 25268 13563 25576 13572
rect 7898 13084 8206 13093
rect 7898 13082 7904 13084
rect 7960 13082 7984 13084
rect 8040 13082 8064 13084
rect 8120 13082 8144 13084
rect 8200 13082 8206 13084
rect 7960 13030 7962 13082
rect 8142 13030 8144 13082
rect 7898 13028 7904 13030
rect 7960 13028 7984 13030
rect 8040 13028 8064 13030
rect 8120 13028 8144 13030
rect 8200 13028 8206 13030
rect 7898 13019 8206 13028
rect 14846 13084 15154 13093
rect 14846 13082 14852 13084
rect 14908 13082 14932 13084
rect 14988 13082 15012 13084
rect 15068 13082 15092 13084
rect 15148 13082 15154 13084
rect 14908 13030 14910 13082
rect 15090 13030 15092 13082
rect 14846 13028 14852 13030
rect 14908 13028 14932 13030
rect 14988 13028 15012 13030
rect 15068 13028 15092 13030
rect 15148 13028 15154 13030
rect 14846 13019 15154 13028
rect 21794 13084 22102 13093
rect 21794 13082 21800 13084
rect 21856 13082 21880 13084
rect 21936 13082 21960 13084
rect 22016 13082 22040 13084
rect 22096 13082 22102 13084
rect 21856 13030 21858 13082
rect 22038 13030 22040 13082
rect 21794 13028 21800 13030
rect 21856 13028 21880 13030
rect 21936 13028 21960 13030
rect 22016 13028 22040 13030
rect 22096 13028 22102 13030
rect 21794 13019 22102 13028
rect 4424 12540 4732 12549
rect 4424 12538 4430 12540
rect 4486 12538 4510 12540
rect 4566 12538 4590 12540
rect 4646 12538 4670 12540
rect 4726 12538 4732 12540
rect 4486 12486 4488 12538
rect 4668 12486 4670 12538
rect 4424 12484 4430 12486
rect 4486 12484 4510 12486
rect 4566 12484 4590 12486
rect 4646 12484 4670 12486
rect 4726 12484 4732 12486
rect 4424 12475 4732 12484
rect 11372 12540 11680 12549
rect 11372 12538 11378 12540
rect 11434 12538 11458 12540
rect 11514 12538 11538 12540
rect 11594 12538 11618 12540
rect 11674 12538 11680 12540
rect 11434 12486 11436 12538
rect 11616 12486 11618 12538
rect 11372 12484 11378 12486
rect 11434 12484 11458 12486
rect 11514 12484 11538 12486
rect 11594 12484 11618 12486
rect 11674 12484 11680 12486
rect 11372 12475 11680 12484
rect 18320 12540 18628 12549
rect 18320 12538 18326 12540
rect 18382 12538 18406 12540
rect 18462 12538 18486 12540
rect 18542 12538 18566 12540
rect 18622 12538 18628 12540
rect 18382 12486 18384 12538
rect 18564 12486 18566 12538
rect 18320 12484 18326 12486
rect 18382 12484 18406 12486
rect 18462 12484 18486 12486
rect 18542 12484 18566 12486
rect 18622 12484 18628 12486
rect 18320 12475 18628 12484
rect 25268 12540 25576 12549
rect 25268 12538 25274 12540
rect 25330 12538 25354 12540
rect 25410 12538 25434 12540
rect 25490 12538 25514 12540
rect 25570 12538 25576 12540
rect 25330 12486 25332 12538
rect 25512 12486 25514 12538
rect 25268 12484 25274 12486
rect 25330 12484 25354 12486
rect 25410 12484 25434 12486
rect 25490 12484 25514 12486
rect 25570 12484 25576 12486
rect 25268 12475 25576 12484
rect 7898 11996 8206 12005
rect 7898 11994 7904 11996
rect 7960 11994 7984 11996
rect 8040 11994 8064 11996
rect 8120 11994 8144 11996
rect 8200 11994 8206 11996
rect 7960 11942 7962 11994
rect 8142 11942 8144 11994
rect 7898 11940 7904 11942
rect 7960 11940 7984 11942
rect 8040 11940 8064 11942
rect 8120 11940 8144 11942
rect 8200 11940 8206 11942
rect 7898 11931 8206 11940
rect 14846 11996 15154 12005
rect 14846 11994 14852 11996
rect 14908 11994 14932 11996
rect 14988 11994 15012 11996
rect 15068 11994 15092 11996
rect 15148 11994 15154 11996
rect 14908 11942 14910 11994
rect 15090 11942 15092 11994
rect 14846 11940 14852 11942
rect 14908 11940 14932 11942
rect 14988 11940 15012 11942
rect 15068 11940 15092 11942
rect 15148 11940 15154 11942
rect 14846 11931 15154 11940
rect 21794 11996 22102 12005
rect 21794 11994 21800 11996
rect 21856 11994 21880 11996
rect 21936 11994 21960 11996
rect 22016 11994 22040 11996
rect 22096 11994 22102 11996
rect 21856 11942 21858 11994
rect 22038 11942 22040 11994
rect 21794 11940 21800 11942
rect 21856 11940 21880 11942
rect 21936 11940 21960 11942
rect 22016 11940 22040 11942
rect 22096 11940 22102 11942
rect 21794 11931 22102 11940
rect 4424 11452 4732 11461
rect 4424 11450 4430 11452
rect 4486 11450 4510 11452
rect 4566 11450 4590 11452
rect 4646 11450 4670 11452
rect 4726 11450 4732 11452
rect 4486 11398 4488 11450
rect 4668 11398 4670 11450
rect 4424 11396 4430 11398
rect 4486 11396 4510 11398
rect 4566 11396 4590 11398
rect 4646 11396 4670 11398
rect 4726 11396 4732 11398
rect 4424 11387 4732 11396
rect 11372 11452 11680 11461
rect 11372 11450 11378 11452
rect 11434 11450 11458 11452
rect 11514 11450 11538 11452
rect 11594 11450 11618 11452
rect 11674 11450 11680 11452
rect 11434 11398 11436 11450
rect 11616 11398 11618 11450
rect 11372 11396 11378 11398
rect 11434 11396 11458 11398
rect 11514 11396 11538 11398
rect 11594 11396 11618 11398
rect 11674 11396 11680 11398
rect 11372 11387 11680 11396
rect 18320 11452 18628 11461
rect 18320 11450 18326 11452
rect 18382 11450 18406 11452
rect 18462 11450 18486 11452
rect 18542 11450 18566 11452
rect 18622 11450 18628 11452
rect 18382 11398 18384 11450
rect 18564 11398 18566 11450
rect 18320 11396 18326 11398
rect 18382 11396 18406 11398
rect 18462 11396 18486 11398
rect 18542 11396 18566 11398
rect 18622 11396 18628 11398
rect 18320 11387 18628 11396
rect 25268 11452 25576 11461
rect 25268 11450 25274 11452
rect 25330 11450 25354 11452
rect 25410 11450 25434 11452
rect 25490 11450 25514 11452
rect 25570 11450 25576 11452
rect 25330 11398 25332 11450
rect 25512 11398 25514 11450
rect 25268 11396 25274 11398
rect 25330 11396 25354 11398
rect 25410 11396 25434 11398
rect 25490 11396 25514 11398
rect 25570 11396 25576 11398
rect 25268 11387 25576 11396
rect 7898 10908 8206 10917
rect 7898 10906 7904 10908
rect 7960 10906 7984 10908
rect 8040 10906 8064 10908
rect 8120 10906 8144 10908
rect 8200 10906 8206 10908
rect 7960 10854 7962 10906
rect 8142 10854 8144 10906
rect 7898 10852 7904 10854
rect 7960 10852 7984 10854
rect 8040 10852 8064 10854
rect 8120 10852 8144 10854
rect 8200 10852 8206 10854
rect 7898 10843 8206 10852
rect 14846 10908 15154 10917
rect 14846 10906 14852 10908
rect 14908 10906 14932 10908
rect 14988 10906 15012 10908
rect 15068 10906 15092 10908
rect 15148 10906 15154 10908
rect 14908 10854 14910 10906
rect 15090 10854 15092 10906
rect 14846 10852 14852 10854
rect 14908 10852 14932 10854
rect 14988 10852 15012 10854
rect 15068 10852 15092 10854
rect 15148 10852 15154 10854
rect 14846 10843 15154 10852
rect 21794 10908 22102 10917
rect 21794 10906 21800 10908
rect 21856 10906 21880 10908
rect 21936 10906 21960 10908
rect 22016 10906 22040 10908
rect 22096 10906 22102 10908
rect 21856 10854 21858 10906
rect 22038 10854 22040 10906
rect 21794 10852 21800 10854
rect 21856 10852 21880 10854
rect 21936 10852 21960 10854
rect 22016 10852 22040 10854
rect 22096 10852 22102 10854
rect 21794 10843 22102 10852
rect 4424 10364 4732 10373
rect 4424 10362 4430 10364
rect 4486 10362 4510 10364
rect 4566 10362 4590 10364
rect 4646 10362 4670 10364
rect 4726 10362 4732 10364
rect 4486 10310 4488 10362
rect 4668 10310 4670 10362
rect 4424 10308 4430 10310
rect 4486 10308 4510 10310
rect 4566 10308 4590 10310
rect 4646 10308 4670 10310
rect 4726 10308 4732 10310
rect 4424 10299 4732 10308
rect 11372 10364 11680 10373
rect 11372 10362 11378 10364
rect 11434 10362 11458 10364
rect 11514 10362 11538 10364
rect 11594 10362 11618 10364
rect 11674 10362 11680 10364
rect 11434 10310 11436 10362
rect 11616 10310 11618 10362
rect 11372 10308 11378 10310
rect 11434 10308 11458 10310
rect 11514 10308 11538 10310
rect 11594 10308 11618 10310
rect 11674 10308 11680 10310
rect 11372 10299 11680 10308
rect 18320 10364 18628 10373
rect 18320 10362 18326 10364
rect 18382 10362 18406 10364
rect 18462 10362 18486 10364
rect 18542 10362 18566 10364
rect 18622 10362 18628 10364
rect 18382 10310 18384 10362
rect 18564 10310 18566 10362
rect 18320 10308 18326 10310
rect 18382 10308 18406 10310
rect 18462 10308 18486 10310
rect 18542 10308 18566 10310
rect 18622 10308 18628 10310
rect 18320 10299 18628 10308
rect 25268 10364 25576 10373
rect 25268 10362 25274 10364
rect 25330 10362 25354 10364
rect 25410 10362 25434 10364
rect 25490 10362 25514 10364
rect 25570 10362 25576 10364
rect 25330 10310 25332 10362
rect 25512 10310 25514 10362
rect 25268 10308 25274 10310
rect 25330 10308 25354 10310
rect 25410 10308 25434 10310
rect 25490 10308 25514 10310
rect 25570 10308 25576 10310
rect 25268 10299 25576 10308
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 7898 9820 8206 9829
rect 7898 9818 7904 9820
rect 7960 9818 7984 9820
rect 8040 9818 8064 9820
rect 8120 9818 8144 9820
rect 8200 9818 8206 9820
rect 7960 9766 7962 9818
rect 8142 9766 8144 9818
rect 7898 9764 7904 9766
rect 7960 9764 7984 9766
rect 8040 9764 8064 9766
rect 8120 9764 8144 9766
rect 8200 9764 8206 9766
rect 7898 9755 8206 9764
rect 4424 9276 4732 9285
rect 4424 9274 4430 9276
rect 4486 9274 4510 9276
rect 4566 9274 4590 9276
rect 4646 9274 4670 9276
rect 4726 9274 4732 9276
rect 4486 9222 4488 9274
rect 4668 9222 4670 9274
rect 4424 9220 4430 9222
rect 4486 9220 4510 9222
rect 4566 9220 4590 9222
rect 4646 9220 4670 9222
rect 4726 9220 4732 9222
rect 4424 9211 4732 9220
rect 11372 9276 11680 9285
rect 11372 9274 11378 9276
rect 11434 9274 11458 9276
rect 11514 9274 11538 9276
rect 11594 9274 11618 9276
rect 11674 9274 11680 9276
rect 11434 9222 11436 9274
rect 11616 9222 11618 9274
rect 11372 9220 11378 9222
rect 11434 9220 11458 9222
rect 11514 9220 11538 9222
rect 11594 9220 11618 9222
rect 11674 9220 11680 9222
rect 11372 9211 11680 9220
rect 7898 8732 8206 8741
rect 7898 8730 7904 8732
rect 7960 8730 7984 8732
rect 8040 8730 8064 8732
rect 8120 8730 8144 8732
rect 8200 8730 8206 8732
rect 7960 8678 7962 8730
rect 8142 8678 8144 8730
rect 7898 8676 7904 8678
rect 7960 8676 7984 8678
rect 8040 8676 8064 8678
rect 8120 8676 8144 8678
rect 8200 8676 8206 8678
rect 7898 8667 8206 8676
rect 4424 8188 4732 8197
rect 4424 8186 4430 8188
rect 4486 8186 4510 8188
rect 4566 8186 4590 8188
rect 4646 8186 4670 8188
rect 4726 8186 4732 8188
rect 4486 8134 4488 8186
rect 4668 8134 4670 8186
rect 4424 8132 4430 8134
rect 4486 8132 4510 8134
rect 4566 8132 4590 8134
rect 4646 8132 4670 8134
rect 4726 8132 4732 8134
rect 4424 8123 4732 8132
rect 11372 8188 11680 8197
rect 11372 8186 11378 8188
rect 11434 8186 11458 8188
rect 11514 8186 11538 8188
rect 11594 8186 11618 8188
rect 11674 8186 11680 8188
rect 11434 8134 11436 8186
rect 11616 8134 11618 8186
rect 11372 8132 11378 8134
rect 11434 8132 11458 8134
rect 11514 8132 11538 8134
rect 11594 8132 11618 8134
rect 11674 8132 11680 8134
rect 11372 8123 11680 8132
rect 7898 7644 8206 7653
rect 7898 7642 7904 7644
rect 7960 7642 7984 7644
rect 8040 7642 8064 7644
rect 8120 7642 8144 7644
rect 8200 7642 8206 7644
rect 7960 7590 7962 7642
rect 8142 7590 8144 7642
rect 7898 7588 7904 7590
rect 7960 7588 7984 7590
rect 8040 7588 8064 7590
rect 8120 7588 8144 7590
rect 8200 7588 8206 7590
rect 7898 7579 8206 7588
rect 14752 7410 14780 9862
rect 14846 9820 15154 9829
rect 14846 9818 14852 9820
rect 14908 9818 14932 9820
rect 14988 9818 15012 9820
rect 15068 9818 15092 9820
rect 15148 9818 15154 9820
rect 14908 9766 14910 9818
rect 15090 9766 15092 9818
rect 14846 9764 14852 9766
rect 14908 9764 14932 9766
rect 14988 9764 15012 9766
rect 15068 9764 15092 9766
rect 15148 9764 15154 9766
rect 14846 9755 15154 9764
rect 21794 9820 22102 9829
rect 21794 9818 21800 9820
rect 21856 9818 21880 9820
rect 21936 9818 21960 9820
rect 22016 9818 22040 9820
rect 22096 9818 22102 9820
rect 21856 9766 21858 9818
rect 22038 9766 22040 9818
rect 21794 9764 21800 9766
rect 21856 9764 21880 9766
rect 21936 9764 21960 9766
rect 22016 9764 22040 9766
rect 22096 9764 22102 9766
rect 21794 9755 22102 9764
rect 27540 9625 27568 9998
rect 27526 9616 27582 9625
rect 27526 9551 27582 9560
rect 18320 9276 18628 9285
rect 18320 9274 18326 9276
rect 18382 9274 18406 9276
rect 18462 9274 18486 9276
rect 18542 9274 18566 9276
rect 18622 9274 18628 9276
rect 18382 9222 18384 9274
rect 18564 9222 18566 9274
rect 18320 9220 18326 9222
rect 18382 9220 18406 9222
rect 18462 9220 18486 9222
rect 18542 9220 18566 9222
rect 18622 9220 18628 9222
rect 18320 9211 18628 9220
rect 25268 9276 25576 9285
rect 25268 9274 25274 9276
rect 25330 9274 25354 9276
rect 25410 9274 25434 9276
rect 25490 9274 25514 9276
rect 25570 9274 25576 9276
rect 25330 9222 25332 9274
rect 25512 9222 25514 9274
rect 25268 9220 25274 9222
rect 25330 9220 25354 9222
rect 25410 9220 25434 9222
rect 25490 9220 25514 9222
rect 25570 9220 25576 9222
rect 25268 9211 25576 9220
rect 14846 8732 15154 8741
rect 14846 8730 14852 8732
rect 14908 8730 14932 8732
rect 14988 8730 15012 8732
rect 15068 8730 15092 8732
rect 15148 8730 15154 8732
rect 14908 8678 14910 8730
rect 15090 8678 15092 8730
rect 14846 8676 14852 8678
rect 14908 8676 14932 8678
rect 14988 8676 15012 8678
rect 15068 8676 15092 8678
rect 15148 8676 15154 8678
rect 14846 8667 15154 8676
rect 21794 8732 22102 8741
rect 21794 8730 21800 8732
rect 21856 8730 21880 8732
rect 21936 8730 21960 8732
rect 22016 8730 22040 8732
rect 22096 8730 22102 8732
rect 21856 8678 21858 8730
rect 22038 8678 22040 8730
rect 21794 8676 21800 8678
rect 21856 8676 21880 8678
rect 21936 8676 21960 8678
rect 22016 8676 22040 8678
rect 22096 8676 22102 8678
rect 21794 8667 22102 8676
rect 18320 8188 18628 8197
rect 18320 8186 18326 8188
rect 18382 8186 18406 8188
rect 18462 8186 18486 8188
rect 18542 8186 18566 8188
rect 18622 8186 18628 8188
rect 18382 8134 18384 8186
rect 18564 8134 18566 8186
rect 18320 8132 18326 8134
rect 18382 8132 18406 8134
rect 18462 8132 18486 8134
rect 18542 8132 18566 8134
rect 18622 8132 18628 8134
rect 18320 8123 18628 8132
rect 25268 8188 25576 8197
rect 25268 8186 25274 8188
rect 25330 8186 25354 8188
rect 25410 8186 25434 8188
rect 25490 8186 25514 8188
rect 25570 8186 25576 8188
rect 25330 8134 25332 8186
rect 25512 8134 25514 8186
rect 25268 8132 25274 8134
rect 25330 8132 25354 8134
rect 25410 8132 25434 8134
rect 25490 8132 25514 8134
rect 25570 8132 25576 8134
rect 25268 8123 25576 8132
rect 14846 7644 15154 7653
rect 14846 7642 14852 7644
rect 14908 7642 14932 7644
rect 14988 7642 15012 7644
rect 15068 7642 15092 7644
rect 15148 7642 15154 7644
rect 14908 7590 14910 7642
rect 15090 7590 15092 7642
rect 14846 7588 14852 7590
rect 14908 7588 14932 7590
rect 14988 7588 15012 7590
rect 15068 7588 15092 7590
rect 15148 7588 15154 7590
rect 14846 7579 15154 7588
rect 21794 7644 22102 7653
rect 21794 7642 21800 7644
rect 21856 7642 21880 7644
rect 21936 7642 21960 7644
rect 22016 7642 22040 7644
rect 22096 7642 22102 7644
rect 21856 7590 21858 7642
rect 22038 7590 22040 7642
rect 21794 7588 21800 7590
rect 21856 7588 21880 7590
rect 21936 7588 21960 7590
rect 22016 7588 22040 7590
rect 22096 7588 22102 7590
rect 21794 7579 22102 7588
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 4424 7100 4732 7109
rect 4424 7098 4430 7100
rect 4486 7098 4510 7100
rect 4566 7098 4590 7100
rect 4646 7098 4670 7100
rect 4726 7098 4732 7100
rect 4486 7046 4488 7098
rect 4668 7046 4670 7098
rect 4424 7044 4430 7046
rect 4486 7044 4510 7046
rect 4566 7044 4590 7046
rect 4646 7044 4670 7046
rect 4726 7044 4732 7046
rect 4424 7035 4732 7044
rect 4424 6012 4732 6021
rect 4424 6010 4430 6012
rect 4486 6010 4510 6012
rect 4566 6010 4590 6012
rect 4646 6010 4670 6012
rect 4726 6010 4732 6012
rect 4486 5958 4488 6010
rect 4668 5958 4670 6010
rect 4424 5956 4430 5958
rect 4486 5956 4510 5958
rect 4566 5956 4590 5958
rect 4646 5956 4670 5958
rect 4726 5956 4732 5958
rect 4424 5947 4732 5956
rect 4424 4924 4732 4933
rect 4424 4922 4430 4924
rect 4486 4922 4510 4924
rect 4566 4922 4590 4924
rect 4646 4922 4670 4924
rect 4726 4922 4732 4924
rect 4486 4870 4488 4922
rect 4668 4870 4670 4922
rect 4424 4868 4430 4870
rect 4486 4868 4510 4870
rect 4566 4868 4590 4870
rect 4646 4868 4670 4870
rect 4726 4868 4732 4870
rect 4424 4859 4732 4868
rect 4424 3836 4732 3845
rect 4424 3834 4430 3836
rect 4486 3834 4510 3836
rect 4566 3834 4590 3836
rect 4646 3834 4670 3836
rect 4726 3834 4732 3836
rect 4486 3782 4488 3834
rect 4668 3782 4670 3834
rect 4424 3780 4430 3782
rect 4486 3780 4510 3782
rect 4566 3780 4590 3782
rect 4646 3780 4670 3782
rect 4726 3780 4732 3782
rect 4424 3771 4732 3780
rect 4424 2748 4732 2757
rect 4424 2746 4430 2748
rect 4486 2746 4510 2748
rect 4566 2746 4590 2748
rect 4646 2746 4670 2748
rect 4726 2746 4732 2748
rect 4486 2694 4488 2746
rect 4668 2694 4670 2746
rect 4424 2692 4430 2694
rect 4486 2692 4510 2694
rect 4566 2692 4590 2694
rect 4646 2692 4670 2694
rect 4726 2692 4732 2694
rect 4424 2683 4732 2692
rect 7484 2446 7512 7142
rect 11372 7100 11680 7109
rect 11372 7098 11378 7100
rect 11434 7098 11458 7100
rect 11514 7098 11538 7100
rect 11594 7098 11618 7100
rect 11674 7098 11680 7100
rect 11434 7046 11436 7098
rect 11616 7046 11618 7098
rect 11372 7044 11378 7046
rect 11434 7044 11458 7046
rect 11514 7044 11538 7046
rect 11594 7044 11618 7046
rect 11674 7044 11680 7046
rect 11372 7035 11680 7044
rect 18320 7100 18628 7109
rect 18320 7098 18326 7100
rect 18382 7098 18406 7100
rect 18462 7098 18486 7100
rect 18542 7098 18566 7100
rect 18622 7098 18628 7100
rect 18382 7046 18384 7098
rect 18564 7046 18566 7098
rect 18320 7044 18326 7046
rect 18382 7044 18406 7046
rect 18462 7044 18486 7046
rect 18542 7044 18566 7046
rect 18622 7044 18628 7046
rect 18320 7035 18628 7044
rect 25268 7100 25576 7109
rect 25268 7098 25274 7100
rect 25330 7098 25354 7100
rect 25410 7098 25434 7100
rect 25490 7098 25514 7100
rect 25570 7098 25576 7100
rect 25330 7046 25332 7098
rect 25512 7046 25514 7098
rect 25268 7044 25274 7046
rect 25330 7044 25354 7046
rect 25410 7044 25434 7046
rect 25490 7044 25514 7046
rect 25570 7044 25576 7046
rect 25268 7035 25576 7044
rect 7898 6556 8206 6565
rect 7898 6554 7904 6556
rect 7960 6554 7984 6556
rect 8040 6554 8064 6556
rect 8120 6554 8144 6556
rect 8200 6554 8206 6556
rect 7960 6502 7962 6554
rect 8142 6502 8144 6554
rect 7898 6500 7904 6502
rect 7960 6500 7984 6502
rect 8040 6500 8064 6502
rect 8120 6500 8144 6502
rect 8200 6500 8206 6502
rect 7898 6491 8206 6500
rect 14846 6556 15154 6565
rect 14846 6554 14852 6556
rect 14908 6554 14932 6556
rect 14988 6554 15012 6556
rect 15068 6554 15092 6556
rect 15148 6554 15154 6556
rect 14908 6502 14910 6554
rect 15090 6502 15092 6554
rect 14846 6500 14852 6502
rect 14908 6500 14932 6502
rect 14988 6500 15012 6502
rect 15068 6500 15092 6502
rect 15148 6500 15154 6502
rect 14846 6491 15154 6500
rect 21794 6556 22102 6565
rect 21794 6554 21800 6556
rect 21856 6554 21880 6556
rect 21936 6554 21960 6556
rect 22016 6554 22040 6556
rect 22096 6554 22102 6556
rect 21856 6502 21858 6554
rect 22038 6502 22040 6554
rect 21794 6500 21800 6502
rect 21856 6500 21880 6502
rect 21936 6500 21960 6502
rect 22016 6500 22040 6502
rect 22096 6500 22102 6502
rect 21794 6491 22102 6500
rect 11372 6012 11680 6021
rect 11372 6010 11378 6012
rect 11434 6010 11458 6012
rect 11514 6010 11538 6012
rect 11594 6010 11618 6012
rect 11674 6010 11680 6012
rect 11434 5958 11436 6010
rect 11616 5958 11618 6010
rect 11372 5956 11378 5958
rect 11434 5956 11458 5958
rect 11514 5956 11538 5958
rect 11594 5956 11618 5958
rect 11674 5956 11680 5958
rect 11372 5947 11680 5956
rect 18320 6012 18628 6021
rect 18320 6010 18326 6012
rect 18382 6010 18406 6012
rect 18462 6010 18486 6012
rect 18542 6010 18566 6012
rect 18622 6010 18628 6012
rect 18382 5958 18384 6010
rect 18564 5958 18566 6010
rect 18320 5956 18326 5958
rect 18382 5956 18406 5958
rect 18462 5956 18486 5958
rect 18542 5956 18566 5958
rect 18622 5956 18628 5958
rect 18320 5947 18628 5956
rect 25268 6012 25576 6021
rect 25268 6010 25274 6012
rect 25330 6010 25354 6012
rect 25410 6010 25434 6012
rect 25490 6010 25514 6012
rect 25570 6010 25576 6012
rect 25330 5958 25332 6010
rect 25512 5958 25514 6010
rect 25268 5956 25274 5958
rect 25330 5956 25354 5958
rect 25410 5956 25434 5958
rect 25490 5956 25514 5958
rect 25570 5956 25576 5958
rect 25268 5947 25576 5956
rect 7898 5468 8206 5477
rect 7898 5466 7904 5468
rect 7960 5466 7984 5468
rect 8040 5466 8064 5468
rect 8120 5466 8144 5468
rect 8200 5466 8206 5468
rect 7960 5414 7962 5466
rect 8142 5414 8144 5466
rect 7898 5412 7904 5414
rect 7960 5412 7984 5414
rect 8040 5412 8064 5414
rect 8120 5412 8144 5414
rect 8200 5412 8206 5414
rect 7898 5403 8206 5412
rect 14846 5468 15154 5477
rect 14846 5466 14852 5468
rect 14908 5466 14932 5468
rect 14988 5466 15012 5468
rect 15068 5466 15092 5468
rect 15148 5466 15154 5468
rect 14908 5414 14910 5466
rect 15090 5414 15092 5466
rect 14846 5412 14852 5414
rect 14908 5412 14932 5414
rect 14988 5412 15012 5414
rect 15068 5412 15092 5414
rect 15148 5412 15154 5414
rect 14846 5403 15154 5412
rect 21794 5468 22102 5477
rect 21794 5466 21800 5468
rect 21856 5466 21880 5468
rect 21936 5466 21960 5468
rect 22016 5466 22040 5468
rect 22096 5466 22102 5468
rect 21856 5414 21858 5466
rect 22038 5414 22040 5466
rect 21794 5412 21800 5414
rect 21856 5412 21880 5414
rect 21936 5412 21960 5414
rect 22016 5412 22040 5414
rect 22096 5412 22102 5414
rect 21794 5403 22102 5412
rect 11372 4924 11680 4933
rect 11372 4922 11378 4924
rect 11434 4922 11458 4924
rect 11514 4922 11538 4924
rect 11594 4922 11618 4924
rect 11674 4922 11680 4924
rect 11434 4870 11436 4922
rect 11616 4870 11618 4922
rect 11372 4868 11378 4870
rect 11434 4868 11458 4870
rect 11514 4868 11538 4870
rect 11594 4868 11618 4870
rect 11674 4868 11680 4870
rect 11372 4859 11680 4868
rect 18320 4924 18628 4933
rect 18320 4922 18326 4924
rect 18382 4922 18406 4924
rect 18462 4922 18486 4924
rect 18542 4922 18566 4924
rect 18622 4922 18628 4924
rect 18382 4870 18384 4922
rect 18564 4870 18566 4922
rect 18320 4868 18326 4870
rect 18382 4868 18406 4870
rect 18462 4868 18486 4870
rect 18542 4868 18566 4870
rect 18622 4868 18628 4870
rect 18320 4859 18628 4868
rect 25268 4924 25576 4933
rect 25268 4922 25274 4924
rect 25330 4922 25354 4924
rect 25410 4922 25434 4924
rect 25490 4922 25514 4924
rect 25570 4922 25576 4924
rect 25330 4870 25332 4922
rect 25512 4870 25514 4922
rect 25268 4868 25274 4870
rect 25330 4868 25354 4870
rect 25410 4868 25434 4870
rect 25490 4868 25514 4870
rect 25570 4868 25576 4870
rect 25268 4859 25576 4868
rect 7898 4380 8206 4389
rect 7898 4378 7904 4380
rect 7960 4378 7984 4380
rect 8040 4378 8064 4380
rect 8120 4378 8144 4380
rect 8200 4378 8206 4380
rect 7960 4326 7962 4378
rect 8142 4326 8144 4378
rect 7898 4324 7904 4326
rect 7960 4324 7984 4326
rect 8040 4324 8064 4326
rect 8120 4324 8144 4326
rect 8200 4324 8206 4326
rect 7898 4315 8206 4324
rect 14846 4380 15154 4389
rect 14846 4378 14852 4380
rect 14908 4378 14932 4380
rect 14988 4378 15012 4380
rect 15068 4378 15092 4380
rect 15148 4378 15154 4380
rect 14908 4326 14910 4378
rect 15090 4326 15092 4378
rect 14846 4324 14852 4326
rect 14908 4324 14932 4326
rect 14988 4324 15012 4326
rect 15068 4324 15092 4326
rect 15148 4324 15154 4326
rect 14846 4315 15154 4324
rect 21794 4380 22102 4389
rect 21794 4378 21800 4380
rect 21856 4378 21880 4380
rect 21936 4378 21960 4380
rect 22016 4378 22040 4380
rect 22096 4378 22102 4380
rect 21856 4326 21858 4378
rect 22038 4326 22040 4378
rect 21794 4324 21800 4326
rect 21856 4324 21880 4326
rect 21936 4324 21960 4326
rect 22016 4324 22040 4326
rect 22096 4324 22102 4326
rect 21794 4315 22102 4324
rect 11372 3836 11680 3845
rect 11372 3834 11378 3836
rect 11434 3834 11458 3836
rect 11514 3834 11538 3836
rect 11594 3834 11618 3836
rect 11674 3834 11680 3836
rect 11434 3782 11436 3834
rect 11616 3782 11618 3834
rect 11372 3780 11378 3782
rect 11434 3780 11458 3782
rect 11514 3780 11538 3782
rect 11594 3780 11618 3782
rect 11674 3780 11680 3782
rect 11372 3771 11680 3780
rect 18320 3836 18628 3845
rect 18320 3834 18326 3836
rect 18382 3834 18406 3836
rect 18462 3834 18486 3836
rect 18542 3834 18566 3836
rect 18622 3834 18628 3836
rect 18382 3782 18384 3834
rect 18564 3782 18566 3834
rect 18320 3780 18326 3782
rect 18382 3780 18406 3782
rect 18462 3780 18486 3782
rect 18542 3780 18566 3782
rect 18622 3780 18628 3782
rect 18320 3771 18628 3780
rect 25268 3836 25576 3845
rect 25268 3834 25274 3836
rect 25330 3834 25354 3836
rect 25410 3834 25434 3836
rect 25490 3834 25514 3836
rect 25570 3834 25576 3836
rect 25330 3782 25332 3834
rect 25512 3782 25514 3834
rect 25268 3780 25274 3782
rect 25330 3780 25354 3782
rect 25410 3780 25434 3782
rect 25490 3780 25514 3782
rect 25570 3780 25576 3782
rect 25268 3771 25576 3780
rect 7898 3292 8206 3301
rect 7898 3290 7904 3292
rect 7960 3290 7984 3292
rect 8040 3290 8064 3292
rect 8120 3290 8144 3292
rect 8200 3290 8206 3292
rect 7960 3238 7962 3290
rect 8142 3238 8144 3290
rect 7898 3236 7904 3238
rect 7960 3236 7984 3238
rect 8040 3236 8064 3238
rect 8120 3236 8144 3238
rect 8200 3236 8206 3238
rect 7898 3227 8206 3236
rect 14846 3292 15154 3301
rect 14846 3290 14852 3292
rect 14908 3290 14932 3292
rect 14988 3290 15012 3292
rect 15068 3290 15092 3292
rect 15148 3290 15154 3292
rect 14908 3238 14910 3290
rect 15090 3238 15092 3290
rect 14846 3236 14852 3238
rect 14908 3236 14932 3238
rect 14988 3236 15012 3238
rect 15068 3236 15092 3238
rect 15148 3236 15154 3238
rect 14846 3227 15154 3236
rect 21794 3292 22102 3301
rect 21794 3290 21800 3292
rect 21856 3290 21880 3292
rect 21936 3290 21960 3292
rect 22016 3290 22040 3292
rect 22096 3290 22102 3292
rect 21856 3238 21858 3290
rect 22038 3238 22040 3290
rect 21794 3236 21800 3238
rect 21856 3236 21880 3238
rect 21936 3236 21960 3238
rect 22016 3236 22040 3238
rect 22096 3236 22102 3238
rect 21794 3227 22102 3236
rect 11372 2748 11680 2757
rect 11372 2746 11378 2748
rect 11434 2746 11458 2748
rect 11514 2746 11538 2748
rect 11594 2746 11618 2748
rect 11674 2746 11680 2748
rect 11434 2694 11436 2746
rect 11616 2694 11618 2746
rect 11372 2692 11378 2694
rect 11434 2692 11458 2694
rect 11514 2692 11538 2694
rect 11594 2692 11618 2694
rect 11674 2692 11680 2694
rect 11372 2683 11680 2692
rect 18320 2748 18628 2757
rect 18320 2746 18326 2748
rect 18382 2746 18406 2748
rect 18462 2746 18486 2748
rect 18542 2746 18566 2748
rect 18622 2746 18628 2748
rect 18382 2694 18384 2746
rect 18564 2694 18566 2746
rect 18320 2692 18326 2694
rect 18382 2692 18406 2694
rect 18462 2692 18486 2694
rect 18542 2692 18566 2694
rect 18622 2692 18628 2694
rect 18320 2683 18628 2692
rect 25268 2748 25576 2757
rect 25268 2746 25274 2748
rect 25330 2746 25354 2748
rect 25410 2746 25434 2748
rect 25490 2746 25514 2748
rect 25570 2746 25576 2748
rect 25330 2694 25332 2746
rect 25512 2694 25514 2746
rect 25268 2692 25274 2694
rect 25330 2692 25354 2694
rect 25410 2692 25434 2694
rect 25490 2692 25514 2694
rect 25570 2692 25576 2694
rect 25268 2683 25576 2692
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 800 7144 2246
rect 7898 2204 8206 2213
rect 7898 2202 7904 2204
rect 7960 2202 7984 2204
rect 8040 2202 8064 2204
rect 8120 2202 8144 2204
rect 8200 2202 8206 2204
rect 7960 2150 7962 2202
rect 8142 2150 8144 2202
rect 7898 2148 7904 2150
rect 7960 2148 7984 2150
rect 8040 2148 8064 2150
rect 8120 2148 8144 2150
rect 8200 2148 8206 2150
rect 7898 2139 8206 2148
rect 14846 2204 15154 2213
rect 14846 2202 14852 2204
rect 14908 2202 14932 2204
rect 14988 2202 15012 2204
rect 15068 2202 15092 2204
rect 15148 2202 15154 2204
rect 14908 2150 14910 2202
rect 15090 2150 15092 2202
rect 14846 2148 14852 2150
rect 14908 2148 14932 2150
rect 14988 2148 15012 2150
rect 15068 2148 15092 2150
rect 15148 2148 15154 2150
rect 14846 2139 15154 2148
rect 21794 2204 22102 2213
rect 21794 2202 21800 2204
rect 21856 2202 21880 2204
rect 21936 2202 21960 2204
rect 22016 2202 22040 2204
rect 22096 2202 22102 2204
rect 21856 2150 21858 2202
rect 22038 2150 22040 2202
rect 21794 2148 21800 2150
rect 21856 2148 21880 2150
rect 21936 2148 21960 2150
rect 22016 2148 22040 2150
rect 22096 2148 22102 2150
rect 21794 2139 22102 2148
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 29642 0 29698 800
<< via2 >>
rect 4430 27770 4486 27772
rect 4510 27770 4566 27772
rect 4590 27770 4646 27772
rect 4670 27770 4726 27772
rect 4430 27718 4476 27770
rect 4476 27718 4486 27770
rect 4510 27718 4540 27770
rect 4540 27718 4552 27770
rect 4552 27718 4566 27770
rect 4590 27718 4604 27770
rect 4604 27718 4616 27770
rect 4616 27718 4646 27770
rect 4670 27718 4680 27770
rect 4680 27718 4726 27770
rect 4430 27716 4486 27718
rect 4510 27716 4566 27718
rect 4590 27716 4646 27718
rect 4670 27716 4726 27718
rect 11378 27770 11434 27772
rect 11458 27770 11514 27772
rect 11538 27770 11594 27772
rect 11618 27770 11674 27772
rect 11378 27718 11424 27770
rect 11424 27718 11434 27770
rect 11458 27718 11488 27770
rect 11488 27718 11500 27770
rect 11500 27718 11514 27770
rect 11538 27718 11552 27770
rect 11552 27718 11564 27770
rect 11564 27718 11594 27770
rect 11618 27718 11628 27770
rect 11628 27718 11674 27770
rect 11378 27716 11434 27718
rect 11458 27716 11514 27718
rect 11538 27716 11594 27718
rect 11618 27716 11674 27718
rect 18326 27770 18382 27772
rect 18406 27770 18462 27772
rect 18486 27770 18542 27772
rect 18566 27770 18622 27772
rect 18326 27718 18372 27770
rect 18372 27718 18382 27770
rect 18406 27718 18436 27770
rect 18436 27718 18448 27770
rect 18448 27718 18462 27770
rect 18486 27718 18500 27770
rect 18500 27718 18512 27770
rect 18512 27718 18542 27770
rect 18566 27718 18576 27770
rect 18576 27718 18622 27770
rect 18326 27716 18382 27718
rect 18406 27716 18462 27718
rect 18486 27716 18542 27718
rect 18566 27716 18622 27718
rect 25274 27770 25330 27772
rect 25354 27770 25410 27772
rect 25434 27770 25490 27772
rect 25514 27770 25570 27772
rect 25274 27718 25320 27770
rect 25320 27718 25330 27770
rect 25354 27718 25384 27770
rect 25384 27718 25396 27770
rect 25396 27718 25410 27770
rect 25434 27718 25448 27770
rect 25448 27718 25460 27770
rect 25460 27718 25490 27770
rect 25514 27718 25524 27770
rect 25524 27718 25570 27770
rect 25274 27716 25330 27718
rect 25354 27716 25410 27718
rect 25434 27716 25490 27718
rect 25514 27716 25570 27718
rect 7904 27226 7960 27228
rect 7984 27226 8040 27228
rect 8064 27226 8120 27228
rect 8144 27226 8200 27228
rect 7904 27174 7950 27226
rect 7950 27174 7960 27226
rect 7984 27174 8014 27226
rect 8014 27174 8026 27226
rect 8026 27174 8040 27226
rect 8064 27174 8078 27226
rect 8078 27174 8090 27226
rect 8090 27174 8120 27226
rect 8144 27174 8154 27226
rect 8154 27174 8200 27226
rect 7904 27172 7960 27174
rect 7984 27172 8040 27174
rect 8064 27172 8120 27174
rect 8144 27172 8200 27174
rect 14852 27226 14908 27228
rect 14932 27226 14988 27228
rect 15012 27226 15068 27228
rect 15092 27226 15148 27228
rect 14852 27174 14898 27226
rect 14898 27174 14908 27226
rect 14932 27174 14962 27226
rect 14962 27174 14974 27226
rect 14974 27174 14988 27226
rect 15012 27174 15026 27226
rect 15026 27174 15038 27226
rect 15038 27174 15068 27226
rect 15092 27174 15102 27226
rect 15102 27174 15148 27226
rect 14852 27172 14908 27174
rect 14932 27172 14988 27174
rect 15012 27172 15068 27174
rect 15092 27172 15148 27174
rect 21800 27226 21856 27228
rect 21880 27226 21936 27228
rect 21960 27226 22016 27228
rect 22040 27226 22096 27228
rect 21800 27174 21846 27226
rect 21846 27174 21856 27226
rect 21880 27174 21910 27226
rect 21910 27174 21922 27226
rect 21922 27174 21936 27226
rect 21960 27174 21974 27226
rect 21974 27174 21986 27226
rect 21986 27174 22016 27226
rect 22040 27174 22050 27226
rect 22050 27174 22096 27226
rect 21800 27172 21856 27174
rect 21880 27172 21936 27174
rect 21960 27172 22016 27174
rect 22040 27172 22096 27174
rect 4430 26682 4486 26684
rect 4510 26682 4566 26684
rect 4590 26682 4646 26684
rect 4670 26682 4726 26684
rect 4430 26630 4476 26682
rect 4476 26630 4486 26682
rect 4510 26630 4540 26682
rect 4540 26630 4552 26682
rect 4552 26630 4566 26682
rect 4590 26630 4604 26682
rect 4604 26630 4616 26682
rect 4616 26630 4646 26682
rect 4670 26630 4680 26682
rect 4680 26630 4726 26682
rect 4430 26628 4486 26630
rect 4510 26628 4566 26630
rect 4590 26628 4646 26630
rect 4670 26628 4726 26630
rect 11378 26682 11434 26684
rect 11458 26682 11514 26684
rect 11538 26682 11594 26684
rect 11618 26682 11674 26684
rect 11378 26630 11424 26682
rect 11424 26630 11434 26682
rect 11458 26630 11488 26682
rect 11488 26630 11500 26682
rect 11500 26630 11514 26682
rect 11538 26630 11552 26682
rect 11552 26630 11564 26682
rect 11564 26630 11594 26682
rect 11618 26630 11628 26682
rect 11628 26630 11674 26682
rect 11378 26628 11434 26630
rect 11458 26628 11514 26630
rect 11538 26628 11594 26630
rect 11618 26628 11674 26630
rect 18326 26682 18382 26684
rect 18406 26682 18462 26684
rect 18486 26682 18542 26684
rect 18566 26682 18622 26684
rect 18326 26630 18372 26682
rect 18372 26630 18382 26682
rect 18406 26630 18436 26682
rect 18436 26630 18448 26682
rect 18448 26630 18462 26682
rect 18486 26630 18500 26682
rect 18500 26630 18512 26682
rect 18512 26630 18542 26682
rect 18566 26630 18576 26682
rect 18576 26630 18622 26682
rect 18326 26628 18382 26630
rect 18406 26628 18462 26630
rect 18486 26628 18542 26630
rect 18566 26628 18622 26630
rect 25274 26682 25330 26684
rect 25354 26682 25410 26684
rect 25434 26682 25490 26684
rect 25514 26682 25570 26684
rect 25274 26630 25320 26682
rect 25320 26630 25330 26682
rect 25354 26630 25384 26682
rect 25384 26630 25396 26682
rect 25396 26630 25410 26682
rect 25434 26630 25448 26682
rect 25448 26630 25460 26682
rect 25460 26630 25490 26682
rect 25514 26630 25524 26682
rect 25524 26630 25570 26682
rect 25274 26628 25330 26630
rect 25354 26628 25410 26630
rect 25434 26628 25490 26630
rect 25514 26628 25570 26630
rect 7904 26138 7960 26140
rect 7984 26138 8040 26140
rect 8064 26138 8120 26140
rect 8144 26138 8200 26140
rect 7904 26086 7950 26138
rect 7950 26086 7960 26138
rect 7984 26086 8014 26138
rect 8014 26086 8026 26138
rect 8026 26086 8040 26138
rect 8064 26086 8078 26138
rect 8078 26086 8090 26138
rect 8090 26086 8120 26138
rect 8144 26086 8154 26138
rect 8154 26086 8200 26138
rect 7904 26084 7960 26086
rect 7984 26084 8040 26086
rect 8064 26084 8120 26086
rect 8144 26084 8200 26086
rect 14852 26138 14908 26140
rect 14932 26138 14988 26140
rect 15012 26138 15068 26140
rect 15092 26138 15148 26140
rect 14852 26086 14898 26138
rect 14898 26086 14908 26138
rect 14932 26086 14962 26138
rect 14962 26086 14974 26138
rect 14974 26086 14988 26138
rect 15012 26086 15026 26138
rect 15026 26086 15038 26138
rect 15038 26086 15068 26138
rect 15092 26086 15102 26138
rect 15102 26086 15148 26138
rect 14852 26084 14908 26086
rect 14932 26084 14988 26086
rect 15012 26084 15068 26086
rect 15092 26084 15148 26086
rect 21800 26138 21856 26140
rect 21880 26138 21936 26140
rect 21960 26138 22016 26140
rect 22040 26138 22096 26140
rect 21800 26086 21846 26138
rect 21846 26086 21856 26138
rect 21880 26086 21910 26138
rect 21910 26086 21922 26138
rect 21922 26086 21936 26138
rect 21960 26086 21974 26138
rect 21974 26086 21986 26138
rect 21986 26086 22016 26138
rect 22040 26086 22050 26138
rect 22050 26086 22096 26138
rect 21800 26084 21856 26086
rect 21880 26084 21936 26086
rect 21960 26084 22016 26086
rect 22040 26084 22096 26086
rect 4430 25594 4486 25596
rect 4510 25594 4566 25596
rect 4590 25594 4646 25596
rect 4670 25594 4726 25596
rect 4430 25542 4476 25594
rect 4476 25542 4486 25594
rect 4510 25542 4540 25594
rect 4540 25542 4552 25594
rect 4552 25542 4566 25594
rect 4590 25542 4604 25594
rect 4604 25542 4616 25594
rect 4616 25542 4646 25594
rect 4670 25542 4680 25594
rect 4680 25542 4726 25594
rect 4430 25540 4486 25542
rect 4510 25540 4566 25542
rect 4590 25540 4646 25542
rect 4670 25540 4726 25542
rect 11378 25594 11434 25596
rect 11458 25594 11514 25596
rect 11538 25594 11594 25596
rect 11618 25594 11674 25596
rect 11378 25542 11424 25594
rect 11424 25542 11434 25594
rect 11458 25542 11488 25594
rect 11488 25542 11500 25594
rect 11500 25542 11514 25594
rect 11538 25542 11552 25594
rect 11552 25542 11564 25594
rect 11564 25542 11594 25594
rect 11618 25542 11628 25594
rect 11628 25542 11674 25594
rect 11378 25540 11434 25542
rect 11458 25540 11514 25542
rect 11538 25540 11594 25542
rect 11618 25540 11674 25542
rect 18326 25594 18382 25596
rect 18406 25594 18462 25596
rect 18486 25594 18542 25596
rect 18566 25594 18622 25596
rect 18326 25542 18372 25594
rect 18372 25542 18382 25594
rect 18406 25542 18436 25594
rect 18436 25542 18448 25594
rect 18448 25542 18462 25594
rect 18486 25542 18500 25594
rect 18500 25542 18512 25594
rect 18512 25542 18542 25594
rect 18566 25542 18576 25594
rect 18576 25542 18622 25594
rect 18326 25540 18382 25542
rect 18406 25540 18462 25542
rect 18486 25540 18542 25542
rect 18566 25540 18622 25542
rect 25274 25594 25330 25596
rect 25354 25594 25410 25596
rect 25434 25594 25490 25596
rect 25514 25594 25570 25596
rect 25274 25542 25320 25594
rect 25320 25542 25330 25594
rect 25354 25542 25384 25594
rect 25384 25542 25396 25594
rect 25396 25542 25410 25594
rect 25434 25542 25448 25594
rect 25448 25542 25460 25594
rect 25460 25542 25490 25594
rect 25514 25542 25524 25594
rect 25524 25542 25570 25594
rect 25274 25540 25330 25542
rect 25354 25540 25410 25542
rect 25434 25540 25490 25542
rect 25514 25540 25570 25542
rect 7904 25050 7960 25052
rect 7984 25050 8040 25052
rect 8064 25050 8120 25052
rect 8144 25050 8200 25052
rect 7904 24998 7950 25050
rect 7950 24998 7960 25050
rect 7984 24998 8014 25050
rect 8014 24998 8026 25050
rect 8026 24998 8040 25050
rect 8064 24998 8078 25050
rect 8078 24998 8090 25050
rect 8090 24998 8120 25050
rect 8144 24998 8154 25050
rect 8154 24998 8200 25050
rect 7904 24996 7960 24998
rect 7984 24996 8040 24998
rect 8064 24996 8120 24998
rect 8144 24996 8200 24998
rect 14852 25050 14908 25052
rect 14932 25050 14988 25052
rect 15012 25050 15068 25052
rect 15092 25050 15148 25052
rect 14852 24998 14898 25050
rect 14898 24998 14908 25050
rect 14932 24998 14962 25050
rect 14962 24998 14974 25050
rect 14974 24998 14988 25050
rect 15012 24998 15026 25050
rect 15026 24998 15038 25050
rect 15038 24998 15068 25050
rect 15092 24998 15102 25050
rect 15102 24998 15148 25050
rect 14852 24996 14908 24998
rect 14932 24996 14988 24998
rect 15012 24996 15068 24998
rect 15092 24996 15148 24998
rect 21800 25050 21856 25052
rect 21880 25050 21936 25052
rect 21960 25050 22016 25052
rect 22040 25050 22096 25052
rect 21800 24998 21846 25050
rect 21846 24998 21856 25050
rect 21880 24998 21910 25050
rect 21910 24998 21922 25050
rect 21922 24998 21936 25050
rect 21960 24998 21974 25050
rect 21974 24998 21986 25050
rect 21986 24998 22016 25050
rect 22040 24998 22050 25050
rect 22050 24998 22096 25050
rect 21800 24996 21856 24998
rect 21880 24996 21936 24998
rect 21960 24996 22016 24998
rect 22040 24996 22096 24998
rect 4430 24506 4486 24508
rect 4510 24506 4566 24508
rect 4590 24506 4646 24508
rect 4670 24506 4726 24508
rect 4430 24454 4476 24506
rect 4476 24454 4486 24506
rect 4510 24454 4540 24506
rect 4540 24454 4552 24506
rect 4552 24454 4566 24506
rect 4590 24454 4604 24506
rect 4604 24454 4616 24506
rect 4616 24454 4646 24506
rect 4670 24454 4680 24506
rect 4680 24454 4726 24506
rect 4430 24452 4486 24454
rect 4510 24452 4566 24454
rect 4590 24452 4646 24454
rect 4670 24452 4726 24454
rect 11378 24506 11434 24508
rect 11458 24506 11514 24508
rect 11538 24506 11594 24508
rect 11618 24506 11674 24508
rect 11378 24454 11424 24506
rect 11424 24454 11434 24506
rect 11458 24454 11488 24506
rect 11488 24454 11500 24506
rect 11500 24454 11514 24506
rect 11538 24454 11552 24506
rect 11552 24454 11564 24506
rect 11564 24454 11594 24506
rect 11618 24454 11628 24506
rect 11628 24454 11674 24506
rect 11378 24452 11434 24454
rect 11458 24452 11514 24454
rect 11538 24452 11594 24454
rect 11618 24452 11674 24454
rect 18326 24506 18382 24508
rect 18406 24506 18462 24508
rect 18486 24506 18542 24508
rect 18566 24506 18622 24508
rect 18326 24454 18372 24506
rect 18372 24454 18382 24506
rect 18406 24454 18436 24506
rect 18436 24454 18448 24506
rect 18448 24454 18462 24506
rect 18486 24454 18500 24506
rect 18500 24454 18512 24506
rect 18512 24454 18542 24506
rect 18566 24454 18576 24506
rect 18576 24454 18622 24506
rect 18326 24452 18382 24454
rect 18406 24452 18462 24454
rect 18486 24452 18542 24454
rect 18566 24452 18622 24454
rect 25274 24506 25330 24508
rect 25354 24506 25410 24508
rect 25434 24506 25490 24508
rect 25514 24506 25570 24508
rect 25274 24454 25320 24506
rect 25320 24454 25330 24506
rect 25354 24454 25384 24506
rect 25384 24454 25396 24506
rect 25396 24454 25410 24506
rect 25434 24454 25448 24506
rect 25448 24454 25460 24506
rect 25460 24454 25490 24506
rect 25514 24454 25524 24506
rect 25524 24454 25570 24506
rect 25274 24452 25330 24454
rect 25354 24452 25410 24454
rect 25434 24452 25490 24454
rect 25514 24452 25570 24454
rect 7904 23962 7960 23964
rect 7984 23962 8040 23964
rect 8064 23962 8120 23964
rect 8144 23962 8200 23964
rect 7904 23910 7950 23962
rect 7950 23910 7960 23962
rect 7984 23910 8014 23962
rect 8014 23910 8026 23962
rect 8026 23910 8040 23962
rect 8064 23910 8078 23962
rect 8078 23910 8090 23962
rect 8090 23910 8120 23962
rect 8144 23910 8154 23962
rect 8154 23910 8200 23962
rect 7904 23908 7960 23910
rect 7984 23908 8040 23910
rect 8064 23908 8120 23910
rect 8144 23908 8200 23910
rect 14852 23962 14908 23964
rect 14932 23962 14988 23964
rect 15012 23962 15068 23964
rect 15092 23962 15148 23964
rect 14852 23910 14898 23962
rect 14898 23910 14908 23962
rect 14932 23910 14962 23962
rect 14962 23910 14974 23962
rect 14974 23910 14988 23962
rect 15012 23910 15026 23962
rect 15026 23910 15038 23962
rect 15038 23910 15068 23962
rect 15092 23910 15102 23962
rect 15102 23910 15148 23962
rect 14852 23908 14908 23910
rect 14932 23908 14988 23910
rect 15012 23908 15068 23910
rect 15092 23908 15148 23910
rect 21800 23962 21856 23964
rect 21880 23962 21936 23964
rect 21960 23962 22016 23964
rect 22040 23962 22096 23964
rect 21800 23910 21846 23962
rect 21846 23910 21856 23962
rect 21880 23910 21910 23962
rect 21910 23910 21922 23962
rect 21922 23910 21936 23962
rect 21960 23910 21974 23962
rect 21974 23910 21986 23962
rect 21986 23910 22016 23962
rect 22040 23910 22050 23962
rect 22050 23910 22096 23962
rect 21800 23908 21856 23910
rect 21880 23908 21936 23910
rect 21960 23908 22016 23910
rect 22040 23908 22096 23910
rect 4430 23418 4486 23420
rect 4510 23418 4566 23420
rect 4590 23418 4646 23420
rect 4670 23418 4726 23420
rect 4430 23366 4476 23418
rect 4476 23366 4486 23418
rect 4510 23366 4540 23418
rect 4540 23366 4552 23418
rect 4552 23366 4566 23418
rect 4590 23366 4604 23418
rect 4604 23366 4616 23418
rect 4616 23366 4646 23418
rect 4670 23366 4680 23418
rect 4680 23366 4726 23418
rect 4430 23364 4486 23366
rect 4510 23364 4566 23366
rect 4590 23364 4646 23366
rect 4670 23364 4726 23366
rect 11378 23418 11434 23420
rect 11458 23418 11514 23420
rect 11538 23418 11594 23420
rect 11618 23418 11674 23420
rect 11378 23366 11424 23418
rect 11424 23366 11434 23418
rect 11458 23366 11488 23418
rect 11488 23366 11500 23418
rect 11500 23366 11514 23418
rect 11538 23366 11552 23418
rect 11552 23366 11564 23418
rect 11564 23366 11594 23418
rect 11618 23366 11628 23418
rect 11628 23366 11674 23418
rect 11378 23364 11434 23366
rect 11458 23364 11514 23366
rect 11538 23364 11594 23366
rect 11618 23364 11674 23366
rect 18326 23418 18382 23420
rect 18406 23418 18462 23420
rect 18486 23418 18542 23420
rect 18566 23418 18622 23420
rect 18326 23366 18372 23418
rect 18372 23366 18382 23418
rect 18406 23366 18436 23418
rect 18436 23366 18448 23418
rect 18448 23366 18462 23418
rect 18486 23366 18500 23418
rect 18500 23366 18512 23418
rect 18512 23366 18542 23418
rect 18566 23366 18576 23418
rect 18576 23366 18622 23418
rect 18326 23364 18382 23366
rect 18406 23364 18462 23366
rect 18486 23364 18542 23366
rect 18566 23364 18622 23366
rect 25274 23418 25330 23420
rect 25354 23418 25410 23420
rect 25434 23418 25490 23420
rect 25514 23418 25570 23420
rect 25274 23366 25320 23418
rect 25320 23366 25330 23418
rect 25354 23366 25384 23418
rect 25384 23366 25396 23418
rect 25396 23366 25410 23418
rect 25434 23366 25448 23418
rect 25448 23366 25460 23418
rect 25460 23366 25490 23418
rect 25514 23366 25524 23418
rect 25524 23366 25570 23418
rect 25274 23364 25330 23366
rect 25354 23364 25410 23366
rect 25434 23364 25490 23366
rect 25514 23364 25570 23366
rect 7904 22874 7960 22876
rect 7984 22874 8040 22876
rect 8064 22874 8120 22876
rect 8144 22874 8200 22876
rect 7904 22822 7950 22874
rect 7950 22822 7960 22874
rect 7984 22822 8014 22874
rect 8014 22822 8026 22874
rect 8026 22822 8040 22874
rect 8064 22822 8078 22874
rect 8078 22822 8090 22874
rect 8090 22822 8120 22874
rect 8144 22822 8154 22874
rect 8154 22822 8200 22874
rect 7904 22820 7960 22822
rect 7984 22820 8040 22822
rect 8064 22820 8120 22822
rect 8144 22820 8200 22822
rect 14852 22874 14908 22876
rect 14932 22874 14988 22876
rect 15012 22874 15068 22876
rect 15092 22874 15148 22876
rect 14852 22822 14898 22874
rect 14898 22822 14908 22874
rect 14932 22822 14962 22874
rect 14962 22822 14974 22874
rect 14974 22822 14988 22874
rect 15012 22822 15026 22874
rect 15026 22822 15038 22874
rect 15038 22822 15068 22874
rect 15092 22822 15102 22874
rect 15102 22822 15148 22874
rect 14852 22820 14908 22822
rect 14932 22820 14988 22822
rect 15012 22820 15068 22822
rect 15092 22820 15148 22822
rect 21800 22874 21856 22876
rect 21880 22874 21936 22876
rect 21960 22874 22016 22876
rect 22040 22874 22096 22876
rect 21800 22822 21846 22874
rect 21846 22822 21856 22874
rect 21880 22822 21910 22874
rect 21910 22822 21922 22874
rect 21922 22822 21936 22874
rect 21960 22822 21974 22874
rect 21974 22822 21986 22874
rect 21986 22822 22016 22874
rect 22040 22822 22050 22874
rect 22050 22822 22096 22874
rect 21800 22820 21856 22822
rect 21880 22820 21936 22822
rect 21960 22820 22016 22822
rect 22040 22820 22096 22822
rect 4430 22330 4486 22332
rect 4510 22330 4566 22332
rect 4590 22330 4646 22332
rect 4670 22330 4726 22332
rect 4430 22278 4476 22330
rect 4476 22278 4486 22330
rect 4510 22278 4540 22330
rect 4540 22278 4552 22330
rect 4552 22278 4566 22330
rect 4590 22278 4604 22330
rect 4604 22278 4616 22330
rect 4616 22278 4646 22330
rect 4670 22278 4680 22330
rect 4680 22278 4726 22330
rect 4430 22276 4486 22278
rect 4510 22276 4566 22278
rect 4590 22276 4646 22278
rect 4670 22276 4726 22278
rect 11378 22330 11434 22332
rect 11458 22330 11514 22332
rect 11538 22330 11594 22332
rect 11618 22330 11674 22332
rect 11378 22278 11424 22330
rect 11424 22278 11434 22330
rect 11458 22278 11488 22330
rect 11488 22278 11500 22330
rect 11500 22278 11514 22330
rect 11538 22278 11552 22330
rect 11552 22278 11564 22330
rect 11564 22278 11594 22330
rect 11618 22278 11628 22330
rect 11628 22278 11674 22330
rect 11378 22276 11434 22278
rect 11458 22276 11514 22278
rect 11538 22276 11594 22278
rect 11618 22276 11674 22278
rect 18326 22330 18382 22332
rect 18406 22330 18462 22332
rect 18486 22330 18542 22332
rect 18566 22330 18622 22332
rect 18326 22278 18372 22330
rect 18372 22278 18382 22330
rect 18406 22278 18436 22330
rect 18436 22278 18448 22330
rect 18448 22278 18462 22330
rect 18486 22278 18500 22330
rect 18500 22278 18512 22330
rect 18512 22278 18542 22330
rect 18566 22278 18576 22330
rect 18576 22278 18622 22330
rect 18326 22276 18382 22278
rect 18406 22276 18462 22278
rect 18486 22276 18542 22278
rect 18566 22276 18622 22278
rect 25274 22330 25330 22332
rect 25354 22330 25410 22332
rect 25434 22330 25490 22332
rect 25514 22330 25570 22332
rect 25274 22278 25320 22330
rect 25320 22278 25330 22330
rect 25354 22278 25384 22330
rect 25384 22278 25396 22330
rect 25396 22278 25410 22330
rect 25434 22278 25448 22330
rect 25448 22278 25460 22330
rect 25460 22278 25490 22330
rect 25514 22278 25524 22330
rect 25524 22278 25570 22330
rect 25274 22276 25330 22278
rect 25354 22276 25410 22278
rect 25434 22276 25490 22278
rect 25514 22276 25570 22278
rect 7904 21786 7960 21788
rect 7984 21786 8040 21788
rect 8064 21786 8120 21788
rect 8144 21786 8200 21788
rect 7904 21734 7950 21786
rect 7950 21734 7960 21786
rect 7984 21734 8014 21786
rect 8014 21734 8026 21786
rect 8026 21734 8040 21786
rect 8064 21734 8078 21786
rect 8078 21734 8090 21786
rect 8090 21734 8120 21786
rect 8144 21734 8154 21786
rect 8154 21734 8200 21786
rect 7904 21732 7960 21734
rect 7984 21732 8040 21734
rect 8064 21732 8120 21734
rect 8144 21732 8200 21734
rect 14852 21786 14908 21788
rect 14932 21786 14988 21788
rect 15012 21786 15068 21788
rect 15092 21786 15148 21788
rect 14852 21734 14898 21786
rect 14898 21734 14908 21786
rect 14932 21734 14962 21786
rect 14962 21734 14974 21786
rect 14974 21734 14988 21786
rect 15012 21734 15026 21786
rect 15026 21734 15038 21786
rect 15038 21734 15068 21786
rect 15092 21734 15102 21786
rect 15102 21734 15148 21786
rect 14852 21732 14908 21734
rect 14932 21732 14988 21734
rect 15012 21732 15068 21734
rect 15092 21732 15148 21734
rect 21800 21786 21856 21788
rect 21880 21786 21936 21788
rect 21960 21786 22016 21788
rect 22040 21786 22096 21788
rect 21800 21734 21846 21786
rect 21846 21734 21856 21786
rect 21880 21734 21910 21786
rect 21910 21734 21922 21786
rect 21922 21734 21936 21786
rect 21960 21734 21974 21786
rect 21974 21734 21986 21786
rect 21986 21734 22016 21786
rect 22040 21734 22050 21786
rect 22050 21734 22096 21786
rect 21800 21732 21856 21734
rect 21880 21732 21936 21734
rect 21960 21732 22016 21734
rect 22040 21732 22096 21734
rect 4430 21242 4486 21244
rect 4510 21242 4566 21244
rect 4590 21242 4646 21244
rect 4670 21242 4726 21244
rect 4430 21190 4476 21242
rect 4476 21190 4486 21242
rect 4510 21190 4540 21242
rect 4540 21190 4552 21242
rect 4552 21190 4566 21242
rect 4590 21190 4604 21242
rect 4604 21190 4616 21242
rect 4616 21190 4646 21242
rect 4670 21190 4680 21242
rect 4680 21190 4726 21242
rect 4430 21188 4486 21190
rect 4510 21188 4566 21190
rect 4590 21188 4646 21190
rect 4670 21188 4726 21190
rect 11378 21242 11434 21244
rect 11458 21242 11514 21244
rect 11538 21242 11594 21244
rect 11618 21242 11674 21244
rect 11378 21190 11424 21242
rect 11424 21190 11434 21242
rect 11458 21190 11488 21242
rect 11488 21190 11500 21242
rect 11500 21190 11514 21242
rect 11538 21190 11552 21242
rect 11552 21190 11564 21242
rect 11564 21190 11594 21242
rect 11618 21190 11628 21242
rect 11628 21190 11674 21242
rect 11378 21188 11434 21190
rect 11458 21188 11514 21190
rect 11538 21188 11594 21190
rect 11618 21188 11674 21190
rect 18326 21242 18382 21244
rect 18406 21242 18462 21244
rect 18486 21242 18542 21244
rect 18566 21242 18622 21244
rect 18326 21190 18372 21242
rect 18372 21190 18382 21242
rect 18406 21190 18436 21242
rect 18436 21190 18448 21242
rect 18448 21190 18462 21242
rect 18486 21190 18500 21242
rect 18500 21190 18512 21242
rect 18512 21190 18542 21242
rect 18566 21190 18576 21242
rect 18576 21190 18622 21242
rect 18326 21188 18382 21190
rect 18406 21188 18462 21190
rect 18486 21188 18542 21190
rect 18566 21188 18622 21190
rect 25274 21242 25330 21244
rect 25354 21242 25410 21244
rect 25434 21242 25490 21244
rect 25514 21242 25570 21244
rect 25274 21190 25320 21242
rect 25320 21190 25330 21242
rect 25354 21190 25384 21242
rect 25384 21190 25396 21242
rect 25396 21190 25410 21242
rect 25434 21190 25448 21242
rect 25448 21190 25460 21242
rect 25460 21190 25490 21242
rect 25514 21190 25524 21242
rect 25524 21190 25570 21242
rect 25274 21188 25330 21190
rect 25354 21188 25410 21190
rect 25434 21188 25490 21190
rect 25514 21188 25570 21190
rect 7904 20698 7960 20700
rect 7984 20698 8040 20700
rect 8064 20698 8120 20700
rect 8144 20698 8200 20700
rect 7904 20646 7950 20698
rect 7950 20646 7960 20698
rect 7984 20646 8014 20698
rect 8014 20646 8026 20698
rect 8026 20646 8040 20698
rect 8064 20646 8078 20698
rect 8078 20646 8090 20698
rect 8090 20646 8120 20698
rect 8144 20646 8154 20698
rect 8154 20646 8200 20698
rect 7904 20644 7960 20646
rect 7984 20644 8040 20646
rect 8064 20644 8120 20646
rect 8144 20644 8200 20646
rect 14852 20698 14908 20700
rect 14932 20698 14988 20700
rect 15012 20698 15068 20700
rect 15092 20698 15148 20700
rect 14852 20646 14898 20698
rect 14898 20646 14908 20698
rect 14932 20646 14962 20698
rect 14962 20646 14974 20698
rect 14974 20646 14988 20698
rect 15012 20646 15026 20698
rect 15026 20646 15038 20698
rect 15038 20646 15068 20698
rect 15092 20646 15102 20698
rect 15102 20646 15148 20698
rect 14852 20644 14908 20646
rect 14932 20644 14988 20646
rect 15012 20644 15068 20646
rect 15092 20644 15148 20646
rect 21800 20698 21856 20700
rect 21880 20698 21936 20700
rect 21960 20698 22016 20700
rect 22040 20698 22096 20700
rect 21800 20646 21846 20698
rect 21846 20646 21856 20698
rect 21880 20646 21910 20698
rect 21910 20646 21922 20698
rect 21922 20646 21936 20698
rect 21960 20646 21974 20698
rect 21974 20646 21986 20698
rect 21986 20646 22016 20698
rect 22040 20646 22050 20698
rect 22050 20646 22096 20698
rect 21800 20644 21856 20646
rect 21880 20644 21936 20646
rect 21960 20644 22016 20646
rect 22040 20644 22096 20646
rect 4430 20154 4486 20156
rect 4510 20154 4566 20156
rect 4590 20154 4646 20156
rect 4670 20154 4726 20156
rect 4430 20102 4476 20154
rect 4476 20102 4486 20154
rect 4510 20102 4540 20154
rect 4540 20102 4552 20154
rect 4552 20102 4566 20154
rect 4590 20102 4604 20154
rect 4604 20102 4616 20154
rect 4616 20102 4646 20154
rect 4670 20102 4680 20154
rect 4680 20102 4726 20154
rect 4430 20100 4486 20102
rect 4510 20100 4566 20102
rect 4590 20100 4646 20102
rect 4670 20100 4726 20102
rect 11378 20154 11434 20156
rect 11458 20154 11514 20156
rect 11538 20154 11594 20156
rect 11618 20154 11674 20156
rect 11378 20102 11424 20154
rect 11424 20102 11434 20154
rect 11458 20102 11488 20154
rect 11488 20102 11500 20154
rect 11500 20102 11514 20154
rect 11538 20102 11552 20154
rect 11552 20102 11564 20154
rect 11564 20102 11594 20154
rect 11618 20102 11628 20154
rect 11628 20102 11674 20154
rect 11378 20100 11434 20102
rect 11458 20100 11514 20102
rect 11538 20100 11594 20102
rect 11618 20100 11674 20102
rect 18326 20154 18382 20156
rect 18406 20154 18462 20156
rect 18486 20154 18542 20156
rect 18566 20154 18622 20156
rect 18326 20102 18372 20154
rect 18372 20102 18382 20154
rect 18406 20102 18436 20154
rect 18436 20102 18448 20154
rect 18448 20102 18462 20154
rect 18486 20102 18500 20154
rect 18500 20102 18512 20154
rect 18512 20102 18542 20154
rect 18566 20102 18576 20154
rect 18576 20102 18622 20154
rect 18326 20100 18382 20102
rect 18406 20100 18462 20102
rect 18486 20100 18542 20102
rect 18566 20100 18622 20102
rect 25274 20154 25330 20156
rect 25354 20154 25410 20156
rect 25434 20154 25490 20156
rect 25514 20154 25570 20156
rect 25274 20102 25320 20154
rect 25320 20102 25330 20154
rect 25354 20102 25384 20154
rect 25384 20102 25396 20154
rect 25396 20102 25410 20154
rect 25434 20102 25448 20154
rect 25448 20102 25460 20154
rect 25460 20102 25490 20154
rect 25514 20102 25524 20154
rect 25524 20102 25570 20154
rect 25274 20100 25330 20102
rect 25354 20100 25410 20102
rect 25434 20100 25490 20102
rect 25514 20100 25570 20102
rect 7904 19610 7960 19612
rect 7984 19610 8040 19612
rect 8064 19610 8120 19612
rect 8144 19610 8200 19612
rect 7904 19558 7950 19610
rect 7950 19558 7960 19610
rect 7984 19558 8014 19610
rect 8014 19558 8026 19610
rect 8026 19558 8040 19610
rect 8064 19558 8078 19610
rect 8078 19558 8090 19610
rect 8090 19558 8120 19610
rect 8144 19558 8154 19610
rect 8154 19558 8200 19610
rect 7904 19556 7960 19558
rect 7984 19556 8040 19558
rect 8064 19556 8120 19558
rect 8144 19556 8200 19558
rect 14852 19610 14908 19612
rect 14932 19610 14988 19612
rect 15012 19610 15068 19612
rect 15092 19610 15148 19612
rect 14852 19558 14898 19610
rect 14898 19558 14908 19610
rect 14932 19558 14962 19610
rect 14962 19558 14974 19610
rect 14974 19558 14988 19610
rect 15012 19558 15026 19610
rect 15026 19558 15038 19610
rect 15038 19558 15068 19610
rect 15092 19558 15102 19610
rect 15102 19558 15148 19610
rect 14852 19556 14908 19558
rect 14932 19556 14988 19558
rect 15012 19556 15068 19558
rect 15092 19556 15148 19558
rect 21800 19610 21856 19612
rect 21880 19610 21936 19612
rect 21960 19610 22016 19612
rect 22040 19610 22096 19612
rect 21800 19558 21846 19610
rect 21846 19558 21856 19610
rect 21880 19558 21910 19610
rect 21910 19558 21922 19610
rect 21922 19558 21936 19610
rect 21960 19558 21974 19610
rect 21974 19558 21986 19610
rect 21986 19558 22016 19610
rect 22040 19558 22050 19610
rect 22050 19558 22096 19610
rect 21800 19556 21856 19558
rect 21880 19556 21936 19558
rect 21960 19556 22016 19558
rect 22040 19556 22096 19558
rect 4430 19066 4486 19068
rect 4510 19066 4566 19068
rect 4590 19066 4646 19068
rect 4670 19066 4726 19068
rect 4430 19014 4476 19066
rect 4476 19014 4486 19066
rect 4510 19014 4540 19066
rect 4540 19014 4552 19066
rect 4552 19014 4566 19066
rect 4590 19014 4604 19066
rect 4604 19014 4616 19066
rect 4616 19014 4646 19066
rect 4670 19014 4680 19066
rect 4680 19014 4726 19066
rect 4430 19012 4486 19014
rect 4510 19012 4566 19014
rect 4590 19012 4646 19014
rect 4670 19012 4726 19014
rect 11378 19066 11434 19068
rect 11458 19066 11514 19068
rect 11538 19066 11594 19068
rect 11618 19066 11674 19068
rect 11378 19014 11424 19066
rect 11424 19014 11434 19066
rect 11458 19014 11488 19066
rect 11488 19014 11500 19066
rect 11500 19014 11514 19066
rect 11538 19014 11552 19066
rect 11552 19014 11564 19066
rect 11564 19014 11594 19066
rect 11618 19014 11628 19066
rect 11628 19014 11674 19066
rect 11378 19012 11434 19014
rect 11458 19012 11514 19014
rect 11538 19012 11594 19014
rect 11618 19012 11674 19014
rect 18326 19066 18382 19068
rect 18406 19066 18462 19068
rect 18486 19066 18542 19068
rect 18566 19066 18622 19068
rect 18326 19014 18372 19066
rect 18372 19014 18382 19066
rect 18406 19014 18436 19066
rect 18436 19014 18448 19066
rect 18448 19014 18462 19066
rect 18486 19014 18500 19066
rect 18500 19014 18512 19066
rect 18512 19014 18542 19066
rect 18566 19014 18576 19066
rect 18576 19014 18622 19066
rect 18326 19012 18382 19014
rect 18406 19012 18462 19014
rect 18486 19012 18542 19014
rect 18566 19012 18622 19014
rect 25274 19066 25330 19068
rect 25354 19066 25410 19068
rect 25434 19066 25490 19068
rect 25514 19066 25570 19068
rect 25274 19014 25320 19066
rect 25320 19014 25330 19066
rect 25354 19014 25384 19066
rect 25384 19014 25396 19066
rect 25396 19014 25410 19066
rect 25434 19014 25448 19066
rect 25448 19014 25460 19066
rect 25460 19014 25490 19066
rect 25514 19014 25524 19066
rect 25524 19014 25570 19066
rect 25274 19012 25330 19014
rect 25354 19012 25410 19014
rect 25434 19012 25490 19014
rect 25514 19012 25570 19014
rect 7904 18522 7960 18524
rect 7984 18522 8040 18524
rect 8064 18522 8120 18524
rect 8144 18522 8200 18524
rect 7904 18470 7950 18522
rect 7950 18470 7960 18522
rect 7984 18470 8014 18522
rect 8014 18470 8026 18522
rect 8026 18470 8040 18522
rect 8064 18470 8078 18522
rect 8078 18470 8090 18522
rect 8090 18470 8120 18522
rect 8144 18470 8154 18522
rect 8154 18470 8200 18522
rect 7904 18468 7960 18470
rect 7984 18468 8040 18470
rect 8064 18468 8120 18470
rect 8144 18468 8200 18470
rect 14852 18522 14908 18524
rect 14932 18522 14988 18524
rect 15012 18522 15068 18524
rect 15092 18522 15148 18524
rect 14852 18470 14898 18522
rect 14898 18470 14908 18522
rect 14932 18470 14962 18522
rect 14962 18470 14974 18522
rect 14974 18470 14988 18522
rect 15012 18470 15026 18522
rect 15026 18470 15038 18522
rect 15038 18470 15068 18522
rect 15092 18470 15102 18522
rect 15102 18470 15148 18522
rect 14852 18468 14908 18470
rect 14932 18468 14988 18470
rect 15012 18468 15068 18470
rect 15092 18468 15148 18470
rect 21800 18522 21856 18524
rect 21880 18522 21936 18524
rect 21960 18522 22016 18524
rect 22040 18522 22096 18524
rect 21800 18470 21846 18522
rect 21846 18470 21856 18522
rect 21880 18470 21910 18522
rect 21910 18470 21922 18522
rect 21922 18470 21936 18522
rect 21960 18470 21974 18522
rect 21974 18470 21986 18522
rect 21986 18470 22016 18522
rect 22040 18470 22050 18522
rect 22050 18470 22096 18522
rect 21800 18468 21856 18470
rect 21880 18468 21936 18470
rect 21960 18468 22016 18470
rect 22040 18468 22096 18470
rect 4430 17978 4486 17980
rect 4510 17978 4566 17980
rect 4590 17978 4646 17980
rect 4670 17978 4726 17980
rect 4430 17926 4476 17978
rect 4476 17926 4486 17978
rect 4510 17926 4540 17978
rect 4540 17926 4552 17978
rect 4552 17926 4566 17978
rect 4590 17926 4604 17978
rect 4604 17926 4616 17978
rect 4616 17926 4646 17978
rect 4670 17926 4680 17978
rect 4680 17926 4726 17978
rect 4430 17924 4486 17926
rect 4510 17924 4566 17926
rect 4590 17924 4646 17926
rect 4670 17924 4726 17926
rect 11378 17978 11434 17980
rect 11458 17978 11514 17980
rect 11538 17978 11594 17980
rect 11618 17978 11674 17980
rect 11378 17926 11424 17978
rect 11424 17926 11434 17978
rect 11458 17926 11488 17978
rect 11488 17926 11500 17978
rect 11500 17926 11514 17978
rect 11538 17926 11552 17978
rect 11552 17926 11564 17978
rect 11564 17926 11594 17978
rect 11618 17926 11628 17978
rect 11628 17926 11674 17978
rect 11378 17924 11434 17926
rect 11458 17924 11514 17926
rect 11538 17924 11594 17926
rect 11618 17924 11674 17926
rect 18326 17978 18382 17980
rect 18406 17978 18462 17980
rect 18486 17978 18542 17980
rect 18566 17978 18622 17980
rect 18326 17926 18372 17978
rect 18372 17926 18382 17978
rect 18406 17926 18436 17978
rect 18436 17926 18448 17978
rect 18448 17926 18462 17978
rect 18486 17926 18500 17978
rect 18500 17926 18512 17978
rect 18512 17926 18542 17978
rect 18566 17926 18576 17978
rect 18576 17926 18622 17978
rect 18326 17924 18382 17926
rect 18406 17924 18462 17926
rect 18486 17924 18542 17926
rect 18566 17924 18622 17926
rect 25274 17978 25330 17980
rect 25354 17978 25410 17980
rect 25434 17978 25490 17980
rect 25514 17978 25570 17980
rect 25274 17926 25320 17978
rect 25320 17926 25330 17978
rect 25354 17926 25384 17978
rect 25384 17926 25396 17978
rect 25396 17926 25410 17978
rect 25434 17926 25448 17978
rect 25448 17926 25460 17978
rect 25460 17926 25490 17978
rect 25514 17926 25524 17978
rect 25524 17926 25570 17978
rect 25274 17924 25330 17926
rect 25354 17924 25410 17926
rect 25434 17924 25490 17926
rect 25514 17924 25570 17926
rect 7904 17434 7960 17436
rect 7984 17434 8040 17436
rect 8064 17434 8120 17436
rect 8144 17434 8200 17436
rect 7904 17382 7950 17434
rect 7950 17382 7960 17434
rect 7984 17382 8014 17434
rect 8014 17382 8026 17434
rect 8026 17382 8040 17434
rect 8064 17382 8078 17434
rect 8078 17382 8090 17434
rect 8090 17382 8120 17434
rect 8144 17382 8154 17434
rect 8154 17382 8200 17434
rect 7904 17380 7960 17382
rect 7984 17380 8040 17382
rect 8064 17380 8120 17382
rect 8144 17380 8200 17382
rect 14852 17434 14908 17436
rect 14932 17434 14988 17436
rect 15012 17434 15068 17436
rect 15092 17434 15148 17436
rect 14852 17382 14898 17434
rect 14898 17382 14908 17434
rect 14932 17382 14962 17434
rect 14962 17382 14974 17434
rect 14974 17382 14988 17434
rect 15012 17382 15026 17434
rect 15026 17382 15038 17434
rect 15038 17382 15068 17434
rect 15092 17382 15102 17434
rect 15102 17382 15148 17434
rect 14852 17380 14908 17382
rect 14932 17380 14988 17382
rect 15012 17380 15068 17382
rect 15092 17380 15148 17382
rect 21800 17434 21856 17436
rect 21880 17434 21936 17436
rect 21960 17434 22016 17436
rect 22040 17434 22096 17436
rect 21800 17382 21846 17434
rect 21846 17382 21856 17434
rect 21880 17382 21910 17434
rect 21910 17382 21922 17434
rect 21922 17382 21936 17434
rect 21960 17382 21974 17434
rect 21974 17382 21986 17434
rect 21986 17382 22016 17434
rect 22040 17382 22050 17434
rect 22050 17382 22096 17434
rect 21800 17380 21856 17382
rect 21880 17380 21936 17382
rect 21960 17380 22016 17382
rect 22040 17380 22096 17382
rect 4430 16890 4486 16892
rect 4510 16890 4566 16892
rect 4590 16890 4646 16892
rect 4670 16890 4726 16892
rect 4430 16838 4476 16890
rect 4476 16838 4486 16890
rect 4510 16838 4540 16890
rect 4540 16838 4552 16890
rect 4552 16838 4566 16890
rect 4590 16838 4604 16890
rect 4604 16838 4616 16890
rect 4616 16838 4646 16890
rect 4670 16838 4680 16890
rect 4680 16838 4726 16890
rect 4430 16836 4486 16838
rect 4510 16836 4566 16838
rect 4590 16836 4646 16838
rect 4670 16836 4726 16838
rect 11378 16890 11434 16892
rect 11458 16890 11514 16892
rect 11538 16890 11594 16892
rect 11618 16890 11674 16892
rect 11378 16838 11424 16890
rect 11424 16838 11434 16890
rect 11458 16838 11488 16890
rect 11488 16838 11500 16890
rect 11500 16838 11514 16890
rect 11538 16838 11552 16890
rect 11552 16838 11564 16890
rect 11564 16838 11594 16890
rect 11618 16838 11628 16890
rect 11628 16838 11674 16890
rect 11378 16836 11434 16838
rect 11458 16836 11514 16838
rect 11538 16836 11594 16838
rect 11618 16836 11674 16838
rect 18326 16890 18382 16892
rect 18406 16890 18462 16892
rect 18486 16890 18542 16892
rect 18566 16890 18622 16892
rect 18326 16838 18372 16890
rect 18372 16838 18382 16890
rect 18406 16838 18436 16890
rect 18436 16838 18448 16890
rect 18448 16838 18462 16890
rect 18486 16838 18500 16890
rect 18500 16838 18512 16890
rect 18512 16838 18542 16890
rect 18566 16838 18576 16890
rect 18576 16838 18622 16890
rect 18326 16836 18382 16838
rect 18406 16836 18462 16838
rect 18486 16836 18542 16838
rect 18566 16836 18622 16838
rect 25274 16890 25330 16892
rect 25354 16890 25410 16892
rect 25434 16890 25490 16892
rect 25514 16890 25570 16892
rect 25274 16838 25320 16890
rect 25320 16838 25330 16890
rect 25354 16838 25384 16890
rect 25384 16838 25396 16890
rect 25396 16838 25410 16890
rect 25434 16838 25448 16890
rect 25448 16838 25460 16890
rect 25460 16838 25490 16890
rect 25514 16838 25524 16890
rect 25524 16838 25570 16890
rect 25274 16836 25330 16838
rect 25354 16836 25410 16838
rect 25434 16836 25490 16838
rect 25514 16836 25570 16838
rect 7904 16346 7960 16348
rect 7984 16346 8040 16348
rect 8064 16346 8120 16348
rect 8144 16346 8200 16348
rect 7904 16294 7950 16346
rect 7950 16294 7960 16346
rect 7984 16294 8014 16346
rect 8014 16294 8026 16346
rect 8026 16294 8040 16346
rect 8064 16294 8078 16346
rect 8078 16294 8090 16346
rect 8090 16294 8120 16346
rect 8144 16294 8154 16346
rect 8154 16294 8200 16346
rect 7904 16292 7960 16294
rect 7984 16292 8040 16294
rect 8064 16292 8120 16294
rect 8144 16292 8200 16294
rect 14852 16346 14908 16348
rect 14932 16346 14988 16348
rect 15012 16346 15068 16348
rect 15092 16346 15148 16348
rect 14852 16294 14898 16346
rect 14898 16294 14908 16346
rect 14932 16294 14962 16346
rect 14962 16294 14974 16346
rect 14974 16294 14988 16346
rect 15012 16294 15026 16346
rect 15026 16294 15038 16346
rect 15038 16294 15068 16346
rect 15092 16294 15102 16346
rect 15102 16294 15148 16346
rect 14852 16292 14908 16294
rect 14932 16292 14988 16294
rect 15012 16292 15068 16294
rect 15092 16292 15148 16294
rect 21800 16346 21856 16348
rect 21880 16346 21936 16348
rect 21960 16346 22016 16348
rect 22040 16346 22096 16348
rect 21800 16294 21846 16346
rect 21846 16294 21856 16346
rect 21880 16294 21910 16346
rect 21910 16294 21922 16346
rect 21922 16294 21936 16346
rect 21960 16294 21974 16346
rect 21974 16294 21986 16346
rect 21986 16294 22016 16346
rect 22040 16294 22050 16346
rect 22050 16294 22096 16346
rect 21800 16292 21856 16294
rect 21880 16292 21936 16294
rect 21960 16292 22016 16294
rect 22040 16292 22096 16294
rect 4430 15802 4486 15804
rect 4510 15802 4566 15804
rect 4590 15802 4646 15804
rect 4670 15802 4726 15804
rect 4430 15750 4476 15802
rect 4476 15750 4486 15802
rect 4510 15750 4540 15802
rect 4540 15750 4552 15802
rect 4552 15750 4566 15802
rect 4590 15750 4604 15802
rect 4604 15750 4616 15802
rect 4616 15750 4646 15802
rect 4670 15750 4680 15802
rect 4680 15750 4726 15802
rect 4430 15748 4486 15750
rect 4510 15748 4566 15750
rect 4590 15748 4646 15750
rect 4670 15748 4726 15750
rect 11378 15802 11434 15804
rect 11458 15802 11514 15804
rect 11538 15802 11594 15804
rect 11618 15802 11674 15804
rect 11378 15750 11424 15802
rect 11424 15750 11434 15802
rect 11458 15750 11488 15802
rect 11488 15750 11500 15802
rect 11500 15750 11514 15802
rect 11538 15750 11552 15802
rect 11552 15750 11564 15802
rect 11564 15750 11594 15802
rect 11618 15750 11628 15802
rect 11628 15750 11674 15802
rect 11378 15748 11434 15750
rect 11458 15748 11514 15750
rect 11538 15748 11594 15750
rect 11618 15748 11674 15750
rect 18326 15802 18382 15804
rect 18406 15802 18462 15804
rect 18486 15802 18542 15804
rect 18566 15802 18622 15804
rect 18326 15750 18372 15802
rect 18372 15750 18382 15802
rect 18406 15750 18436 15802
rect 18436 15750 18448 15802
rect 18448 15750 18462 15802
rect 18486 15750 18500 15802
rect 18500 15750 18512 15802
rect 18512 15750 18542 15802
rect 18566 15750 18576 15802
rect 18576 15750 18622 15802
rect 18326 15748 18382 15750
rect 18406 15748 18462 15750
rect 18486 15748 18542 15750
rect 18566 15748 18622 15750
rect 25274 15802 25330 15804
rect 25354 15802 25410 15804
rect 25434 15802 25490 15804
rect 25514 15802 25570 15804
rect 25274 15750 25320 15802
rect 25320 15750 25330 15802
rect 25354 15750 25384 15802
rect 25384 15750 25396 15802
rect 25396 15750 25410 15802
rect 25434 15750 25448 15802
rect 25448 15750 25460 15802
rect 25460 15750 25490 15802
rect 25514 15750 25524 15802
rect 25524 15750 25570 15802
rect 25274 15748 25330 15750
rect 25354 15748 25410 15750
rect 25434 15748 25490 15750
rect 25514 15748 25570 15750
rect 7904 15258 7960 15260
rect 7984 15258 8040 15260
rect 8064 15258 8120 15260
rect 8144 15258 8200 15260
rect 7904 15206 7950 15258
rect 7950 15206 7960 15258
rect 7984 15206 8014 15258
rect 8014 15206 8026 15258
rect 8026 15206 8040 15258
rect 8064 15206 8078 15258
rect 8078 15206 8090 15258
rect 8090 15206 8120 15258
rect 8144 15206 8154 15258
rect 8154 15206 8200 15258
rect 7904 15204 7960 15206
rect 7984 15204 8040 15206
rect 8064 15204 8120 15206
rect 8144 15204 8200 15206
rect 14852 15258 14908 15260
rect 14932 15258 14988 15260
rect 15012 15258 15068 15260
rect 15092 15258 15148 15260
rect 14852 15206 14898 15258
rect 14898 15206 14908 15258
rect 14932 15206 14962 15258
rect 14962 15206 14974 15258
rect 14974 15206 14988 15258
rect 15012 15206 15026 15258
rect 15026 15206 15038 15258
rect 15038 15206 15068 15258
rect 15092 15206 15102 15258
rect 15102 15206 15148 15258
rect 14852 15204 14908 15206
rect 14932 15204 14988 15206
rect 15012 15204 15068 15206
rect 15092 15204 15148 15206
rect 21800 15258 21856 15260
rect 21880 15258 21936 15260
rect 21960 15258 22016 15260
rect 22040 15258 22096 15260
rect 21800 15206 21846 15258
rect 21846 15206 21856 15258
rect 21880 15206 21910 15258
rect 21910 15206 21922 15258
rect 21922 15206 21936 15258
rect 21960 15206 21974 15258
rect 21974 15206 21986 15258
rect 21986 15206 22016 15258
rect 22040 15206 22050 15258
rect 22050 15206 22096 15258
rect 21800 15204 21856 15206
rect 21880 15204 21936 15206
rect 21960 15204 22016 15206
rect 22040 15204 22096 15206
rect 4430 14714 4486 14716
rect 4510 14714 4566 14716
rect 4590 14714 4646 14716
rect 4670 14714 4726 14716
rect 4430 14662 4476 14714
rect 4476 14662 4486 14714
rect 4510 14662 4540 14714
rect 4540 14662 4552 14714
rect 4552 14662 4566 14714
rect 4590 14662 4604 14714
rect 4604 14662 4616 14714
rect 4616 14662 4646 14714
rect 4670 14662 4680 14714
rect 4680 14662 4726 14714
rect 4430 14660 4486 14662
rect 4510 14660 4566 14662
rect 4590 14660 4646 14662
rect 4670 14660 4726 14662
rect 11378 14714 11434 14716
rect 11458 14714 11514 14716
rect 11538 14714 11594 14716
rect 11618 14714 11674 14716
rect 11378 14662 11424 14714
rect 11424 14662 11434 14714
rect 11458 14662 11488 14714
rect 11488 14662 11500 14714
rect 11500 14662 11514 14714
rect 11538 14662 11552 14714
rect 11552 14662 11564 14714
rect 11564 14662 11594 14714
rect 11618 14662 11628 14714
rect 11628 14662 11674 14714
rect 11378 14660 11434 14662
rect 11458 14660 11514 14662
rect 11538 14660 11594 14662
rect 11618 14660 11674 14662
rect 18326 14714 18382 14716
rect 18406 14714 18462 14716
rect 18486 14714 18542 14716
rect 18566 14714 18622 14716
rect 18326 14662 18372 14714
rect 18372 14662 18382 14714
rect 18406 14662 18436 14714
rect 18436 14662 18448 14714
rect 18448 14662 18462 14714
rect 18486 14662 18500 14714
rect 18500 14662 18512 14714
rect 18512 14662 18542 14714
rect 18566 14662 18576 14714
rect 18576 14662 18622 14714
rect 18326 14660 18382 14662
rect 18406 14660 18462 14662
rect 18486 14660 18542 14662
rect 18566 14660 18622 14662
rect 25274 14714 25330 14716
rect 25354 14714 25410 14716
rect 25434 14714 25490 14716
rect 25514 14714 25570 14716
rect 25274 14662 25320 14714
rect 25320 14662 25330 14714
rect 25354 14662 25384 14714
rect 25384 14662 25396 14714
rect 25396 14662 25410 14714
rect 25434 14662 25448 14714
rect 25448 14662 25460 14714
rect 25460 14662 25490 14714
rect 25514 14662 25524 14714
rect 25524 14662 25570 14714
rect 25274 14660 25330 14662
rect 25354 14660 25410 14662
rect 25434 14660 25490 14662
rect 25514 14660 25570 14662
rect 7904 14170 7960 14172
rect 7984 14170 8040 14172
rect 8064 14170 8120 14172
rect 8144 14170 8200 14172
rect 7904 14118 7950 14170
rect 7950 14118 7960 14170
rect 7984 14118 8014 14170
rect 8014 14118 8026 14170
rect 8026 14118 8040 14170
rect 8064 14118 8078 14170
rect 8078 14118 8090 14170
rect 8090 14118 8120 14170
rect 8144 14118 8154 14170
rect 8154 14118 8200 14170
rect 7904 14116 7960 14118
rect 7984 14116 8040 14118
rect 8064 14116 8120 14118
rect 8144 14116 8200 14118
rect 14852 14170 14908 14172
rect 14932 14170 14988 14172
rect 15012 14170 15068 14172
rect 15092 14170 15148 14172
rect 14852 14118 14898 14170
rect 14898 14118 14908 14170
rect 14932 14118 14962 14170
rect 14962 14118 14974 14170
rect 14974 14118 14988 14170
rect 15012 14118 15026 14170
rect 15026 14118 15038 14170
rect 15038 14118 15068 14170
rect 15092 14118 15102 14170
rect 15102 14118 15148 14170
rect 14852 14116 14908 14118
rect 14932 14116 14988 14118
rect 15012 14116 15068 14118
rect 15092 14116 15148 14118
rect 21800 14170 21856 14172
rect 21880 14170 21936 14172
rect 21960 14170 22016 14172
rect 22040 14170 22096 14172
rect 21800 14118 21846 14170
rect 21846 14118 21856 14170
rect 21880 14118 21910 14170
rect 21910 14118 21922 14170
rect 21922 14118 21936 14170
rect 21960 14118 21974 14170
rect 21974 14118 21986 14170
rect 21986 14118 22016 14170
rect 22040 14118 22050 14170
rect 22050 14118 22096 14170
rect 21800 14116 21856 14118
rect 21880 14116 21936 14118
rect 21960 14116 22016 14118
rect 22040 14116 22096 14118
rect 28170 13640 28226 13696
rect 4430 13626 4486 13628
rect 4510 13626 4566 13628
rect 4590 13626 4646 13628
rect 4670 13626 4726 13628
rect 4430 13574 4476 13626
rect 4476 13574 4486 13626
rect 4510 13574 4540 13626
rect 4540 13574 4552 13626
rect 4552 13574 4566 13626
rect 4590 13574 4604 13626
rect 4604 13574 4616 13626
rect 4616 13574 4646 13626
rect 4670 13574 4680 13626
rect 4680 13574 4726 13626
rect 4430 13572 4486 13574
rect 4510 13572 4566 13574
rect 4590 13572 4646 13574
rect 4670 13572 4726 13574
rect 11378 13626 11434 13628
rect 11458 13626 11514 13628
rect 11538 13626 11594 13628
rect 11618 13626 11674 13628
rect 11378 13574 11424 13626
rect 11424 13574 11434 13626
rect 11458 13574 11488 13626
rect 11488 13574 11500 13626
rect 11500 13574 11514 13626
rect 11538 13574 11552 13626
rect 11552 13574 11564 13626
rect 11564 13574 11594 13626
rect 11618 13574 11628 13626
rect 11628 13574 11674 13626
rect 11378 13572 11434 13574
rect 11458 13572 11514 13574
rect 11538 13572 11594 13574
rect 11618 13572 11674 13574
rect 18326 13626 18382 13628
rect 18406 13626 18462 13628
rect 18486 13626 18542 13628
rect 18566 13626 18622 13628
rect 18326 13574 18372 13626
rect 18372 13574 18382 13626
rect 18406 13574 18436 13626
rect 18436 13574 18448 13626
rect 18448 13574 18462 13626
rect 18486 13574 18500 13626
rect 18500 13574 18512 13626
rect 18512 13574 18542 13626
rect 18566 13574 18576 13626
rect 18576 13574 18622 13626
rect 18326 13572 18382 13574
rect 18406 13572 18462 13574
rect 18486 13572 18542 13574
rect 18566 13572 18622 13574
rect 25274 13626 25330 13628
rect 25354 13626 25410 13628
rect 25434 13626 25490 13628
rect 25514 13626 25570 13628
rect 25274 13574 25320 13626
rect 25320 13574 25330 13626
rect 25354 13574 25384 13626
rect 25384 13574 25396 13626
rect 25396 13574 25410 13626
rect 25434 13574 25448 13626
rect 25448 13574 25460 13626
rect 25460 13574 25490 13626
rect 25514 13574 25524 13626
rect 25524 13574 25570 13626
rect 25274 13572 25330 13574
rect 25354 13572 25410 13574
rect 25434 13572 25490 13574
rect 25514 13572 25570 13574
rect 7904 13082 7960 13084
rect 7984 13082 8040 13084
rect 8064 13082 8120 13084
rect 8144 13082 8200 13084
rect 7904 13030 7950 13082
rect 7950 13030 7960 13082
rect 7984 13030 8014 13082
rect 8014 13030 8026 13082
rect 8026 13030 8040 13082
rect 8064 13030 8078 13082
rect 8078 13030 8090 13082
rect 8090 13030 8120 13082
rect 8144 13030 8154 13082
rect 8154 13030 8200 13082
rect 7904 13028 7960 13030
rect 7984 13028 8040 13030
rect 8064 13028 8120 13030
rect 8144 13028 8200 13030
rect 14852 13082 14908 13084
rect 14932 13082 14988 13084
rect 15012 13082 15068 13084
rect 15092 13082 15148 13084
rect 14852 13030 14898 13082
rect 14898 13030 14908 13082
rect 14932 13030 14962 13082
rect 14962 13030 14974 13082
rect 14974 13030 14988 13082
rect 15012 13030 15026 13082
rect 15026 13030 15038 13082
rect 15038 13030 15068 13082
rect 15092 13030 15102 13082
rect 15102 13030 15148 13082
rect 14852 13028 14908 13030
rect 14932 13028 14988 13030
rect 15012 13028 15068 13030
rect 15092 13028 15148 13030
rect 21800 13082 21856 13084
rect 21880 13082 21936 13084
rect 21960 13082 22016 13084
rect 22040 13082 22096 13084
rect 21800 13030 21846 13082
rect 21846 13030 21856 13082
rect 21880 13030 21910 13082
rect 21910 13030 21922 13082
rect 21922 13030 21936 13082
rect 21960 13030 21974 13082
rect 21974 13030 21986 13082
rect 21986 13030 22016 13082
rect 22040 13030 22050 13082
rect 22050 13030 22096 13082
rect 21800 13028 21856 13030
rect 21880 13028 21936 13030
rect 21960 13028 22016 13030
rect 22040 13028 22096 13030
rect 4430 12538 4486 12540
rect 4510 12538 4566 12540
rect 4590 12538 4646 12540
rect 4670 12538 4726 12540
rect 4430 12486 4476 12538
rect 4476 12486 4486 12538
rect 4510 12486 4540 12538
rect 4540 12486 4552 12538
rect 4552 12486 4566 12538
rect 4590 12486 4604 12538
rect 4604 12486 4616 12538
rect 4616 12486 4646 12538
rect 4670 12486 4680 12538
rect 4680 12486 4726 12538
rect 4430 12484 4486 12486
rect 4510 12484 4566 12486
rect 4590 12484 4646 12486
rect 4670 12484 4726 12486
rect 11378 12538 11434 12540
rect 11458 12538 11514 12540
rect 11538 12538 11594 12540
rect 11618 12538 11674 12540
rect 11378 12486 11424 12538
rect 11424 12486 11434 12538
rect 11458 12486 11488 12538
rect 11488 12486 11500 12538
rect 11500 12486 11514 12538
rect 11538 12486 11552 12538
rect 11552 12486 11564 12538
rect 11564 12486 11594 12538
rect 11618 12486 11628 12538
rect 11628 12486 11674 12538
rect 11378 12484 11434 12486
rect 11458 12484 11514 12486
rect 11538 12484 11594 12486
rect 11618 12484 11674 12486
rect 18326 12538 18382 12540
rect 18406 12538 18462 12540
rect 18486 12538 18542 12540
rect 18566 12538 18622 12540
rect 18326 12486 18372 12538
rect 18372 12486 18382 12538
rect 18406 12486 18436 12538
rect 18436 12486 18448 12538
rect 18448 12486 18462 12538
rect 18486 12486 18500 12538
rect 18500 12486 18512 12538
rect 18512 12486 18542 12538
rect 18566 12486 18576 12538
rect 18576 12486 18622 12538
rect 18326 12484 18382 12486
rect 18406 12484 18462 12486
rect 18486 12484 18542 12486
rect 18566 12484 18622 12486
rect 25274 12538 25330 12540
rect 25354 12538 25410 12540
rect 25434 12538 25490 12540
rect 25514 12538 25570 12540
rect 25274 12486 25320 12538
rect 25320 12486 25330 12538
rect 25354 12486 25384 12538
rect 25384 12486 25396 12538
rect 25396 12486 25410 12538
rect 25434 12486 25448 12538
rect 25448 12486 25460 12538
rect 25460 12486 25490 12538
rect 25514 12486 25524 12538
rect 25524 12486 25570 12538
rect 25274 12484 25330 12486
rect 25354 12484 25410 12486
rect 25434 12484 25490 12486
rect 25514 12484 25570 12486
rect 7904 11994 7960 11996
rect 7984 11994 8040 11996
rect 8064 11994 8120 11996
rect 8144 11994 8200 11996
rect 7904 11942 7950 11994
rect 7950 11942 7960 11994
rect 7984 11942 8014 11994
rect 8014 11942 8026 11994
rect 8026 11942 8040 11994
rect 8064 11942 8078 11994
rect 8078 11942 8090 11994
rect 8090 11942 8120 11994
rect 8144 11942 8154 11994
rect 8154 11942 8200 11994
rect 7904 11940 7960 11942
rect 7984 11940 8040 11942
rect 8064 11940 8120 11942
rect 8144 11940 8200 11942
rect 14852 11994 14908 11996
rect 14932 11994 14988 11996
rect 15012 11994 15068 11996
rect 15092 11994 15148 11996
rect 14852 11942 14898 11994
rect 14898 11942 14908 11994
rect 14932 11942 14962 11994
rect 14962 11942 14974 11994
rect 14974 11942 14988 11994
rect 15012 11942 15026 11994
rect 15026 11942 15038 11994
rect 15038 11942 15068 11994
rect 15092 11942 15102 11994
rect 15102 11942 15148 11994
rect 14852 11940 14908 11942
rect 14932 11940 14988 11942
rect 15012 11940 15068 11942
rect 15092 11940 15148 11942
rect 21800 11994 21856 11996
rect 21880 11994 21936 11996
rect 21960 11994 22016 11996
rect 22040 11994 22096 11996
rect 21800 11942 21846 11994
rect 21846 11942 21856 11994
rect 21880 11942 21910 11994
rect 21910 11942 21922 11994
rect 21922 11942 21936 11994
rect 21960 11942 21974 11994
rect 21974 11942 21986 11994
rect 21986 11942 22016 11994
rect 22040 11942 22050 11994
rect 22050 11942 22096 11994
rect 21800 11940 21856 11942
rect 21880 11940 21936 11942
rect 21960 11940 22016 11942
rect 22040 11940 22096 11942
rect 4430 11450 4486 11452
rect 4510 11450 4566 11452
rect 4590 11450 4646 11452
rect 4670 11450 4726 11452
rect 4430 11398 4476 11450
rect 4476 11398 4486 11450
rect 4510 11398 4540 11450
rect 4540 11398 4552 11450
rect 4552 11398 4566 11450
rect 4590 11398 4604 11450
rect 4604 11398 4616 11450
rect 4616 11398 4646 11450
rect 4670 11398 4680 11450
rect 4680 11398 4726 11450
rect 4430 11396 4486 11398
rect 4510 11396 4566 11398
rect 4590 11396 4646 11398
rect 4670 11396 4726 11398
rect 11378 11450 11434 11452
rect 11458 11450 11514 11452
rect 11538 11450 11594 11452
rect 11618 11450 11674 11452
rect 11378 11398 11424 11450
rect 11424 11398 11434 11450
rect 11458 11398 11488 11450
rect 11488 11398 11500 11450
rect 11500 11398 11514 11450
rect 11538 11398 11552 11450
rect 11552 11398 11564 11450
rect 11564 11398 11594 11450
rect 11618 11398 11628 11450
rect 11628 11398 11674 11450
rect 11378 11396 11434 11398
rect 11458 11396 11514 11398
rect 11538 11396 11594 11398
rect 11618 11396 11674 11398
rect 18326 11450 18382 11452
rect 18406 11450 18462 11452
rect 18486 11450 18542 11452
rect 18566 11450 18622 11452
rect 18326 11398 18372 11450
rect 18372 11398 18382 11450
rect 18406 11398 18436 11450
rect 18436 11398 18448 11450
rect 18448 11398 18462 11450
rect 18486 11398 18500 11450
rect 18500 11398 18512 11450
rect 18512 11398 18542 11450
rect 18566 11398 18576 11450
rect 18576 11398 18622 11450
rect 18326 11396 18382 11398
rect 18406 11396 18462 11398
rect 18486 11396 18542 11398
rect 18566 11396 18622 11398
rect 25274 11450 25330 11452
rect 25354 11450 25410 11452
rect 25434 11450 25490 11452
rect 25514 11450 25570 11452
rect 25274 11398 25320 11450
rect 25320 11398 25330 11450
rect 25354 11398 25384 11450
rect 25384 11398 25396 11450
rect 25396 11398 25410 11450
rect 25434 11398 25448 11450
rect 25448 11398 25460 11450
rect 25460 11398 25490 11450
rect 25514 11398 25524 11450
rect 25524 11398 25570 11450
rect 25274 11396 25330 11398
rect 25354 11396 25410 11398
rect 25434 11396 25490 11398
rect 25514 11396 25570 11398
rect 7904 10906 7960 10908
rect 7984 10906 8040 10908
rect 8064 10906 8120 10908
rect 8144 10906 8200 10908
rect 7904 10854 7950 10906
rect 7950 10854 7960 10906
rect 7984 10854 8014 10906
rect 8014 10854 8026 10906
rect 8026 10854 8040 10906
rect 8064 10854 8078 10906
rect 8078 10854 8090 10906
rect 8090 10854 8120 10906
rect 8144 10854 8154 10906
rect 8154 10854 8200 10906
rect 7904 10852 7960 10854
rect 7984 10852 8040 10854
rect 8064 10852 8120 10854
rect 8144 10852 8200 10854
rect 14852 10906 14908 10908
rect 14932 10906 14988 10908
rect 15012 10906 15068 10908
rect 15092 10906 15148 10908
rect 14852 10854 14898 10906
rect 14898 10854 14908 10906
rect 14932 10854 14962 10906
rect 14962 10854 14974 10906
rect 14974 10854 14988 10906
rect 15012 10854 15026 10906
rect 15026 10854 15038 10906
rect 15038 10854 15068 10906
rect 15092 10854 15102 10906
rect 15102 10854 15148 10906
rect 14852 10852 14908 10854
rect 14932 10852 14988 10854
rect 15012 10852 15068 10854
rect 15092 10852 15148 10854
rect 21800 10906 21856 10908
rect 21880 10906 21936 10908
rect 21960 10906 22016 10908
rect 22040 10906 22096 10908
rect 21800 10854 21846 10906
rect 21846 10854 21856 10906
rect 21880 10854 21910 10906
rect 21910 10854 21922 10906
rect 21922 10854 21936 10906
rect 21960 10854 21974 10906
rect 21974 10854 21986 10906
rect 21986 10854 22016 10906
rect 22040 10854 22050 10906
rect 22050 10854 22096 10906
rect 21800 10852 21856 10854
rect 21880 10852 21936 10854
rect 21960 10852 22016 10854
rect 22040 10852 22096 10854
rect 4430 10362 4486 10364
rect 4510 10362 4566 10364
rect 4590 10362 4646 10364
rect 4670 10362 4726 10364
rect 4430 10310 4476 10362
rect 4476 10310 4486 10362
rect 4510 10310 4540 10362
rect 4540 10310 4552 10362
rect 4552 10310 4566 10362
rect 4590 10310 4604 10362
rect 4604 10310 4616 10362
rect 4616 10310 4646 10362
rect 4670 10310 4680 10362
rect 4680 10310 4726 10362
rect 4430 10308 4486 10310
rect 4510 10308 4566 10310
rect 4590 10308 4646 10310
rect 4670 10308 4726 10310
rect 11378 10362 11434 10364
rect 11458 10362 11514 10364
rect 11538 10362 11594 10364
rect 11618 10362 11674 10364
rect 11378 10310 11424 10362
rect 11424 10310 11434 10362
rect 11458 10310 11488 10362
rect 11488 10310 11500 10362
rect 11500 10310 11514 10362
rect 11538 10310 11552 10362
rect 11552 10310 11564 10362
rect 11564 10310 11594 10362
rect 11618 10310 11628 10362
rect 11628 10310 11674 10362
rect 11378 10308 11434 10310
rect 11458 10308 11514 10310
rect 11538 10308 11594 10310
rect 11618 10308 11674 10310
rect 18326 10362 18382 10364
rect 18406 10362 18462 10364
rect 18486 10362 18542 10364
rect 18566 10362 18622 10364
rect 18326 10310 18372 10362
rect 18372 10310 18382 10362
rect 18406 10310 18436 10362
rect 18436 10310 18448 10362
rect 18448 10310 18462 10362
rect 18486 10310 18500 10362
rect 18500 10310 18512 10362
rect 18512 10310 18542 10362
rect 18566 10310 18576 10362
rect 18576 10310 18622 10362
rect 18326 10308 18382 10310
rect 18406 10308 18462 10310
rect 18486 10308 18542 10310
rect 18566 10308 18622 10310
rect 25274 10362 25330 10364
rect 25354 10362 25410 10364
rect 25434 10362 25490 10364
rect 25514 10362 25570 10364
rect 25274 10310 25320 10362
rect 25320 10310 25330 10362
rect 25354 10310 25384 10362
rect 25384 10310 25396 10362
rect 25396 10310 25410 10362
rect 25434 10310 25448 10362
rect 25448 10310 25460 10362
rect 25460 10310 25490 10362
rect 25514 10310 25524 10362
rect 25524 10310 25570 10362
rect 25274 10308 25330 10310
rect 25354 10308 25410 10310
rect 25434 10308 25490 10310
rect 25514 10308 25570 10310
rect 7904 9818 7960 9820
rect 7984 9818 8040 9820
rect 8064 9818 8120 9820
rect 8144 9818 8200 9820
rect 7904 9766 7950 9818
rect 7950 9766 7960 9818
rect 7984 9766 8014 9818
rect 8014 9766 8026 9818
rect 8026 9766 8040 9818
rect 8064 9766 8078 9818
rect 8078 9766 8090 9818
rect 8090 9766 8120 9818
rect 8144 9766 8154 9818
rect 8154 9766 8200 9818
rect 7904 9764 7960 9766
rect 7984 9764 8040 9766
rect 8064 9764 8120 9766
rect 8144 9764 8200 9766
rect 4430 9274 4486 9276
rect 4510 9274 4566 9276
rect 4590 9274 4646 9276
rect 4670 9274 4726 9276
rect 4430 9222 4476 9274
rect 4476 9222 4486 9274
rect 4510 9222 4540 9274
rect 4540 9222 4552 9274
rect 4552 9222 4566 9274
rect 4590 9222 4604 9274
rect 4604 9222 4616 9274
rect 4616 9222 4646 9274
rect 4670 9222 4680 9274
rect 4680 9222 4726 9274
rect 4430 9220 4486 9222
rect 4510 9220 4566 9222
rect 4590 9220 4646 9222
rect 4670 9220 4726 9222
rect 11378 9274 11434 9276
rect 11458 9274 11514 9276
rect 11538 9274 11594 9276
rect 11618 9274 11674 9276
rect 11378 9222 11424 9274
rect 11424 9222 11434 9274
rect 11458 9222 11488 9274
rect 11488 9222 11500 9274
rect 11500 9222 11514 9274
rect 11538 9222 11552 9274
rect 11552 9222 11564 9274
rect 11564 9222 11594 9274
rect 11618 9222 11628 9274
rect 11628 9222 11674 9274
rect 11378 9220 11434 9222
rect 11458 9220 11514 9222
rect 11538 9220 11594 9222
rect 11618 9220 11674 9222
rect 7904 8730 7960 8732
rect 7984 8730 8040 8732
rect 8064 8730 8120 8732
rect 8144 8730 8200 8732
rect 7904 8678 7950 8730
rect 7950 8678 7960 8730
rect 7984 8678 8014 8730
rect 8014 8678 8026 8730
rect 8026 8678 8040 8730
rect 8064 8678 8078 8730
rect 8078 8678 8090 8730
rect 8090 8678 8120 8730
rect 8144 8678 8154 8730
rect 8154 8678 8200 8730
rect 7904 8676 7960 8678
rect 7984 8676 8040 8678
rect 8064 8676 8120 8678
rect 8144 8676 8200 8678
rect 4430 8186 4486 8188
rect 4510 8186 4566 8188
rect 4590 8186 4646 8188
rect 4670 8186 4726 8188
rect 4430 8134 4476 8186
rect 4476 8134 4486 8186
rect 4510 8134 4540 8186
rect 4540 8134 4552 8186
rect 4552 8134 4566 8186
rect 4590 8134 4604 8186
rect 4604 8134 4616 8186
rect 4616 8134 4646 8186
rect 4670 8134 4680 8186
rect 4680 8134 4726 8186
rect 4430 8132 4486 8134
rect 4510 8132 4566 8134
rect 4590 8132 4646 8134
rect 4670 8132 4726 8134
rect 11378 8186 11434 8188
rect 11458 8186 11514 8188
rect 11538 8186 11594 8188
rect 11618 8186 11674 8188
rect 11378 8134 11424 8186
rect 11424 8134 11434 8186
rect 11458 8134 11488 8186
rect 11488 8134 11500 8186
rect 11500 8134 11514 8186
rect 11538 8134 11552 8186
rect 11552 8134 11564 8186
rect 11564 8134 11594 8186
rect 11618 8134 11628 8186
rect 11628 8134 11674 8186
rect 11378 8132 11434 8134
rect 11458 8132 11514 8134
rect 11538 8132 11594 8134
rect 11618 8132 11674 8134
rect 7904 7642 7960 7644
rect 7984 7642 8040 7644
rect 8064 7642 8120 7644
rect 8144 7642 8200 7644
rect 7904 7590 7950 7642
rect 7950 7590 7960 7642
rect 7984 7590 8014 7642
rect 8014 7590 8026 7642
rect 8026 7590 8040 7642
rect 8064 7590 8078 7642
rect 8078 7590 8090 7642
rect 8090 7590 8120 7642
rect 8144 7590 8154 7642
rect 8154 7590 8200 7642
rect 7904 7588 7960 7590
rect 7984 7588 8040 7590
rect 8064 7588 8120 7590
rect 8144 7588 8200 7590
rect 14852 9818 14908 9820
rect 14932 9818 14988 9820
rect 15012 9818 15068 9820
rect 15092 9818 15148 9820
rect 14852 9766 14898 9818
rect 14898 9766 14908 9818
rect 14932 9766 14962 9818
rect 14962 9766 14974 9818
rect 14974 9766 14988 9818
rect 15012 9766 15026 9818
rect 15026 9766 15038 9818
rect 15038 9766 15068 9818
rect 15092 9766 15102 9818
rect 15102 9766 15148 9818
rect 14852 9764 14908 9766
rect 14932 9764 14988 9766
rect 15012 9764 15068 9766
rect 15092 9764 15148 9766
rect 21800 9818 21856 9820
rect 21880 9818 21936 9820
rect 21960 9818 22016 9820
rect 22040 9818 22096 9820
rect 21800 9766 21846 9818
rect 21846 9766 21856 9818
rect 21880 9766 21910 9818
rect 21910 9766 21922 9818
rect 21922 9766 21936 9818
rect 21960 9766 21974 9818
rect 21974 9766 21986 9818
rect 21986 9766 22016 9818
rect 22040 9766 22050 9818
rect 22050 9766 22096 9818
rect 21800 9764 21856 9766
rect 21880 9764 21936 9766
rect 21960 9764 22016 9766
rect 22040 9764 22096 9766
rect 27526 9560 27582 9616
rect 18326 9274 18382 9276
rect 18406 9274 18462 9276
rect 18486 9274 18542 9276
rect 18566 9274 18622 9276
rect 18326 9222 18372 9274
rect 18372 9222 18382 9274
rect 18406 9222 18436 9274
rect 18436 9222 18448 9274
rect 18448 9222 18462 9274
rect 18486 9222 18500 9274
rect 18500 9222 18512 9274
rect 18512 9222 18542 9274
rect 18566 9222 18576 9274
rect 18576 9222 18622 9274
rect 18326 9220 18382 9222
rect 18406 9220 18462 9222
rect 18486 9220 18542 9222
rect 18566 9220 18622 9222
rect 25274 9274 25330 9276
rect 25354 9274 25410 9276
rect 25434 9274 25490 9276
rect 25514 9274 25570 9276
rect 25274 9222 25320 9274
rect 25320 9222 25330 9274
rect 25354 9222 25384 9274
rect 25384 9222 25396 9274
rect 25396 9222 25410 9274
rect 25434 9222 25448 9274
rect 25448 9222 25460 9274
rect 25460 9222 25490 9274
rect 25514 9222 25524 9274
rect 25524 9222 25570 9274
rect 25274 9220 25330 9222
rect 25354 9220 25410 9222
rect 25434 9220 25490 9222
rect 25514 9220 25570 9222
rect 14852 8730 14908 8732
rect 14932 8730 14988 8732
rect 15012 8730 15068 8732
rect 15092 8730 15148 8732
rect 14852 8678 14898 8730
rect 14898 8678 14908 8730
rect 14932 8678 14962 8730
rect 14962 8678 14974 8730
rect 14974 8678 14988 8730
rect 15012 8678 15026 8730
rect 15026 8678 15038 8730
rect 15038 8678 15068 8730
rect 15092 8678 15102 8730
rect 15102 8678 15148 8730
rect 14852 8676 14908 8678
rect 14932 8676 14988 8678
rect 15012 8676 15068 8678
rect 15092 8676 15148 8678
rect 21800 8730 21856 8732
rect 21880 8730 21936 8732
rect 21960 8730 22016 8732
rect 22040 8730 22096 8732
rect 21800 8678 21846 8730
rect 21846 8678 21856 8730
rect 21880 8678 21910 8730
rect 21910 8678 21922 8730
rect 21922 8678 21936 8730
rect 21960 8678 21974 8730
rect 21974 8678 21986 8730
rect 21986 8678 22016 8730
rect 22040 8678 22050 8730
rect 22050 8678 22096 8730
rect 21800 8676 21856 8678
rect 21880 8676 21936 8678
rect 21960 8676 22016 8678
rect 22040 8676 22096 8678
rect 18326 8186 18382 8188
rect 18406 8186 18462 8188
rect 18486 8186 18542 8188
rect 18566 8186 18622 8188
rect 18326 8134 18372 8186
rect 18372 8134 18382 8186
rect 18406 8134 18436 8186
rect 18436 8134 18448 8186
rect 18448 8134 18462 8186
rect 18486 8134 18500 8186
rect 18500 8134 18512 8186
rect 18512 8134 18542 8186
rect 18566 8134 18576 8186
rect 18576 8134 18622 8186
rect 18326 8132 18382 8134
rect 18406 8132 18462 8134
rect 18486 8132 18542 8134
rect 18566 8132 18622 8134
rect 25274 8186 25330 8188
rect 25354 8186 25410 8188
rect 25434 8186 25490 8188
rect 25514 8186 25570 8188
rect 25274 8134 25320 8186
rect 25320 8134 25330 8186
rect 25354 8134 25384 8186
rect 25384 8134 25396 8186
rect 25396 8134 25410 8186
rect 25434 8134 25448 8186
rect 25448 8134 25460 8186
rect 25460 8134 25490 8186
rect 25514 8134 25524 8186
rect 25524 8134 25570 8186
rect 25274 8132 25330 8134
rect 25354 8132 25410 8134
rect 25434 8132 25490 8134
rect 25514 8132 25570 8134
rect 14852 7642 14908 7644
rect 14932 7642 14988 7644
rect 15012 7642 15068 7644
rect 15092 7642 15148 7644
rect 14852 7590 14898 7642
rect 14898 7590 14908 7642
rect 14932 7590 14962 7642
rect 14962 7590 14974 7642
rect 14974 7590 14988 7642
rect 15012 7590 15026 7642
rect 15026 7590 15038 7642
rect 15038 7590 15068 7642
rect 15092 7590 15102 7642
rect 15102 7590 15148 7642
rect 14852 7588 14908 7590
rect 14932 7588 14988 7590
rect 15012 7588 15068 7590
rect 15092 7588 15148 7590
rect 21800 7642 21856 7644
rect 21880 7642 21936 7644
rect 21960 7642 22016 7644
rect 22040 7642 22096 7644
rect 21800 7590 21846 7642
rect 21846 7590 21856 7642
rect 21880 7590 21910 7642
rect 21910 7590 21922 7642
rect 21922 7590 21936 7642
rect 21960 7590 21974 7642
rect 21974 7590 21986 7642
rect 21986 7590 22016 7642
rect 22040 7590 22050 7642
rect 22050 7590 22096 7642
rect 21800 7588 21856 7590
rect 21880 7588 21936 7590
rect 21960 7588 22016 7590
rect 22040 7588 22096 7590
rect 4430 7098 4486 7100
rect 4510 7098 4566 7100
rect 4590 7098 4646 7100
rect 4670 7098 4726 7100
rect 4430 7046 4476 7098
rect 4476 7046 4486 7098
rect 4510 7046 4540 7098
rect 4540 7046 4552 7098
rect 4552 7046 4566 7098
rect 4590 7046 4604 7098
rect 4604 7046 4616 7098
rect 4616 7046 4646 7098
rect 4670 7046 4680 7098
rect 4680 7046 4726 7098
rect 4430 7044 4486 7046
rect 4510 7044 4566 7046
rect 4590 7044 4646 7046
rect 4670 7044 4726 7046
rect 4430 6010 4486 6012
rect 4510 6010 4566 6012
rect 4590 6010 4646 6012
rect 4670 6010 4726 6012
rect 4430 5958 4476 6010
rect 4476 5958 4486 6010
rect 4510 5958 4540 6010
rect 4540 5958 4552 6010
rect 4552 5958 4566 6010
rect 4590 5958 4604 6010
rect 4604 5958 4616 6010
rect 4616 5958 4646 6010
rect 4670 5958 4680 6010
rect 4680 5958 4726 6010
rect 4430 5956 4486 5958
rect 4510 5956 4566 5958
rect 4590 5956 4646 5958
rect 4670 5956 4726 5958
rect 4430 4922 4486 4924
rect 4510 4922 4566 4924
rect 4590 4922 4646 4924
rect 4670 4922 4726 4924
rect 4430 4870 4476 4922
rect 4476 4870 4486 4922
rect 4510 4870 4540 4922
rect 4540 4870 4552 4922
rect 4552 4870 4566 4922
rect 4590 4870 4604 4922
rect 4604 4870 4616 4922
rect 4616 4870 4646 4922
rect 4670 4870 4680 4922
rect 4680 4870 4726 4922
rect 4430 4868 4486 4870
rect 4510 4868 4566 4870
rect 4590 4868 4646 4870
rect 4670 4868 4726 4870
rect 4430 3834 4486 3836
rect 4510 3834 4566 3836
rect 4590 3834 4646 3836
rect 4670 3834 4726 3836
rect 4430 3782 4476 3834
rect 4476 3782 4486 3834
rect 4510 3782 4540 3834
rect 4540 3782 4552 3834
rect 4552 3782 4566 3834
rect 4590 3782 4604 3834
rect 4604 3782 4616 3834
rect 4616 3782 4646 3834
rect 4670 3782 4680 3834
rect 4680 3782 4726 3834
rect 4430 3780 4486 3782
rect 4510 3780 4566 3782
rect 4590 3780 4646 3782
rect 4670 3780 4726 3782
rect 4430 2746 4486 2748
rect 4510 2746 4566 2748
rect 4590 2746 4646 2748
rect 4670 2746 4726 2748
rect 4430 2694 4476 2746
rect 4476 2694 4486 2746
rect 4510 2694 4540 2746
rect 4540 2694 4552 2746
rect 4552 2694 4566 2746
rect 4590 2694 4604 2746
rect 4604 2694 4616 2746
rect 4616 2694 4646 2746
rect 4670 2694 4680 2746
rect 4680 2694 4726 2746
rect 4430 2692 4486 2694
rect 4510 2692 4566 2694
rect 4590 2692 4646 2694
rect 4670 2692 4726 2694
rect 11378 7098 11434 7100
rect 11458 7098 11514 7100
rect 11538 7098 11594 7100
rect 11618 7098 11674 7100
rect 11378 7046 11424 7098
rect 11424 7046 11434 7098
rect 11458 7046 11488 7098
rect 11488 7046 11500 7098
rect 11500 7046 11514 7098
rect 11538 7046 11552 7098
rect 11552 7046 11564 7098
rect 11564 7046 11594 7098
rect 11618 7046 11628 7098
rect 11628 7046 11674 7098
rect 11378 7044 11434 7046
rect 11458 7044 11514 7046
rect 11538 7044 11594 7046
rect 11618 7044 11674 7046
rect 18326 7098 18382 7100
rect 18406 7098 18462 7100
rect 18486 7098 18542 7100
rect 18566 7098 18622 7100
rect 18326 7046 18372 7098
rect 18372 7046 18382 7098
rect 18406 7046 18436 7098
rect 18436 7046 18448 7098
rect 18448 7046 18462 7098
rect 18486 7046 18500 7098
rect 18500 7046 18512 7098
rect 18512 7046 18542 7098
rect 18566 7046 18576 7098
rect 18576 7046 18622 7098
rect 18326 7044 18382 7046
rect 18406 7044 18462 7046
rect 18486 7044 18542 7046
rect 18566 7044 18622 7046
rect 25274 7098 25330 7100
rect 25354 7098 25410 7100
rect 25434 7098 25490 7100
rect 25514 7098 25570 7100
rect 25274 7046 25320 7098
rect 25320 7046 25330 7098
rect 25354 7046 25384 7098
rect 25384 7046 25396 7098
rect 25396 7046 25410 7098
rect 25434 7046 25448 7098
rect 25448 7046 25460 7098
rect 25460 7046 25490 7098
rect 25514 7046 25524 7098
rect 25524 7046 25570 7098
rect 25274 7044 25330 7046
rect 25354 7044 25410 7046
rect 25434 7044 25490 7046
rect 25514 7044 25570 7046
rect 7904 6554 7960 6556
rect 7984 6554 8040 6556
rect 8064 6554 8120 6556
rect 8144 6554 8200 6556
rect 7904 6502 7950 6554
rect 7950 6502 7960 6554
rect 7984 6502 8014 6554
rect 8014 6502 8026 6554
rect 8026 6502 8040 6554
rect 8064 6502 8078 6554
rect 8078 6502 8090 6554
rect 8090 6502 8120 6554
rect 8144 6502 8154 6554
rect 8154 6502 8200 6554
rect 7904 6500 7960 6502
rect 7984 6500 8040 6502
rect 8064 6500 8120 6502
rect 8144 6500 8200 6502
rect 14852 6554 14908 6556
rect 14932 6554 14988 6556
rect 15012 6554 15068 6556
rect 15092 6554 15148 6556
rect 14852 6502 14898 6554
rect 14898 6502 14908 6554
rect 14932 6502 14962 6554
rect 14962 6502 14974 6554
rect 14974 6502 14988 6554
rect 15012 6502 15026 6554
rect 15026 6502 15038 6554
rect 15038 6502 15068 6554
rect 15092 6502 15102 6554
rect 15102 6502 15148 6554
rect 14852 6500 14908 6502
rect 14932 6500 14988 6502
rect 15012 6500 15068 6502
rect 15092 6500 15148 6502
rect 21800 6554 21856 6556
rect 21880 6554 21936 6556
rect 21960 6554 22016 6556
rect 22040 6554 22096 6556
rect 21800 6502 21846 6554
rect 21846 6502 21856 6554
rect 21880 6502 21910 6554
rect 21910 6502 21922 6554
rect 21922 6502 21936 6554
rect 21960 6502 21974 6554
rect 21974 6502 21986 6554
rect 21986 6502 22016 6554
rect 22040 6502 22050 6554
rect 22050 6502 22096 6554
rect 21800 6500 21856 6502
rect 21880 6500 21936 6502
rect 21960 6500 22016 6502
rect 22040 6500 22096 6502
rect 11378 6010 11434 6012
rect 11458 6010 11514 6012
rect 11538 6010 11594 6012
rect 11618 6010 11674 6012
rect 11378 5958 11424 6010
rect 11424 5958 11434 6010
rect 11458 5958 11488 6010
rect 11488 5958 11500 6010
rect 11500 5958 11514 6010
rect 11538 5958 11552 6010
rect 11552 5958 11564 6010
rect 11564 5958 11594 6010
rect 11618 5958 11628 6010
rect 11628 5958 11674 6010
rect 11378 5956 11434 5958
rect 11458 5956 11514 5958
rect 11538 5956 11594 5958
rect 11618 5956 11674 5958
rect 18326 6010 18382 6012
rect 18406 6010 18462 6012
rect 18486 6010 18542 6012
rect 18566 6010 18622 6012
rect 18326 5958 18372 6010
rect 18372 5958 18382 6010
rect 18406 5958 18436 6010
rect 18436 5958 18448 6010
rect 18448 5958 18462 6010
rect 18486 5958 18500 6010
rect 18500 5958 18512 6010
rect 18512 5958 18542 6010
rect 18566 5958 18576 6010
rect 18576 5958 18622 6010
rect 18326 5956 18382 5958
rect 18406 5956 18462 5958
rect 18486 5956 18542 5958
rect 18566 5956 18622 5958
rect 25274 6010 25330 6012
rect 25354 6010 25410 6012
rect 25434 6010 25490 6012
rect 25514 6010 25570 6012
rect 25274 5958 25320 6010
rect 25320 5958 25330 6010
rect 25354 5958 25384 6010
rect 25384 5958 25396 6010
rect 25396 5958 25410 6010
rect 25434 5958 25448 6010
rect 25448 5958 25460 6010
rect 25460 5958 25490 6010
rect 25514 5958 25524 6010
rect 25524 5958 25570 6010
rect 25274 5956 25330 5958
rect 25354 5956 25410 5958
rect 25434 5956 25490 5958
rect 25514 5956 25570 5958
rect 7904 5466 7960 5468
rect 7984 5466 8040 5468
rect 8064 5466 8120 5468
rect 8144 5466 8200 5468
rect 7904 5414 7950 5466
rect 7950 5414 7960 5466
rect 7984 5414 8014 5466
rect 8014 5414 8026 5466
rect 8026 5414 8040 5466
rect 8064 5414 8078 5466
rect 8078 5414 8090 5466
rect 8090 5414 8120 5466
rect 8144 5414 8154 5466
rect 8154 5414 8200 5466
rect 7904 5412 7960 5414
rect 7984 5412 8040 5414
rect 8064 5412 8120 5414
rect 8144 5412 8200 5414
rect 14852 5466 14908 5468
rect 14932 5466 14988 5468
rect 15012 5466 15068 5468
rect 15092 5466 15148 5468
rect 14852 5414 14898 5466
rect 14898 5414 14908 5466
rect 14932 5414 14962 5466
rect 14962 5414 14974 5466
rect 14974 5414 14988 5466
rect 15012 5414 15026 5466
rect 15026 5414 15038 5466
rect 15038 5414 15068 5466
rect 15092 5414 15102 5466
rect 15102 5414 15148 5466
rect 14852 5412 14908 5414
rect 14932 5412 14988 5414
rect 15012 5412 15068 5414
rect 15092 5412 15148 5414
rect 21800 5466 21856 5468
rect 21880 5466 21936 5468
rect 21960 5466 22016 5468
rect 22040 5466 22096 5468
rect 21800 5414 21846 5466
rect 21846 5414 21856 5466
rect 21880 5414 21910 5466
rect 21910 5414 21922 5466
rect 21922 5414 21936 5466
rect 21960 5414 21974 5466
rect 21974 5414 21986 5466
rect 21986 5414 22016 5466
rect 22040 5414 22050 5466
rect 22050 5414 22096 5466
rect 21800 5412 21856 5414
rect 21880 5412 21936 5414
rect 21960 5412 22016 5414
rect 22040 5412 22096 5414
rect 11378 4922 11434 4924
rect 11458 4922 11514 4924
rect 11538 4922 11594 4924
rect 11618 4922 11674 4924
rect 11378 4870 11424 4922
rect 11424 4870 11434 4922
rect 11458 4870 11488 4922
rect 11488 4870 11500 4922
rect 11500 4870 11514 4922
rect 11538 4870 11552 4922
rect 11552 4870 11564 4922
rect 11564 4870 11594 4922
rect 11618 4870 11628 4922
rect 11628 4870 11674 4922
rect 11378 4868 11434 4870
rect 11458 4868 11514 4870
rect 11538 4868 11594 4870
rect 11618 4868 11674 4870
rect 18326 4922 18382 4924
rect 18406 4922 18462 4924
rect 18486 4922 18542 4924
rect 18566 4922 18622 4924
rect 18326 4870 18372 4922
rect 18372 4870 18382 4922
rect 18406 4870 18436 4922
rect 18436 4870 18448 4922
rect 18448 4870 18462 4922
rect 18486 4870 18500 4922
rect 18500 4870 18512 4922
rect 18512 4870 18542 4922
rect 18566 4870 18576 4922
rect 18576 4870 18622 4922
rect 18326 4868 18382 4870
rect 18406 4868 18462 4870
rect 18486 4868 18542 4870
rect 18566 4868 18622 4870
rect 25274 4922 25330 4924
rect 25354 4922 25410 4924
rect 25434 4922 25490 4924
rect 25514 4922 25570 4924
rect 25274 4870 25320 4922
rect 25320 4870 25330 4922
rect 25354 4870 25384 4922
rect 25384 4870 25396 4922
rect 25396 4870 25410 4922
rect 25434 4870 25448 4922
rect 25448 4870 25460 4922
rect 25460 4870 25490 4922
rect 25514 4870 25524 4922
rect 25524 4870 25570 4922
rect 25274 4868 25330 4870
rect 25354 4868 25410 4870
rect 25434 4868 25490 4870
rect 25514 4868 25570 4870
rect 7904 4378 7960 4380
rect 7984 4378 8040 4380
rect 8064 4378 8120 4380
rect 8144 4378 8200 4380
rect 7904 4326 7950 4378
rect 7950 4326 7960 4378
rect 7984 4326 8014 4378
rect 8014 4326 8026 4378
rect 8026 4326 8040 4378
rect 8064 4326 8078 4378
rect 8078 4326 8090 4378
rect 8090 4326 8120 4378
rect 8144 4326 8154 4378
rect 8154 4326 8200 4378
rect 7904 4324 7960 4326
rect 7984 4324 8040 4326
rect 8064 4324 8120 4326
rect 8144 4324 8200 4326
rect 14852 4378 14908 4380
rect 14932 4378 14988 4380
rect 15012 4378 15068 4380
rect 15092 4378 15148 4380
rect 14852 4326 14898 4378
rect 14898 4326 14908 4378
rect 14932 4326 14962 4378
rect 14962 4326 14974 4378
rect 14974 4326 14988 4378
rect 15012 4326 15026 4378
rect 15026 4326 15038 4378
rect 15038 4326 15068 4378
rect 15092 4326 15102 4378
rect 15102 4326 15148 4378
rect 14852 4324 14908 4326
rect 14932 4324 14988 4326
rect 15012 4324 15068 4326
rect 15092 4324 15148 4326
rect 21800 4378 21856 4380
rect 21880 4378 21936 4380
rect 21960 4378 22016 4380
rect 22040 4378 22096 4380
rect 21800 4326 21846 4378
rect 21846 4326 21856 4378
rect 21880 4326 21910 4378
rect 21910 4326 21922 4378
rect 21922 4326 21936 4378
rect 21960 4326 21974 4378
rect 21974 4326 21986 4378
rect 21986 4326 22016 4378
rect 22040 4326 22050 4378
rect 22050 4326 22096 4378
rect 21800 4324 21856 4326
rect 21880 4324 21936 4326
rect 21960 4324 22016 4326
rect 22040 4324 22096 4326
rect 11378 3834 11434 3836
rect 11458 3834 11514 3836
rect 11538 3834 11594 3836
rect 11618 3834 11674 3836
rect 11378 3782 11424 3834
rect 11424 3782 11434 3834
rect 11458 3782 11488 3834
rect 11488 3782 11500 3834
rect 11500 3782 11514 3834
rect 11538 3782 11552 3834
rect 11552 3782 11564 3834
rect 11564 3782 11594 3834
rect 11618 3782 11628 3834
rect 11628 3782 11674 3834
rect 11378 3780 11434 3782
rect 11458 3780 11514 3782
rect 11538 3780 11594 3782
rect 11618 3780 11674 3782
rect 18326 3834 18382 3836
rect 18406 3834 18462 3836
rect 18486 3834 18542 3836
rect 18566 3834 18622 3836
rect 18326 3782 18372 3834
rect 18372 3782 18382 3834
rect 18406 3782 18436 3834
rect 18436 3782 18448 3834
rect 18448 3782 18462 3834
rect 18486 3782 18500 3834
rect 18500 3782 18512 3834
rect 18512 3782 18542 3834
rect 18566 3782 18576 3834
rect 18576 3782 18622 3834
rect 18326 3780 18382 3782
rect 18406 3780 18462 3782
rect 18486 3780 18542 3782
rect 18566 3780 18622 3782
rect 25274 3834 25330 3836
rect 25354 3834 25410 3836
rect 25434 3834 25490 3836
rect 25514 3834 25570 3836
rect 25274 3782 25320 3834
rect 25320 3782 25330 3834
rect 25354 3782 25384 3834
rect 25384 3782 25396 3834
rect 25396 3782 25410 3834
rect 25434 3782 25448 3834
rect 25448 3782 25460 3834
rect 25460 3782 25490 3834
rect 25514 3782 25524 3834
rect 25524 3782 25570 3834
rect 25274 3780 25330 3782
rect 25354 3780 25410 3782
rect 25434 3780 25490 3782
rect 25514 3780 25570 3782
rect 7904 3290 7960 3292
rect 7984 3290 8040 3292
rect 8064 3290 8120 3292
rect 8144 3290 8200 3292
rect 7904 3238 7950 3290
rect 7950 3238 7960 3290
rect 7984 3238 8014 3290
rect 8014 3238 8026 3290
rect 8026 3238 8040 3290
rect 8064 3238 8078 3290
rect 8078 3238 8090 3290
rect 8090 3238 8120 3290
rect 8144 3238 8154 3290
rect 8154 3238 8200 3290
rect 7904 3236 7960 3238
rect 7984 3236 8040 3238
rect 8064 3236 8120 3238
rect 8144 3236 8200 3238
rect 14852 3290 14908 3292
rect 14932 3290 14988 3292
rect 15012 3290 15068 3292
rect 15092 3290 15148 3292
rect 14852 3238 14898 3290
rect 14898 3238 14908 3290
rect 14932 3238 14962 3290
rect 14962 3238 14974 3290
rect 14974 3238 14988 3290
rect 15012 3238 15026 3290
rect 15026 3238 15038 3290
rect 15038 3238 15068 3290
rect 15092 3238 15102 3290
rect 15102 3238 15148 3290
rect 14852 3236 14908 3238
rect 14932 3236 14988 3238
rect 15012 3236 15068 3238
rect 15092 3236 15148 3238
rect 21800 3290 21856 3292
rect 21880 3290 21936 3292
rect 21960 3290 22016 3292
rect 22040 3290 22096 3292
rect 21800 3238 21846 3290
rect 21846 3238 21856 3290
rect 21880 3238 21910 3290
rect 21910 3238 21922 3290
rect 21922 3238 21936 3290
rect 21960 3238 21974 3290
rect 21974 3238 21986 3290
rect 21986 3238 22016 3290
rect 22040 3238 22050 3290
rect 22050 3238 22096 3290
rect 21800 3236 21856 3238
rect 21880 3236 21936 3238
rect 21960 3236 22016 3238
rect 22040 3236 22096 3238
rect 11378 2746 11434 2748
rect 11458 2746 11514 2748
rect 11538 2746 11594 2748
rect 11618 2746 11674 2748
rect 11378 2694 11424 2746
rect 11424 2694 11434 2746
rect 11458 2694 11488 2746
rect 11488 2694 11500 2746
rect 11500 2694 11514 2746
rect 11538 2694 11552 2746
rect 11552 2694 11564 2746
rect 11564 2694 11594 2746
rect 11618 2694 11628 2746
rect 11628 2694 11674 2746
rect 11378 2692 11434 2694
rect 11458 2692 11514 2694
rect 11538 2692 11594 2694
rect 11618 2692 11674 2694
rect 18326 2746 18382 2748
rect 18406 2746 18462 2748
rect 18486 2746 18542 2748
rect 18566 2746 18622 2748
rect 18326 2694 18372 2746
rect 18372 2694 18382 2746
rect 18406 2694 18436 2746
rect 18436 2694 18448 2746
rect 18448 2694 18462 2746
rect 18486 2694 18500 2746
rect 18500 2694 18512 2746
rect 18512 2694 18542 2746
rect 18566 2694 18576 2746
rect 18576 2694 18622 2746
rect 18326 2692 18382 2694
rect 18406 2692 18462 2694
rect 18486 2692 18542 2694
rect 18566 2692 18622 2694
rect 25274 2746 25330 2748
rect 25354 2746 25410 2748
rect 25434 2746 25490 2748
rect 25514 2746 25570 2748
rect 25274 2694 25320 2746
rect 25320 2694 25330 2746
rect 25354 2694 25384 2746
rect 25384 2694 25396 2746
rect 25396 2694 25410 2746
rect 25434 2694 25448 2746
rect 25448 2694 25460 2746
rect 25460 2694 25490 2746
rect 25514 2694 25524 2746
rect 25524 2694 25570 2746
rect 25274 2692 25330 2694
rect 25354 2692 25410 2694
rect 25434 2692 25490 2694
rect 25514 2692 25570 2694
rect 7904 2202 7960 2204
rect 7984 2202 8040 2204
rect 8064 2202 8120 2204
rect 8144 2202 8200 2204
rect 7904 2150 7950 2202
rect 7950 2150 7960 2202
rect 7984 2150 8014 2202
rect 8014 2150 8026 2202
rect 8026 2150 8040 2202
rect 8064 2150 8078 2202
rect 8078 2150 8090 2202
rect 8090 2150 8120 2202
rect 8144 2150 8154 2202
rect 8154 2150 8200 2202
rect 7904 2148 7960 2150
rect 7984 2148 8040 2150
rect 8064 2148 8120 2150
rect 8144 2148 8200 2150
rect 14852 2202 14908 2204
rect 14932 2202 14988 2204
rect 15012 2202 15068 2204
rect 15092 2202 15148 2204
rect 14852 2150 14898 2202
rect 14898 2150 14908 2202
rect 14932 2150 14962 2202
rect 14962 2150 14974 2202
rect 14974 2150 14988 2202
rect 15012 2150 15026 2202
rect 15026 2150 15038 2202
rect 15038 2150 15068 2202
rect 15092 2150 15102 2202
rect 15102 2150 15148 2202
rect 14852 2148 14908 2150
rect 14932 2148 14988 2150
rect 15012 2148 15068 2150
rect 15092 2148 15148 2150
rect 21800 2202 21856 2204
rect 21880 2202 21936 2204
rect 21960 2202 22016 2204
rect 22040 2202 22096 2204
rect 21800 2150 21846 2202
rect 21846 2150 21856 2202
rect 21880 2150 21910 2202
rect 21910 2150 21922 2202
rect 21922 2150 21936 2202
rect 21960 2150 21974 2202
rect 21974 2150 21986 2202
rect 21986 2150 22016 2202
rect 22040 2150 22050 2202
rect 22050 2150 22096 2202
rect 21800 2148 21856 2150
rect 21880 2148 21936 2150
rect 21960 2148 22016 2150
rect 22040 2148 22096 2150
<< metal3 >>
rect 0 29248 800 29368
rect 29200 28568 30000 28688
rect 0 27888 800 28008
rect 29200 27888 30000 28008
rect 4420 27776 4736 27777
rect 4420 27712 4426 27776
rect 4490 27712 4506 27776
rect 4570 27712 4586 27776
rect 4650 27712 4666 27776
rect 4730 27712 4736 27776
rect 4420 27711 4736 27712
rect 11368 27776 11684 27777
rect 11368 27712 11374 27776
rect 11438 27712 11454 27776
rect 11518 27712 11534 27776
rect 11598 27712 11614 27776
rect 11678 27712 11684 27776
rect 11368 27711 11684 27712
rect 18316 27776 18632 27777
rect 18316 27712 18322 27776
rect 18386 27712 18402 27776
rect 18466 27712 18482 27776
rect 18546 27712 18562 27776
rect 18626 27712 18632 27776
rect 18316 27711 18632 27712
rect 25264 27776 25580 27777
rect 25264 27712 25270 27776
rect 25334 27712 25350 27776
rect 25414 27712 25430 27776
rect 25494 27712 25510 27776
rect 25574 27712 25580 27776
rect 25264 27711 25580 27712
rect 0 27208 800 27328
rect 7894 27232 8210 27233
rect 7894 27168 7900 27232
rect 7964 27168 7980 27232
rect 8044 27168 8060 27232
rect 8124 27168 8140 27232
rect 8204 27168 8210 27232
rect 7894 27167 8210 27168
rect 14842 27232 15158 27233
rect 14842 27168 14848 27232
rect 14912 27168 14928 27232
rect 14992 27168 15008 27232
rect 15072 27168 15088 27232
rect 15152 27168 15158 27232
rect 14842 27167 15158 27168
rect 21790 27232 22106 27233
rect 21790 27168 21796 27232
rect 21860 27168 21876 27232
rect 21940 27168 21956 27232
rect 22020 27168 22036 27232
rect 22100 27168 22106 27232
rect 21790 27167 22106 27168
rect 4420 26688 4736 26689
rect 0 26528 800 26648
rect 4420 26624 4426 26688
rect 4490 26624 4506 26688
rect 4570 26624 4586 26688
rect 4650 26624 4666 26688
rect 4730 26624 4736 26688
rect 4420 26623 4736 26624
rect 11368 26688 11684 26689
rect 11368 26624 11374 26688
rect 11438 26624 11454 26688
rect 11518 26624 11534 26688
rect 11598 26624 11614 26688
rect 11678 26624 11684 26688
rect 11368 26623 11684 26624
rect 18316 26688 18632 26689
rect 18316 26624 18322 26688
rect 18386 26624 18402 26688
rect 18466 26624 18482 26688
rect 18546 26624 18562 26688
rect 18626 26624 18632 26688
rect 18316 26623 18632 26624
rect 25264 26688 25580 26689
rect 25264 26624 25270 26688
rect 25334 26624 25350 26688
rect 25414 26624 25430 26688
rect 25494 26624 25510 26688
rect 25574 26624 25580 26688
rect 25264 26623 25580 26624
rect 29200 26528 30000 26648
rect 7894 26144 8210 26145
rect 7894 26080 7900 26144
rect 7964 26080 7980 26144
rect 8044 26080 8060 26144
rect 8124 26080 8140 26144
rect 8204 26080 8210 26144
rect 7894 26079 8210 26080
rect 14842 26144 15158 26145
rect 14842 26080 14848 26144
rect 14912 26080 14928 26144
rect 14992 26080 15008 26144
rect 15072 26080 15088 26144
rect 15152 26080 15158 26144
rect 14842 26079 15158 26080
rect 21790 26144 22106 26145
rect 21790 26080 21796 26144
rect 21860 26080 21876 26144
rect 21940 26080 21956 26144
rect 22020 26080 22036 26144
rect 22100 26080 22106 26144
rect 21790 26079 22106 26080
rect 29200 25848 30000 25968
rect 4420 25600 4736 25601
rect 4420 25536 4426 25600
rect 4490 25536 4506 25600
rect 4570 25536 4586 25600
rect 4650 25536 4666 25600
rect 4730 25536 4736 25600
rect 4420 25535 4736 25536
rect 11368 25600 11684 25601
rect 11368 25536 11374 25600
rect 11438 25536 11454 25600
rect 11518 25536 11534 25600
rect 11598 25536 11614 25600
rect 11678 25536 11684 25600
rect 11368 25535 11684 25536
rect 18316 25600 18632 25601
rect 18316 25536 18322 25600
rect 18386 25536 18402 25600
rect 18466 25536 18482 25600
rect 18546 25536 18562 25600
rect 18626 25536 18632 25600
rect 18316 25535 18632 25536
rect 25264 25600 25580 25601
rect 25264 25536 25270 25600
rect 25334 25536 25350 25600
rect 25414 25536 25430 25600
rect 25494 25536 25510 25600
rect 25574 25536 25580 25600
rect 25264 25535 25580 25536
rect 0 25168 800 25288
rect 29200 25168 30000 25288
rect 7894 25056 8210 25057
rect 7894 24992 7900 25056
rect 7964 24992 7980 25056
rect 8044 24992 8060 25056
rect 8124 24992 8140 25056
rect 8204 24992 8210 25056
rect 7894 24991 8210 24992
rect 14842 25056 15158 25057
rect 14842 24992 14848 25056
rect 14912 24992 14928 25056
rect 14992 24992 15008 25056
rect 15072 24992 15088 25056
rect 15152 24992 15158 25056
rect 14842 24991 15158 24992
rect 21790 25056 22106 25057
rect 21790 24992 21796 25056
rect 21860 24992 21876 25056
rect 21940 24992 21956 25056
rect 22020 24992 22036 25056
rect 22100 24992 22106 25056
rect 21790 24991 22106 24992
rect 0 24488 800 24608
rect 4420 24512 4736 24513
rect 4420 24448 4426 24512
rect 4490 24448 4506 24512
rect 4570 24448 4586 24512
rect 4650 24448 4666 24512
rect 4730 24448 4736 24512
rect 4420 24447 4736 24448
rect 11368 24512 11684 24513
rect 11368 24448 11374 24512
rect 11438 24448 11454 24512
rect 11518 24448 11534 24512
rect 11598 24448 11614 24512
rect 11678 24448 11684 24512
rect 11368 24447 11684 24448
rect 18316 24512 18632 24513
rect 18316 24448 18322 24512
rect 18386 24448 18402 24512
rect 18466 24448 18482 24512
rect 18546 24448 18562 24512
rect 18626 24448 18632 24512
rect 18316 24447 18632 24448
rect 25264 24512 25580 24513
rect 25264 24448 25270 24512
rect 25334 24448 25350 24512
rect 25414 24448 25430 24512
rect 25494 24448 25510 24512
rect 25574 24448 25580 24512
rect 25264 24447 25580 24448
rect 7894 23968 8210 23969
rect 7894 23904 7900 23968
rect 7964 23904 7980 23968
rect 8044 23904 8060 23968
rect 8124 23904 8140 23968
rect 8204 23904 8210 23968
rect 7894 23903 8210 23904
rect 14842 23968 15158 23969
rect 14842 23904 14848 23968
rect 14912 23904 14928 23968
rect 14992 23904 15008 23968
rect 15072 23904 15088 23968
rect 15152 23904 15158 23968
rect 14842 23903 15158 23904
rect 21790 23968 22106 23969
rect 21790 23904 21796 23968
rect 21860 23904 21876 23968
rect 21940 23904 21956 23968
rect 22020 23904 22036 23968
rect 22100 23904 22106 23968
rect 21790 23903 22106 23904
rect 29200 23808 30000 23928
rect 4420 23424 4736 23425
rect 4420 23360 4426 23424
rect 4490 23360 4506 23424
rect 4570 23360 4586 23424
rect 4650 23360 4666 23424
rect 4730 23360 4736 23424
rect 4420 23359 4736 23360
rect 11368 23424 11684 23425
rect 11368 23360 11374 23424
rect 11438 23360 11454 23424
rect 11518 23360 11534 23424
rect 11598 23360 11614 23424
rect 11678 23360 11684 23424
rect 11368 23359 11684 23360
rect 18316 23424 18632 23425
rect 18316 23360 18322 23424
rect 18386 23360 18402 23424
rect 18466 23360 18482 23424
rect 18546 23360 18562 23424
rect 18626 23360 18632 23424
rect 18316 23359 18632 23360
rect 25264 23424 25580 23425
rect 25264 23360 25270 23424
rect 25334 23360 25350 23424
rect 25414 23360 25430 23424
rect 25494 23360 25510 23424
rect 25574 23360 25580 23424
rect 25264 23359 25580 23360
rect 0 23128 800 23248
rect 29200 23128 30000 23248
rect 7894 22880 8210 22881
rect 7894 22816 7900 22880
rect 7964 22816 7980 22880
rect 8044 22816 8060 22880
rect 8124 22816 8140 22880
rect 8204 22816 8210 22880
rect 7894 22815 8210 22816
rect 14842 22880 15158 22881
rect 14842 22816 14848 22880
rect 14912 22816 14928 22880
rect 14992 22816 15008 22880
rect 15072 22816 15088 22880
rect 15152 22816 15158 22880
rect 14842 22815 15158 22816
rect 21790 22880 22106 22881
rect 21790 22816 21796 22880
rect 21860 22816 21876 22880
rect 21940 22816 21956 22880
rect 22020 22816 22036 22880
rect 22100 22816 22106 22880
rect 21790 22815 22106 22816
rect 0 22448 800 22568
rect 4420 22336 4736 22337
rect 4420 22272 4426 22336
rect 4490 22272 4506 22336
rect 4570 22272 4586 22336
rect 4650 22272 4666 22336
rect 4730 22272 4736 22336
rect 4420 22271 4736 22272
rect 11368 22336 11684 22337
rect 11368 22272 11374 22336
rect 11438 22272 11454 22336
rect 11518 22272 11534 22336
rect 11598 22272 11614 22336
rect 11678 22272 11684 22336
rect 11368 22271 11684 22272
rect 18316 22336 18632 22337
rect 18316 22272 18322 22336
rect 18386 22272 18402 22336
rect 18466 22272 18482 22336
rect 18546 22272 18562 22336
rect 18626 22272 18632 22336
rect 18316 22271 18632 22272
rect 25264 22336 25580 22337
rect 25264 22272 25270 22336
rect 25334 22272 25350 22336
rect 25414 22272 25430 22336
rect 25494 22272 25510 22336
rect 25574 22272 25580 22336
rect 25264 22271 25580 22272
rect 0 21768 800 21888
rect 7894 21792 8210 21793
rect 7894 21728 7900 21792
rect 7964 21728 7980 21792
rect 8044 21728 8060 21792
rect 8124 21728 8140 21792
rect 8204 21728 8210 21792
rect 7894 21727 8210 21728
rect 14842 21792 15158 21793
rect 14842 21728 14848 21792
rect 14912 21728 14928 21792
rect 14992 21728 15008 21792
rect 15072 21728 15088 21792
rect 15152 21728 15158 21792
rect 14842 21727 15158 21728
rect 21790 21792 22106 21793
rect 21790 21728 21796 21792
rect 21860 21728 21876 21792
rect 21940 21728 21956 21792
rect 22020 21728 22036 21792
rect 22100 21728 22106 21792
rect 29200 21768 30000 21888
rect 21790 21727 22106 21728
rect 4420 21248 4736 21249
rect 4420 21184 4426 21248
rect 4490 21184 4506 21248
rect 4570 21184 4586 21248
rect 4650 21184 4666 21248
rect 4730 21184 4736 21248
rect 4420 21183 4736 21184
rect 11368 21248 11684 21249
rect 11368 21184 11374 21248
rect 11438 21184 11454 21248
rect 11518 21184 11534 21248
rect 11598 21184 11614 21248
rect 11678 21184 11684 21248
rect 11368 21183 11684 21184
rect 18316 21248 18632 21249
rect 18316 21184 18322 21248
rect 18386 21184 18402 21248
rect 18466 21184 18482 21248
rect 18546 21184 18562 21248
rect 18626 21184 18632 21248
rect 18316 21183 18632 21184
rect 25264 21248 25580 21249
rect 25264 21184 25270 21248
rect 25334 21184 25350 21248
rect 25414 21184 25430 21248
rect 25494 21184 25510 21248
rect 25574 21184 25580 21248
rect 25264 21183 25580 21184
rect 29200 21088 30000 21208
rect 7894 20704 8210 20705
rect 7894 20640 7900 20704
rect 7964 20640 7980 20704
rect 8044 20640 8060 20704
rect 8124 20640 8140 20704
rect 8204 20640 8210 20704
rect 7894 20639 8210 20640
rect 14842 20704 15158 20705
rect 14842 20640 14848 20704
rect 14912 20640 14928 20704
rect 14992 20640 15008 20704
rect 15072 20640 15088 20704
rect 15152 20640 15158 20704
rect 14842 20639 15158 20640
rect 21790 20704 22106 20705
rect 21790 20640 21796 20704
rect 21860 20640 21876 20704
rect 21940 20640 21956 20704
rect 22020 20640 22036 20704
rect 22100 20640 22106 20704
rect 21790 20639 22106 20640
rect 0 20408 800 20528
rect 29200 20408 30000 20528
rect 4420 20160 4736 20161
rect 4420 20096 4426 20160
rect 4490 20096 4506 20160
rect 4570 20096 4586 20160
rect 4650 20096 4666 20160
rect 4730 20096 4736 20160
rect 4420 20095 4736 20096
rect 11368 20160 11684 20161
rect 11368 20096 11374 20160
rect 11438 20096 11454 20160
rect 11518 20096 11534 20160
rect 11598 20096 11614 20160
rect 11678 20096 11684 20160
rect 11368 20095 11684 20096
rect 18316 20160 18632 20161
rect 18316 20096 18322 20160
rect 18386 20096 18402 20160
rect 18466 20096 18482 20160
rect 18546 20096 18562 20160
rect 18626 20096 18632 20160
rect 18316 20095 18632 20096
rect 25264 20160 25580 20161
rect 25264 20096 25270 20160
rect 25334 20096 25350 20160
rect 25414 20096 25430 20160
rect 25494 20096 25510 20160
rect 25574 20096 25580 20160
rect 25264 20095 25580 20096
rect 0 19728 800 19848
rect 7894 19616 8210 19617
rect 7894 19552 7900 19616
rect 7964 19552 7980 19616
rect 8044 19552 8060 19616
rect 8124 19552 8140 19616
rect 8204 19552 8210 19616
rect 7894 19551 8210 19552
rect 14842 19616 15158 19617
rect 14842 19552 14848 19616
rect 14912 19552 14928 19616
rect 14992 19552 15008 19616
rect 15072 19552 15088 19616
rect 15152 19552 15158 19616
rect 14842 19551 15158 19552
rect 21790 19616 22106 19617
rect 21790 19552 21796 19616
rect 21860 19552 21876 19616
rect 21940 19552 21956 19616
rect 22020 19552 22036 19616
rect 22100 19552 22106 19616
rect 21790 19551 22106 19552
rect 4420 19072 4736 19073
rect 4420 19008 4426 19072
rect 4490 19008 4506 19072
rect 4570 19008 4586 19072
rect 4650 19008 4666 19072
rect 4730 19008 4736 19072
rect 4420 19007 4736 19008
rect 11368 19072 11684 19073
rect 11368 19008 11374 19072
rect 11438 19008 11454 19072
rect 11518 19008 11534 19072
rect 11598 19008 11614 19072
rect 11678 19008 11684 19072
rect 11368 19007 11684 19008
rect 18316 19072 18632 19073
rect 18316 19008 18322 19072
rect 18386 19008 18402 19072
rect 18466 19008 18482 19072
rect 18546 19008 18562 19072
rect 18626 19008 18632 19072
rect 18316 19007 18632 19008
rect 25264 19072 25580 19073
rect 25264 19008 25270 19072
rect 25334 19008 25350 19072
rect 25414 19008 25430 19072
rect 25494 19008 25510 19072
rect 25574 19008 25580 19072
rect 29200 19048 30000 19168
rect 25264 19007 25580 19008
rect 7894 18528 8210 18529
rect 0 18368 800 18488
rect 7894 18464 7900 18528
rect 7964 18464 7980 18528
rect 8044 18464 8060 18528
rect 8124 18464 8140 18528
rect 8204 18464 8210 18528
rect 7894 18463 8210 18464
rect 14842 18528 15158 18529
rect 14842 18464 14848 18528
rect 14912 18464 14928 18528
rect 14992 18464 15008 18528
rect 15072 18464 15088 18528
rect 15152 18464 15158 18528
rect 14842 18463 15158 18464
rect 21790 18528 22106 18529
rect 21790 18464 21796 18528
rect 21860 18464 21876 18528
rect 21940 18464 21956 18528
rect 22020 18464 22036 18528
rect 22100 18464 22106 18528
rect 21790 18463 22106 18464
rect 29200 18368 30000 18488
rect 4420 17984 4736 17985
rect 4420 17920 4426 17984
rect 4490 17920 4506 17984
rect 4570 17920 4586 17984
rect 4650 17920 4666 17984
rect 4730 17920 4736 17984
rect 4420 17919 4736 17920
rect 11368 17984 11684 17985
rect 11368 17920 11374 17984
rect 11438 17920 11454 17984
rect 11518 17920 11534 17984
rect 11598 17920 11614 17984
rect 11678 17920 11684 17984
rect 11368 17919 11684 17920
rect 18316 17984 18632 17985
rect 18316 17920 18322 17984
rect 18386 17920 18402 17984
rect 18466 17920 18482 17984
rect 18546 17920 18562 17984
rect 18626 17920 18632 17984
rect 18316 17919 18632 17920
rect 25264 17984 25580 17985
rect 25264 17920 25270 17984
rect 25334 17920 25350 17984
rect 25414 17920 25430 17984
rect 25494 17920 25510 17984
rect 25574 17920 25580 17984
rect 25264 17919 25580 17920
rect 0 17688 800 17808
rect 7894 17440 8210 17441
rect 7894 17376 7900 17440
rect 7964 17376 7980 17440
rect 8044 17376 8060 17440
rect 8124 17376 8140 17440
rect 8204 17376 8210 17440
rect 7894 17375 8210 17376
rect 14842 17440 15158 17441
rect 14842 17376 14848 17440
rect 14912 17376 14928 17440
rect 14992 17376 15008 17440
rect 15072 17376 15088 17440
rect 15152 17376 15158 17440
rect 14842 17375 15158 17376
rect 21790 17440 22106 17441
rect 21790 17376 21796 17440
rect 21860 17376 21876 17440
rect 21940 17376 21956 17440
rect 22020 17376 22036 17440
rect 22100 17376 22106 17440
rect 21790 17375 22106 17376
rect 0 17008 800 17128
rect 29200 17008 30000 17128
rect 4420 16896 4736 16897
rect 4420 16832 4426 16896
rect 4490 16832 4506 16896
rect 4570 16832 4586 16896
rect 4650 16832 4666 16896
rect 4730 16832 4736 16896
rect 4420 16831 4736 16832
rect 11368 16896 11684 16897
rect 11368 16832 11374 16896
rect 11438 16832 11454 16896
rect 11518 16832 11534 16896
rect 11598 16832 11614 16896
rect 11678 16832 11684 16896
rect 11368 16831 11684 16832
rect 18316 16896 18632 16897
rect 18316 16832 18322 16896
rect 18386 16832 18402 16896
rect 18466 16832 18482 16896
rect 18546 16832 18562 16896
rect 18626 16832 18632 16896
rect 18316 16831 18632 16832
rect 25264 16896 25580 16897
rect 25264 16832 25270 16896
rect 25334 16832 25350 16896
rect 25414 16832 25430 16896
rect 25494 16832 25510 16896
rect 25574 16832 25580 16896
rect 25264 16831 25580 16832
rect 7894 16352 8210 16353
rect 7894 16288 7900 16352
rect 7964 16288 7980 16352
rect 8044 16288 8060 16352
rect 8124 16288 8140 16352
rect 8204 16288 8210 16352
rect 7894 16287 8210 16288
rect 14842 16352 15158 16353
rect 14842 16288 14848 16352
rect 14912 16288 14928 16352
rect 14992 16288 15008 16352
rect 15072 16288 15088 16352
rect 15152 16288 15158 16352
rect 14842 16287 15158 16288
rect 21790 16352 22106 16353
rect 21790 16288 21796 16352
rect 21860 16288 21876 16352
rect 21940 16288 21956 16352
rect 22020 16288 22036 16352
rect 22100 16288 22106 16352
rect 29200 16328 30000 16448
rect 21790 16287 22106 16288
rect 4420 15808 4736 15809
rect 0 15648 800 15768
rect 4420 15744 4426 15808
rect 4490 15744 4506 15808
rect 4570 15744 4586 15808
rect 4650 15744 4666 15808
rect 4730 15744 4736 15808
rect 4420 15743 4736 15744
rect 11368 15808 11684 15809
rect 11368 15744 11374 15808
rect 11438 15744 11454 15808
rect 11518 15744 11534 15808
rect 11598 15744 11614 15808
rect 11678 15744 11684 15808
rect 11368 15743 11684 15744
rect 18316 15808 18632 15809
rect 18316 15744 18322 15808
rect 18386 15744 18402 15808
rect 18466 15744 18482 15808
rect 18546 15744 18562 15808
rect 18626 15744 18632 15808
rect 18316 15743 18632 15744
rect 25264 15808 25580 15809
rect 25264 15744 25270 15808
rect 25334 15744 25350 15808
rect 25414 15744 25430 15808
rect 25494 15744 25510 15808
rect 25574 15744 25580 15808
rect 25264 15743 25580 15744
rect 29200 15648 30000 15768
rect 7894 15264 8210 15265
rect 7894 15200 7900 15264
rect 7964 15200 7980 15264
rect 8044 15200 8060 15264
rect 8124 15200 8140 15264
rect 8204 15200 8210 15264
rect 7894 15199 8210 15200
rect 14842 15264 15158 15265
rect 14842 15200 14848 15264
rect 14912 15200 14928 15264
rect 14992 15200 15008 15264
rect 15072 15200 15088 15264
rect 15152 15200 15158 15264
rect 14842 15199 15158 15200
rect 21790 15264 22106 15265
rect 21790 15200 21796 15264
rect 21860 15200 21876 15264
rect 21940 15200 21956 15264
rect 22020 15200 22036 15264
rect 22100 15200 22106 15264
rect 21790 15199 22106 15200
rect 0 14968 800 15088
rect 4420 14720 4736 14721
rect 4420 14656 4426 14720
rect 4490 14656 4506 14720
rect 4570 14656 4586 14720
rect 4650 14656 4666 14720
rect 4730 14656 4736 14720
rect 4420 14655 4736 14656
rect 11368 14720 11684 14721
rect 11368 14656 11374 14720
rect 11438 14656 11454 14720
rect 11518 14656 11534 14720
rect 11598 14656 11614 14720
rect 11678 14656 11684 14720
rect 11368 14655 11684 14656
rect 18316 14720 18632 14721
rect 18316 14656 18322 14720
rect 18386 14656 18402 14720
rect 18466 14656 18482 14720
rect 18546 14656 18562 14720
rect 18626 14656 18632 14720
rect 18316 14655 18632 14656
rect 25264 14720 25580 14721
rect 25264 14656 25270 14720
rect 25334 14656 25350 14720
rect 25414 14656 25430 14720
rect 25494 14656 25510 14720
rect 25574 14656 25580 14720
rect 25264 14655 25580 14656
rect 29200 14288 30000 14408
rect 7894 14176 8210 14177
rect 7894 14112 7900 14176
rect 7964 14112 7980 14176
rect 8044 14112 8060 14176
rect 8124 14112 8140 14176
rect 8204 14112 8210 14176
rect 7894 14111 8210 14112
rect 14842 14176 15158 14177
rect 14842 14112 14848 14176
rect 14912 14112 14928 14176
rect 14992 14112 15008 14176
rect 15072 14112 15088 14176
rect 15152 14112 15158 14176
rect 14842 14111 15158 14112
rect 21790 14176 22106 14177
rect 21790 14112 21796 14176
rect 21860 14112 21876 14176
rect 21940 14112 21956 14176
rect 22020 14112 22036 14176
rect 22100 14112 22106 14176
rect 21790 14111 22106 14112
rect 0 13608 800 13728
rect 28165 13698 28231 13701
rect 29200 13698 30000 13728
rect 28165 13696 30000 13698
rect 28165 13640 28170 13696
rect 28226 13640 30000 13696
rect 28165 13638 30000 13640
rect 28165 13635 28231 13638
rect 4420 13632 4736 13633
rect 4420 13568 4426 13632
rect 4490 13568 4506 13632
rect 4570 13568 4586 13632
rect 4650 13568 4666 13632
rect 4730 13568 4736 13632
rect 4420 13567 4736 13568
rect 11368 13632 11684 13633
rect 11368 13568 11374 13632
rect 11438 13568 11454 13632
rect 11518 13568 11534 13632
rect 11598 13568 11614 13632
rect 11678 13568 11684 13632
rect 11368 13567 11684 13568
rect 18316 13632 18632 13633
rect 18316 13568 18322 13632
rect 18386 13568 18402 13632
rect 18466 13568 18482 13632
rect 18546 13568 18562 13632
rect 18626 13568 18632 13632
rect 18316 13567 18632 13568
rect 25264 13632 25580 13633
rect 25264 13568 25270 13632
rect 25334 13568 25350 13632
rect 25414 13568 25430 13632
rect 25494 13568 25510 13632
rect 25574 13568 25580 13632
rect 29200 13608 30000 13638
rect 25264 13567 25580 13568
rect 7894 13088 8210 13089
rect 0 12928 800 13048
rect 7894 13024 7900 13088
rect 7964 13024 7980 13088
rect 8044 13024 8060 13088
rect 8124 13024 8140 13088
rect 8204 13024 8210 13088
rect 7894 13023 8210 13024
rect 14842 13088 15158 13089
rect 14842 13024 14848 13088
rect 14912 13024 14928 13088
rect 14992 13024 15008 13088
rect 15072 13024 15088 13088
rect 15152 13024 15158 13088
rect 14842 13023 15158 13024
rect 21790 13088 22106 13089
rect 21790 13024 21796 13088
rect 21860 13024 21876 13088
rect 21940 13024 21956 13088
rect 22020 13024 22036 13088
rect 22100 13024 22106 13088
rect 21790 13023 22106 13024
rect 4420 12544 4736 12545
rect 4420 12480 4426 12544
rect 4490 12480 4506 12544
rect 4570 12480 4586 12544
rect 4650 12480 4666 12544
rect 4730 12480 4736 12544
rect 4420 12479 4736 12480
rect 11368 12544 11684 12545
rect 11368 12480 11374 12544
rect 11438 12480 11454 12544
rect 11518 12480 11534 12544
rect 11598 12480 11614 12544
rect 11678 12480 11684 12544
rect 11368 12479 11684 12480
rect 18316 12544 18632 12545
rect 18316 12480 18322 12544
rect 18386 12480 18402 12544
rect 18466 12480 18482 12544
rect 18546 12480 18562 12544
rect 18626 12480 18632 12544
rect 18316 12479 18632 12480
rect 25264 12544 25580 12545
rect 25264 12480 25270 12544
rect 25334 12480 25350 12544
rect 25414 12480 25430 12544
rect 25494 12480 25510 12544
rect 25574 12480 25580 12544
rect 25264 12479 25580 12480
rect 0 12248 800 12368
rect 29200 12248 30000 12368
rect 7894 12000 8210 12001
rect 7894 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8210 12000
rect 7894 11935 8210 11936
rect 14842 12000 15158 12001
rect 14842 11936 14848 12000
rect 14912 11936 14928 12000
rect 14992 11936 15008 12000
rect 15072 11936 15088 12000
rect 15152 11936 15158 12000
rect 14842 11935 15158 11936
rect 21790 12000 22106 12001
rect 21790 11936 21796 12000
rect 21860 11936 21876 12000
rect 21940 11936 21956 12000
rect 22020 11936 22036 12000
rect 22100 11936 22106 12000
rect 21790 11935 22106 11936
rect 29200 11568 30000 11688
rect 4420 11456 4736 11457
rect 4420 11392 4426 11456
rect 4490 11392 4506 11456
rect 4570 11392 4586 11456
rect 4650 11392 4666 11456
rect 4730 11392 4736 11456
rect 4420 11391 4736 11392
rect 11368 11456 11684 11457
rect 11368 11392 11374 11456
rect 11438 11392 11454 11456
rect 11518 11392 11534 11456
rect 11598 11392 11614 11456
rect 11678 11392 11684 11456
rect 11368 11391 11684 11392
rect 18316 11456 18632 11457
rect 18316 11392 18322 11456
rect 18386 11392 18402 11456
rect 18466 11392 18482 11456
rect 18546 11392 18562 11456
rect 18626 11392 18632 11456
rect 18316 11391 18632 11392
rect 25264 11456 25580 11457
rect 25264 11392 25270 11456
rect 25334 11392 25350 11456
rect 25414 11392 25430 11456
rect 25494 11392 25510 11456
rect 25574 11392 25580 11456
rect 25264 11391 25580 11392
rect 0 10888 800 11008
rect 7894 10912 8210 10913
rect 7894 10848 7900 10912
rect 7964 10848 7980 10912
rect 8044 10848 8060 10912
rect 8124 10848 8140 10912
rect 8204 10848 8210 10912
rect 7894 10847 8210 10848
rect 14842 10912 15158 10913
rect 14842 10848 14848 10912
rect 14912 10848 14928 10912
rect 14992 10848 15008 10912
rect 15072 10848 15088 10912
rect 15152 10848 15158 10912
rect 14842 10847 15158 10848
rect 21790 10912 22106 10913
rect 21790 10848 21796 10912
rect 21860 10848 21876 10912
rect 21940 10848 21956 10912
rect 22020 10848 22036 10912
rect 22100 10848 22106 10912
rect 21790 10847 22106 10848
rect 4420 10368 4736 10369
rect 0 10208 800 10328
rect 4420 10304 4426 10368
rect 4490 10304 4506 10368
rect 4570 10304 4586 10368
rect 4650 10304 4666 10368
rect 4730 10304 4736 10368
rect 4420 10303 4736 10304
rect 11368 10368 11684 10369
rect 11368 10304 11374 10368
rect 11438 10304 11454 10368
rect 11518 10304 11534 10368
rect 11598 10304 11614 10368
rect 11678 10304 11684 10368
rect 11368 10303 11684 10304
rect 18316 10368 18632 10369
rect 18316 10304 18322 10368
rect 18386 10304 18402 10368
rect 18466 10304 18482 10368
rect 18546 10304 18562 10368
rect 18626 10304 18632 10368
rect 18316 10303 18632 10304
rect 25264 10368 25580 10369
rect 25264 10304 25270 10368
rect 25334 10304 25350 10368
rect 25414 10304 25430 10368
rect 25494 10304 25510 10368
rect 25574 10304 25580 10368
rect 25264 10303 25580 10304
rect 29200 10208 30000 10328
rect 7894 9824 8210 9825
rect 7894 9760 7900 9824
rect 7964 9760 7980 9824
rect 8044 9760 8060 9824
rect 8124 9760 8140 9824
rect 8204 9760 8210 9824
rect 7894 9759 8210 9760
rect 14842 9824 15158 9825
rect 14842 9760 14848 9824
rect 14912 9760 14928 9824
rect 14992 9760 15008 9824
rect 15072 9760 15088 9824
rect 15152 9760 15158 9824
rect 14842 9759 15158 9760
rect 21790 9824 22106 9825
rect 21790 9760 21796 9824
rect 21860 9760 21876 9824
rect 21940 9760 21956 9824
rect 22020 9760 22036 9824
rect 22100 9760 22106 9824
rect 21790 9759 22106 9760
rect 27521 9618 27587 9621
rect 29200 9618 30000 9648
rect 27521 9616 30000 9618
rect 27521 9560 27526 9616
rect 27582 9560 30000 9616
rect 27521 9558 30000 9560
rect 27521 9555 27587 9558
rect 29200 9528 30000 9558
rect 4420 9280 4736 9281
rect 4420 9216 4426 9280
rect 4490 9216 4506 9280
rect 4570 9216 4586 9280
rect 4650 9216 4666 9280
rect 4730 9216 4736 9280
rect 4420 9215 4736 9216
rect 11368 9280 11684 9281
rect 11368 9216 11374 9280
rect 11438 9216 11454 9280
rect 11518 9216 11534 9280
rect 11598 9216 11614 9280
rect 11678 9216 11684 9280
rect 11368 9215 11684 9216
rect 18316 9280 18632 9281
rect 18316 9216 18322 9280
rect 18386 9216 18402 9280
rect 18466 9216 18482 9280
rect 18546 9216 18562 9280
rect 18626 9216 18632 9280
rect 18316 9215 18632 9216
rect 25264 9280 25580 9281
rect 25264 9216 25270 9280
rect 25334 9216 25350 9280
rect 25414 9216 25430 9280
rect 25494 9216 25510 9280
rect 25574 9216 25580 9280
rect 25264 9215 25580 9216
rect 0 8848 800 8968
rect 29200 8848 30000 8968
rect 7894 8736 8210 8737
rect 7894 8672 7900 8736
rect 7964 8672 7980 8736
rect 8044 8672 8060 8736
rect 8124 8672 8140 8736
rect 8204 8672 8210 8736
rect 7894 8671 8210 8672
rect 14842 8736 15158 8737
rect 14842 8672 14848 8736
rect 14912 8672 14928 8736
rect 14992 8672 15008 8736
rect 15072 8672 15088 8736
rect 15152 8672 15158 8736
rect 14842 8671 15158 8672
rect 21790 8736 22106 8737
rect 21790 8672 21796 8736
rect 21860 8672 21876 8736
rect 21940 8672 21956 8736
rect 22020 8672 22036 8736
rect 22100 8672 22106 8736
rect 21790 8671 22106 8672
rect 0 8168 800 8288
rect 4420 8192 4736 8193
rect 4420 8128 4426 8192
rect 4490 8128 4506 8192
rect 4570 8128 4586 8192
rect 4650 8128 4666 8192
rect 4730 8128 4736 8192
rect 4420 8127 4736 8128
rect 11368 8192 11684 8193
rect 11368 8128 11374 8192
rect 11438 8128 11454 8192
rect 11518 8128 11534 8192
rect 11598 8128 11614 8192
rect 11678 8128 11684 8192
rect 11368 8127 11684 8128
rect 18316 8192 18632 8193
rect 18316 8128 18322 8192
rect 18386 8128 18402 8192
rect 18466 8128 18482 8192
rect 18546 8128 18562 8192
rect 18626 8128 18632 8192
rect 18316 8127 18632 8128
rect 25264 8192 25580 8193
rect 25264 8128 25270 8192
rect 25334 8128 25350 8192
rect 25414 8128 25430 8192
rect 25494 8128 25510 8192
rect 25574 8128 25580 8192
rect 25264 8127 25580 8128
rect 7894 7648 8210 7649
rect 0 7488 800 7608
rect 7894 7584 7900 7648
rect 7964 7584 7980 7648
rect 8044 7584 8060 7648
rect 8124 7584 8140 7648
rect 8204 7584 8210 7648
rect 7894 7583 8210 7584
rect 14842 7648 15158 7649
rect 14842 7584 14848 7648
rect 14912 7584 14928 7648
rect 14992 7584 15008 7648
rect 15072 7584 15088 7648
rect 15152 7584 15158 7648
rect 14842 7583 15158 7584
rect 21790 7648 22106 7649
rect 21790 7584 21796 7648
rect 21860 7584 21876 7648
rect 21940 7584 21956 7648
rect 22020 7584 22036 7648
rect 22100 7584 22106 7648
rect 21790 7583 22106 7584
rect 29200 7488 30000 7608
rect 4420 7104 4736 7105
rect 4420 7040 4426 7104
rect 4490 7040 4506 7104
rect 4570 7040 4586 7104
rect 4650 7040 4666 7104
rect 4730 7040 4736 7104
rect 4420 7039 4736 7040
rect 11368 7104 11684 7105
rect 11368 7040 11374 7104
rect 11438 7040 11454 7104
rect 11518 7040 11534 7104
rect 11598 7040 11614 7104
rect 11678 7040 11684 7104
rect 11368 7039 11684 7040
rect 18316 7104 18632 7105
rect 18316 7040 18322 7104
rect 18386 7040 18402 7104
rect 18466 7040 18482 7104
rect 18546 7040 18562 7104
rect 18626 7040 18632 7104
rect 18316 7039 18632 7040
rect 25264 7104 25580 7105
rect 25264 7040 25270 7104
rect 25334 7040 25350 7104
rect 25414 7040 25430 7104
rect 25494 7040 25510 7104
rect 25574 7040 25580 7104
rect 25264 7039 25580 7040
rect 29200 6808 30000 6928
rect 7894 6560 8210 6561
rect 7894 6496 7900 6560
rect 7964 6496 7980 6560
rect 8044 6496 8060 6560
rect 8124 6496 8140 6560
rect 8204 6496 8210 6560
rect 7894 6495 8210 6496
rect 14842 6560 15158 6561
rect 14842 6496 14848 6560
rect 14912 6496 14928 6560
rect 14992 6496 15008 6560
rect 15072 6496 15088 6560
rect 15152 6496 15158 6560
rect 14842 6495 15158 6496
rect 21790 6560 22106 6561
rect 21790 6496 21796 6560
rect 21860 6496 21876 6560
rect 21940 6496 21956 6560
rect 22020 6496 22036 6560
rect 22100 6496 22106 6560
rect 21790 6495 22106 6496
rect 0 6128 800 6248
rect 29200 6128 30000 6248
rect 4420 6016 4736 6017
rect 4420 5952 4426 6016
rect 4490 5952 4506 6016
rect 4570 5952 4586 6016
rect 4650 5952 4666 6016
rect 4730 5952 4736 6016
rect 4420 5951 4736 5952
rect 11368 6016 11684 6017
rect 11368 5952 11374 6016
rect 11438 5952 11454 6016
rect 11518 5952 11534 6016
rect 11598 5952 11614 6016
rect 11678 5952 11684 6016
rect 11368 5951 11684 5952
rect 18316 6016 18632 6017
rect 18316 5952 18322 6016
rect 18386 5952 18402 6016
rect 18466 5952 18482 6016
rect 18546 5952 18562 6016
rect 18626 5952 18632 6016
rect 18316 5951 18632 5952
rect 25264 6016 25580 6017
rect 25264 5952 25270 6016
rect 25334 5952 25350 6016
rect 25414 5952 25430 6016
rect 25494 5952 25510 6016
rect 25574 5952 25580 6016
rect 25264 5951 25580 5952
rect 0 5448 800 5568
rect 7894 5472 8210 5473
rect 7894 5408 7900 5472
rect 7964 5408 7980 5472
rect 8044 5408 8060 5472
rect 8124 5408 8140 5472
rect 8204 5408 8210 5472
rect 7894 5407 8210 5408
rect 14842 5472 15158 5473
rect 14842 5408 14848 5472
rect 14912 5408 14928 5472
rect 14992 5408 15008 5472
rect 15072 5408 15088 5472
rect 15152 5408 15158 5472
rect 14842 5407 15158 5408
rect 21790 5472 22106 5473
rect 21790 5408 21796 5472
rect 21860 5408 21876 5472
rect 21940 5408 21956 5472
rect 22020 5408 22036 5472
rect 22100 5408 22106 5472
rect 21790 5407 22106 5408
rect 4420 4928 4736 4929
rect 4420 4864 4426 4928
rect 4490 4864 4506 4928
rect 4570 4864 4586 4928
rect 4650 4864 4666 4928
rect 4730 4864 4736 4928
rect 4420 4863 4736 4864
rect 11368 4928 11684 4929
rect 11368 4864 11374 4928
rect 11438 4864 11454 4928
rect 11518 4864 11534 4928
rect 11598 4864 11614 4928
rect 11678 4864 11684 4928
rect 11368 4863 11684 4864
rect 18316 4928 18632 4929
rect 18316 4864 18322 4928
rect 18386 4864 18402 4928
rect 18466 4864 18482 4928
rect 18546 4864 18562 4928
rect 18626 4864 18632 4928
rect 18316 4863 18632 4864
rect 25264 4928 25580 4929
rect 25264 4864 25270 4928
rect 25334 4864 25350 4928
rect 25414 4864 25430 4928
rect 25494 4864 25510 4928
rect 25574 4864 25580 4928
rect 25264 4863 25580 4864
rect 29200 4768 30000 4888
rect 7894 4384 8210 4385
rect 7894 4320 7900 4384
rect 7964 4320 7980 4384
rect 8044 4320 8060 4384
rect 8124 4320 8140 4384
rect 8204 4320 8210 4384
rect 7894 4319 8210 4320
rect 14842 4384 15158 4385
rect 14842 4320 14848 4384
rect 14912 4320 14928 4384
rect 14992 4320 15008 4384
rect 15072 4320 15088 4384
rect 15152 4320 15158 4384
rect 14842 4319 15158 4320
rect 21790 4384 22106 4385
rect 21790 4320 21796 4384
rect 21860 4320 21876 4384
rect 21940 4320 21956 4384
rect 22020 4320 22036 4384
rect 22100 4320 22106 4384
rect 21790 4319 22106 4320
rect 0 4088 800 4208
rect 29200 4088 30000 4208
rect 4420 3840 4736 3841
rect 4420 3776 4426 3840
rect 4490 3776 4506 3840
rect 4570 3776 4586 3840
rect 4650 3776 4666 3840
rect 4730 3776 4736 3840
rect 4420 3775 4736 3776
rect 11368 3840 11684 3841
rect 11368 3776 11374 3840
rect 11438 3776 11454 3840
rect 11518 3776 11534 3840
rect 11598 3776 11614 3840
rect 11678 3776 11684 3840
rect 11368 3775 11684 3776
rect 18316 3840 18632 3841
rect 18316 3776 18322 3840
rect 18386 3776 18402 3840
rect 18466 3776 18482 3840
rect 18546 3776 18562 3840
rect 18626 3776 18632 3840
rect 18316 3775 18632 3776
rect 25264 3840 25580 3841
rect 25264 3776 25270 3840
rect 25334 3776 25350 3840
rect 25414 3776 25430 3840
rect 25494 3776 25510 3840
rect 25574 3776 25580 3840
rect 25264 3775 25580 3776
rect 0 3408 800 3528
rect 7894 3296 8210 3297
rect 7894 3232 7900 3296
rect 7964 3232 7980 3296
rect 8044 3232 8060 3296
rect 8124 3232 8140 3296
rect 8204 3232 8210 3296
rect 7894 3231 8210 3232
rect 14842 3296 15158 3297
rect 14842 3232 14848 3296
rect 14912 3232 14928 3296
rect 14992 3232 15008 3296
rect 15072 3232 15088 3296
rect 15152 3232 15158 3296
rect 14842 3231 15158 3232
rect 21790 3296 22106 3297
rect 21790 3232 21796 3296
rect 21860 3232 21876 3296
rect 21940 3232 21956 3296
rect 22020 3232 22036 3296
rect 22100 3232 22106 3296
rect 21790 3231 22106 3232
rect 0 2728 800 2848
rect 4420 2752 4736 2753
rect 4420 2688 4426 2752
rect 4490 2688 4506 2752
rect 4570 2688 4586 2752
rect 4650 2688 4666 2752
rect 4730 2688 4736 2752
rect 4420 2687 4736 2688
rect 11368 2752 11684 2753
rect 11368 2688 11374 2752
rect 11438 2688 11454 2752
rect 11518 2688 11534 2752
rect 11598 2688 11614 2752
rect 11678 2688 11684 2752
rect 11368 2687 11684 2688
rect 18316 2752 18632 2753
rect 18316 2688 18322 2752
rect 18386 2688 18402 2752
rect 18466 2688 18482 2752
rect 18546 2688 18562 2752
rect 18626 2688 18632 2752
rect 18316 2687 18632 2688
rect 25264 2752 25580 2753
rect 25264 2688 25270 2752
rect 25334 2688 25350 2752
rect 25414 2688 25430 2752
rect 25494 2688 25510 2752
rect 25574 2688 25580 2752
rect 29200 2728 30000 2848
rect 25264 2687 25580 2688
rect 7894 2208 8210 2209
rect 7894 2144 7900 2208
rect 7964 2144 7980 2208
rect 8044 2144 8060 2208
rect 8124 2144 8140 2208
rect 8204 2144 8210 2208
rect 7894 2143 8210 2144
rect 14842 2208 15158 2209
rect 14842 2144 14848 2208
rect 14912 2144 14928 2208
rect 14992 2144 15008 2208
rect 15072 2144 15088 2208
rect 15152 2144 15158 2208
rect 14842 2143 15158 2144
rect 21790 2208 22106 2209
rect 21790 2144 21796 2208
rect 21860 2144 21876 2208
rect 21940 2144 21956 2208
rect 22020 2144 22036 2208
rect 22100 2144 22106 2208
rect 21790 2143 22106 2144
rect 29200 2048 30000 2168
rect 0 1368 800 1488
rect 29200 1368 30000 1488
rect 0 688 800 808
rect 29200 8 30000 128
<< via3 >>
rect 4426 27772 4490 27776
rect 4426 27716 4430 27772
rect 4430 27716 4486 27772
rect 4486 27716 4490 27772
rect 4426 27712 4490 27716
rect 4506 27772 4570 27776
rect 4506 27716 4510 27772
rect 4510 27716 4566 27772
rect 4566 27716 4570 27772
rect 4506 27712 4570 27716
rect 4586 27772 4650 27776
rect 4586 27716 4590 27772
rect 4590 27716 4646 27772
rect 4646 27716 4650 27772
rect 4586 27712 4650 27716
rect 4666 27772 4730 27776
rect 4666 27716 4670 27772
rect 4670 27716 4726 27772
rect 4726 27716 4730 27772
rect 4666 27712 4730 27716
rect 11374 27772 11438 27776
rect 11374 27716 11378 27772
rect 11378 27716 11434 27772
rect 11434 27716 11438 27772
rect 11374 27712 11438 27716
rect 11454 27772 11518 27776
rect 11454 27716 11458 27772
rect 11458 27716 11514 27772
rect 11514 27716 11518 27772
rect 11454 27712 11518 27716
rect 11534 27772 11598 27776
rect 11534 27716 11538 27772
rect 11538 27716 11594 27772
rect 11594 27716 11598 27772
rect 11534 27712 11598 27716
rect 11614 27772 11678 27776
rect 11614 27716 11618 27772
rect 11618 27716 11674 27772
rect 11674 27716 11678 27772
rect 11614 27712 11678 27716
rect 18322 27772 18386 27776
rect 18322 27716 18326 27772
rect 18326 27716 18382 27772
rect 18382 27716 18386 27772
rect 18322 27712 18386 27716
rect 18402 27772 18466 27776
rect 18402 27716 18406 27772
rect 18406 27716 18462 27772
rect 18462 27716 18466 27772
rect 18402 27712 18466 27716
rect 18482 27772 18546 27776
rect 18482 27716 18486 27772
rect 18486 27716 18542 27772
rect 18542 27716 18546 27772
rect 18482 27712 18546 27716
rect 18562 27772 18626 27776
rect 18562 27716 18566 27772
rect 18566 27716 18622 27772
rect 18622 27716 18626 27772
rect 18562 27712 18626 27716
rect 25270 27772 25334 27776
rect 25270 27716 25274 27772
rect 25274 27716 25330 27772
rect 25330 27716 25334 27772
rect 25270 27712 25334 27716
rect 25350 27772 25414 27776
rect 25350 27716 25354 27772
rect 25354 27716 25410 27772
rect 25410 27716 25414 27772
rect 25350 27712 25414 27716
rect 25430 27772 25494 27776
rect 25430 27716 25434 27772
rect 25434 27716 25490 27772
rect 25490 27716 25494 27772
rect 25430 27712 25494 27716
rect 25510 27772 25574 27776
rect 25510 27716 25514 27772
rect 25514 27716 25570 27772
rect 25570 27716 25574 27772
rect 25510 27712 25574 27716
rect 7900 27228 7964 27232
rect 7900 27172 7904 27228
rect 7904 27172 7960 27228
rect 7960 27172 7964 27228
rect 7900 27168 7964 27172
rect 7980 27228 8044 27232
rect 7980 27172 7984 27228
rect 7984 27172 8040 27228
rect 8040 27172 8044 27228
rect 7980 27168 8044 27172
rect 8060 27228 8124 27232
rect 8060 27172 8064 27228
rect 8064 27172 8120 27228
rect 8120 27172 8124 27228
rect 8060 27168 8124 27172
rect 8140 27228 8204 27232
rect 8140 27172 8144 27228
rect 8144 27172 8200 27228
rect 8200 27172 8204 27228
rect 8140 27168 8204 27172
rect 14848 27228 14912 27232
rect 14848 27172 14852 27228
rect 14852 27172 14908 27228
rect 14908 27172 14912 27228
rect 14848 27168 14912 27172
rect 14928 27228 14992 27232
rect 14928 27172 14932 27228
rect 14932 27172 14988 27228
rect 14988 27172 14992 27228
rect 14928 27168 14992 27172
rect 15008 27228 15072 27232
rect 15008 27172 15012 27228
rect 15012 27172 15068 27228
rect 15068 27172 15072 27228
rect 15008 27168 15072 27172
rect 15088 27228 15152 27232
rect 15088 27172 15092 27228
rect 15092 27172 15148 27228
rect 15148 27172 15152 27228
rect 15088 27168 15152 27172
rect 21796 27228 21860 27232
rect 21796 27172 21800 27228
rect 21800 27172 21856 27228
rect 21856 27172 21860 27228
rect 21796 27168 21860 27172
rect 21876 27228 21940 27232
rect 21876 27172 21880 27228
rect 21880 27172 21936 27228
rect 21936 27172 21940 27228
rect 21876 27168 21940 27172
rect 21956 27228 22020 27232
rect 21956 27172 21960 27228
rect 21960 27172 22016 27228
rect 22016 27172 22020 27228
rect 21956 27168 22020 27172
rect 22036 27228 22100 27232
rect 22036 27172 22040 27228
rect 22040 27172 22096 27228
rect 22096 27172 22100 27228
rect 22036 27168 22100 27172
rect 4426 26684 4490 26688
rect 4426 26628 4430 26684
rect 4430 26628 4486 26684
rect 4486 26628 4490 26684
rect 4426 26624 4490 26628
rect 4506 26684 4570 26688
rect 4506 26628 4510 26684
rect 4510 26628 4566 26684
rect 4566 26628 4570 26684
rect 4506 26624 4570 26628
rect 4586 26684 4650 26688
rect 4586 26628 4590 26684
rect 4590 26628 4646 26684
rect 4646 26628 4650 26684
rect 4586 26624 4650 26628
rect 4666 26684 4730 26688
rect 4666 26628 4670 26684
rect 4670 26628 4726 26684
rect 4726 26628 4730 26684
rect 4666 26624 4730 26628
rect 11374 26684 11438 26688
rect 11374 26628 11378 26684
rect 11378 26628 11434 26684
rect 11434 26628 11438 26684
rect 11374 26624 11438 26628
rect 11454 26684 11518 26688
rect 11454 26628 11458 26684
rect 11458 26628 11514 26684
rect 11514 26628 11518 26684
rect 11454 26624 11518 26628
rect 11534 26684 11598 26688
rect 11534 26628 11538 26684
rect 11538 26628 11594 26684
rect 11594 26628 11598 26684
rect 11534 26624 11598 26628
rect 11614 26684 11678 26688
rect 11614 26628 11618 26684
rect 11618 26628 11674 26684
rect 11674 26628 11678 26684
rect 11614 26624 11678 26628
rect 18322 26684 18386 26688
rect 18322 26628 18326 26684
rect 18326 26628 18382 26684
rect 18382 26628 18386 26684
rect 18322 26624 18386 26628
rect 18402 26684 18466 26688
rect 18402 26628 18406 26684
rect 18406 26628 18462 26684
rect 18462 26628 18466 26684
rect 18402 26624 18466 26628
rect 18482 26684 18546 26688
rect 18482 26628 18486 26684
rect 18486 26628 18542 26684
rect 18542 26628 18546 26684
rect 18482 26624 18546 26628
rect 18562 26684 18626 26688
rect 18562 26628 18566 26684
rect 18566 26628 18622 26684
rect 18622 26628 18626 26684
rect 18562 26624 18626 26628
rect 25270 26684 25334 26688
rect 25270 26628 25274 26684
rect 25274 26628 25330 26684
rect 25330 26628 25334 26684
rect 25270 26624 25334 26628
rect 25350 26684 25414 26688
rect 25350 26628 25354 26684
rect 25354 26628 25410 26684
rect 25410 26628 25414 26684
rect 25350 26624 25414 26628
rect 25430 26684 25494 26688
rect 25430 26628 25434 26684
rect 25434 26628 25490 26684
rect 25490 26628 25494 26684
rect 25430 26624 25494 26628
rect 25510 26684 25574 26688
rect 25510 26628 25514 26684
rect 25514 26628 25570 26684
rect 25570 26628 25574 26684
rect 25510 26624 25574 26628
rect 7900 26140 7964 26144
rect 7900 26084 7904 26140
rect 7904 26084 7960 26140
rect 7960 26084 7964 26140
rect 7900 26080 7964 26084
rect 7980 26140 8044 26144
rect 7980 26084 7984 26140
rect 7984 26084 8040 26140
rect 8040 26084 8044 26140
rect 7980 26080 8044 26084
rect 8060 26140 8124 26144
rect 8060 26084 8064 26140
rect 8064 26084 8120 26140
rect 8120 26084 8124 26140
rect 8060 26080 8124 26084
rect 8140 26140 8204 26144
rect 8140 26084 8144 26140
rect 8144 26084 8200 26140
rect 8200 26084 8204 26140
rect 8140 26080 8204 26084
rect 14848 26140 14912 26144
rect 14848 26084 14852 26140
rect 14852 26084 14908 26140
rect 14908 26084 14912 26140
rect 14848 26080 14912 26084
rect 14928 26140 14992 26144
rect 14928 26084 14932 26140
rect 14932 26084 14988 26140
rect 14988 26084 14992 26140
rect 14928 26080 14992 26084
rect 15008 26140 15072 26144
rect 15008 26084 15012 26140
rect 15012 26084 15068 26140
rect 15068 26084 15072 26140
rect 15008 26080 15072 26084
rect 15088 26140 15152 26144
rect 15088 26084 15092 26140
rect 15092 26084 15148 26140
rect 15148 26084 15152 26140
rect 15088 26080 15152 26084
rect 21796 26140 21860 26144
rect 21796 26084 21800 26140
rect 21800 26084 21856 26140
rect 21856 26084 21860 26140
rect 21796 26080 21860 26084
rect 21876 26140 21940 26144
rect 21876 26084 21880 26140
rect 21880 26084 21936 26140
rect 21936 26084 21940 26140
rect 21876 26080 21940 26084
rect 21956 26140 22020 26144
rect 21956 26084 21960 26140
rect 21960 26084 22016 26140
rect 22016 26084 22020 26140
rect 21956 26080 22020 26084
rect 22036 26140 22100 26144
rect 22036 26084 22040 26140
rect 22040 26084 22096 26140
rect 22096 26084 22100 26140
rect 22036 26080 22100 26084
rect 4426 25596 4490 25600
rect 4426 25540 4430 25596
rect 4430 25540 4486 25596
rect 4486 25540 4490 25596
rect 4426 25536 4490 25540
rect 4506 25596 4570 25600
rect 4506 25540 4510 25596
rect 4510 25540 4566 25596
rect 4566 25540 4570 25596
rect 4506 25536 4570 25540
rect 4586 25596 4650 25600
rect 4586 25540 4590 25596
rect 4590 25540 4646 25596
rect 4646 25540 4650 25596
rect 4586 25536 4650 25540
rect 4666 25596 4730 25600
rect 4666 25540 4670 25596
rect 4670 25540 4726 25596
rect 4726 25540 4730 25596
rect 4666 25536 4730 25540
rect 11374 25596 11438 25600
rect 11374 25540 11378 25596
rect 11378 25540 11434 25596
rect 11434 25540 11438 25596
rect 11374 25536 11438 25540
rect 11454 25596 11518 25600
rect 11454 25540 11458 25596
rect 11458 25540 11514 25596
rect 11514 25540 11518 25596
rect 11454 25536 11518 25540
rect 11534 25596 11598 25600
rect 11534 25540 11538 25596
rect 11538 25540 11594 25596
rect 11594 25540 11598 25596
rect 11534 25536 11598 25540
rect 11614 25596 11678 25600
rect 11614 25540 11618 25596
rect 11618 25540 11674 25596
rect 11674 25540 11678 25596
rect 11614 25536 11678 25540
rect 18322 25596 18386 25600
rect 18322 25540 18326 25596
rect 18326 25540 18382 25596
rect 18382 25540 18386 25596
rect 18322 25536 18386 25540
rect 18402 25596 18466 25600
rect 18402 25540 18406 25596
rect 18406 25540 18462 25596
rect 18462 25540 18466 25596
rect 18402 25536 18466 25540
rect 18482 25596 18546 25600
rect 18482 25540 18486 25596
rect 18486 25540 18542 25596
rect 18542 25540 18546 25596
rect 18482 25536 18546 25540
rect 18562 25596 18626 25600
rect 18562 25540 18566 25596
rect 18566 25540 18622 25596
rect 18622 25540 18626 25596
rect 18562 25536 18626 25540
rect 25270 25596 25334 25600
rect 25270 25540 25274 25596
rect 25274 25540 25330 25596
rect 25330 25540 25334 25596
rect 25270 25536 25334 25540
rect 25350 25596 25414 25600
rect 25350 25540 25354 25596
rect 25354 25540 25410 25596
rect 25410 25540 25414 25596
rect 25350 25536 25414 25540
rect 25430 25596 25494 25600
rect 25430 25540 25434 25596
rect 25434 25540 25490 25596
rect 25490 25540 25494 25596
rect 25430 25536 25494 25540
rect 25510 25596 25574 25600
rect 25510 25540 25514 25596
rect 25514 25540 25570 25596
rect 25570 25540 25574 25596
rect 25510 25536 25574 25540
rect 7900 25052 7964 25056
rect 7900 24996 7904 25052
rect 7904 24996 7960 25052
rect 7960 24996 7964 25052
rect 7900 24992 7964 24996
rect 7980 25052 8044 25056
rect 7980 24996 7984 25052
rect 7984 24996 8040 25052
rect 8040 24996 8044 25052
rect 7980 24992 8044 24996
rect 8060 25052 8124 25056
rect 8060 24996 8064 25052
rect 8064 24996 8120 25052
rect 8120 24996 8124 25052
rect 8060 24992 8124 24996
rect 8140 25052 8204 25056
rect 8140 24996 8144 25052
rect 8144 24996 8200 25052
rect 8200 24996 8204 25052
rect 8140 24992 8204 24996
rect 14848 25052 14912 25056
rect 14848 24996 14852 25052
rect 14852 24996 14908 25052
rect 14908 24996 14912 25052
rect 14848 24992 14912 24996
rect 14928 25052 14992 25056
rect 14928 24996 14932 25052
rect 14932 24996 14988 25052
rect 14988 24996 14992 25052
rect 14928 24992 14992 24996
rect 15008 25052 15072 25056
rect 15008 24996 15012 25052
rect 15012 24996 15068 25052
rect 15068 24996 15072 25052
rect 15008 24992 15072 24996
rect 15088 25052 15152 25056
rect 15088 24996 15092 25052
rect 15092 24996 15148 25052
rect 15148 24996 15152 25052
rect 15088 24992 15152 24996
rect 21796 25052 21860 25056
rect 21796 24996 21800 25052
rect 21800 24996 21856 25052
rect 21856 24996 21860 25052
rect 21796 24992 21860 24996
rect 21876 25052 21940 25056
rect 21876 24996 21880 25052
rect 21880 24996 21936 25052
rect 21936 24996 21940 25052
rect 21876 24992 21940 24996
rect 21956 25052 22020 25056
rect 21956 24996 21960 25052
rect 21960 24996 22016 25052
rect 22016 24996 22020 25052
rect 21956 24992 22020 24996
rect 22036 25052 22100 25056
rect 22036 24996 22040 25052
rect 22040 24996 22096 25052
rect 22096 24996 22100 25052
rect 22036 24992 22100 24996
rect 4426 24508 4490 24512
rect 4426 24452 4430 24508
rect 4430 24452 4486 24508
rect 4486 24452 4490 24508
rect 4426 24448 4490 24452
rect 4506 24508 4570 24512
rect 4506 24452 4510 24508
rect 4510 24452 4566 24508
rect 4566 24452 4570 24508
rect 4506 24448 4570 24452
rect 4586 24508 4650 24512
rect 4586 24452 4590 24508
rect 4590 24452 4646 24508
rect 4646 24452 4650 24508
rect 4586 24448 4650 24452
rect 4666 24508 4730 24512
rect 4666 24452 4670 24508
rect 4670 24452 4726 24508
rect 4726 24452 4730 24508
rect 4666 24448 4730 24452
rect 11374 24508 11438 24512
rect 11374 24452 11378 24508
rect 11378 24452 11434 24508
rect 11434 24452 11438 24508
rect 11374 24448 11438 24452
rect 11454 24508 11518 24512
rect 11454 24452 11458 24508
rect 11458 24452 11514 24508
rect 11514 24452 11518 24508
rect 11454 24448 11518 24452
rect 11534 24508 11598 24512
rect 11534 24452 11538 24508
rect 11538 24452 11594 24508
rect 11594 24452 11598 24508
rect 11534 24448 11598 24452
rect 11614 24508 11678 24512
rect 11614 24452 11618 24508
rect 11618 24452 11674 24508
rect 11674 24452 11678 24508
rect 11614 24448 11678 24452
rect 18322 24508 18386 24512
rect 18322 24452 18326 24508
rect 18326 24452 18382 24508
rect 18382 24452 18386 24508
rect 18322 24448 18386 24452
rect 18402 24508 18466 24512
rect 18402 24452 18406 24508
rect 18406 24452 18462 24508
rect 18462 24452 18466 24508
rect 18402 24448 18466 24452
rect 18482 24508 18546 24512
rect 18482 24452 18486 24508
rect 18486 24452 18542 24508
rect 18542 24452 18546 24508
rect 18482 24448 18546 24452
rect 18562 24508 18626 24512
rect 18562 24452 18566 24508
rect 18566 24452 18622 24508
rect 18622 24452 18626 24508
rect 18562 24448 18626 24452
rect 25270 24508 25334 24512
rect 25270 24452 25274 24508
rect 25274 24452 25330 24508
rect 25330 24452 25334 24508
rect 25270 24448 25334 24452
rect 25350 24508 25414 24512
rect 25350 24452 25354 24508
rect 25354 24452 25410 24508
rect 25410 24452 25414 24508
rect 25350 24448 25414 24452
rect 25430 24508 25494 24512
rect 25430 24452 25434 24508
rect 25434 24452 25490 24508
rect 25490 24452 25494 24508
rect 25430 24448 25494 24452
rect 25510 24508 25574 24512
rect 25510 24452 25514 24508
rect 25514 24452 25570 24508
rect 25570 24452 25574 24508
rect 25510 24448 25574 24452
rect 7900 23964 7964 23968
rect 7900 23908 7904 23964
rect 7904 23908 7960 23964
rect 7960 23908 7964 23964
rect 7900 23904 7964 23908
rect 7980 23964 8044 23968
rect 7980 23908 7984 23964
rect 7984 23908 8040 23964
rect 8040 23908 8044 23964
rect 7980 23904 8044 23908
rect 8060 23964 8124 23968
rect 8060 23908 8064 23964
rect 8064 23908 8120 23964
rect 8120 23908 8124 23964
rect 8060 23904 8124 23908
rect 8140 23964 8204 23968
rect 8140 23908 8144 23964
rect 8144 23908 8200 23964
rect 8200 23908 8204 23964
rect 8140 23904 8204 23908
rect 14848 23964 14912 23968
rect 14848 23908 14852 23964
rect 14852 23908 14908 23964
rect 14908 23908 14912 23964
rect 14848 23904 14912 23908
rect 14928 23964 14992 23968
rect 14928 23908 14932 23964
rect 14932 23908 14988 23964
rect 14988 23908 14992 23964
rect 14928 23904 14992 23908
rect 15008 23964 15072 23968
rect 15008 23908 15012 23964
rect 15012 23908 15068 23964
rect 15068 23908 15072 23964
rect 15008 23904 15072 23908
rect 15088 23964 15152 23968
rect 15088 23908 15092 23964
rect 15092 23908 15148 23964
rect 15148 23908 15152 23964
rect 15088 23904 15152 23908
rect 21796 23964 21860 23968
rect 21796 23908 21800 23964
rect 21800 23908 21856 23964
rect 21856 23908 21860 23964
rect 21796 23904 21860 23908
rect 21876 23964 21940 23968
rect 21876 23908 21880 23964
rect 21880 23908 21936 23964
rect 21936 23908 21940 23964
rect 21876 23904 21940 23908
rect 21956 23964 22020 23968
rect 21956 23908 21960 23964
rect 21960 23908 22016 23964
rect 22016 23908 22020 23964
rect 21956 23904 22020 23908
rect 22036 23964 22100 23968
rect 22036 23908 22040 23964
rect 22040 23908 22096 23964
rect 22096 23908 22100 23964
rect 22036 23904 22100 23908
rect 4426 23420 4490 23424
rect 4426 23364 4430 23420
rect 4430 23364 4486 23420
rect 4486 23364 4490 23420
rect 4426 23360 4490 23364
rect 4506 23420 4570 23424
rect 4506 23364 4510 23420
rect 4510 23364 4566 23420
rect 4566 23364 4570 23420
rect 4506 23360 4570 23364
rect 4586 23420 4650 23424
rect 4586 23364 4590 23420
rect 4590 23364 4646 23420
rect 4646 23364 4650 23420
rect 4586 23360 4650 23364
rect 4666 23420 4730 23424
rect 4666 23364 4670 23420
rect 4670 23364 4726 23420
rect 4726 23364 4730 23420
rect 4666 23360 4730 23364
rect 11374 23420 11438 23424
rect 11374 23364 11378 23420
rect 11378 23364 11434 23420
rect 11434 23364 11438 23420
rect 11374 23360 11438 23364
rect 11454 23420 11518 23424
rect 11454 23364 11458 23420
rect 11458 23364 11514 23420
rect 11514 23364 11518 23420
rect 11454 23360 11518 23364
rect 11534 23420 11598 23424
rect 11534 23364 11538 23420
rect 11538 23364 11594 23420
rect 11594 23364 11598 23420
rect 11534 23360 11598 23364
rect 11614 23420 11678 23424
rect 11614 23364 11618 23420
rect 11618 23364 11674 23420
rect 11674 23364 11678 23420
rect 11614 23360 11678 23364
rect 18322 23420 18386 23424
rect 18322 23364 18326 23420
rect 18326 23364 18382 23420
rect 18382 23364 18386 23420
rect 18322 23360 18386 23364
rect 18402 23420 18466 23424
rect 18402 23364 18406 23420
rect 18406 23364 18462 23420
rect 18462 23364 18466 23420
rect 18402 23360 18466 23364
rect 18482 23420 18546 23424
rect 18482 23364 18486 23420
rect 18486 23364 18542 23420
rect 18542 23364 18546 23420
rect 18482 23360 18546 23364
rect 18562 23420 18626 23424
rect 18562 23364 18566 23420
rect 18566 23364 18622 23420
rect 18622 23364 18626 23420
rect 18562 23360 18626 23364
rect 25270 23420 25334 23424
rect 25270 23364 25274 23420
rect 25274 23364 25330 23420
rect 25330 23364 25334 23420
rect 25270 23360 25334 23364
rect 25350 23420 25414 23424
rect 25350 23364 25354 23420
rect 25354 23364 25410 23420
rect 25410 23364 25414 23420
rect 25350 23360 25414 23364
rect 25430 23420 25494 23424
rect 25430 23364 25434 23420
rect 25434 23364 25490 23420
rect 25490 23364 25494 23420
rect 25430 23360 25494 23364
rect 25510 23420 25574 23424
rect 25510 23364 25514 23420
rect 25514 23364 25570 23420
rect 25570 23364 25574 23420
rect 25510 23360 25574 23364
rect 7900 22876 7964 22880
rect 7900 22820 7904 22876
rect 7904 22820 7960 22876
rect 7960 22820 7964 22876
rect 7900 22816 7964 22820
rect 7980 22876 8044 22880
rect 7980 22820 7984 22876
rect 7984 22820 8040 22876
rect 8040 22820 8044 22876
rect 7980 22816 8044 22820
rect 8060 22876 8124 22880
rect 8060 22820 8064 22876
rect 8064 22820 8120 22876
rect 8120 22820 8124 22876
rect 8060 22816 8124 22820
rect 8140 22876 8204 22880
rect 8140 22820 8144 22876
rect 8144 22820 8200 22876
rect 8200 22820 8204 22876
rect 8140 22816 8204 22820
rect 14848 22876 14912 22880
rect 14848 22820 14852 22876
rect 14852 22820 14908 22876
rect 14908 22820 14912 22876
rect 14848 22816 14912 22820
rect 14928 22876 14992 22880
rect 14928 22820 14932 22876
rect 14932 22820 14988 22876
rect 14988 22820 14992 22876
rect 14928 22816 14992 22820
rect 15008 22876 15072 22880
rect 15008 22820 15012 22876
rect 15012 22820 15068 22876
rect 15068 22820 15072 22876
rect 15008 22816 15072 22820
rect 15088 22876 15152 22880
rect 15088 22820 15092 22876
rect 15092 22820 15148 22876
rect 15148 22820 15152 22876
rect 15088 22816 15152 22820
rect 21796 22876 21860 22880
rect 21796 22820 21800 22876
rect 21800 22820 21856 22876
rect 21856 22820 21860 22876
rect 21796 22816 21860 22820
rect 21876 22876 21940 22880
rect 21876 22820 21880 22876
rect 21880 22820 21936 22876
rect 21936 22820 21940 22876
rect 21876 22816 21940 22820
rect 21956 22876 22020 22880
rect 21956 22820 21960 22876
rect 21960 22820 22016 22876
rect 22016 22820 22020 22876
rect 21956 22816 22020 22820
rect 22036 22876 22100 22880
rect 22036 22820 22040 22876
rect 22040 22820 22096 22876
rect 22096 22820 22100 22876
rect 22036 22816 22100 22820
rect 4426 22332 4490 22336
rect 4426 22276 4430 22332
rect 4430 22276 4486 22332
rect 4486 22276 4490 22332
rect 4426 22272 4490 22276
rect 4506 22332 4570 22336
rect 4506 22276 4510 22332
rect 4510 22276 4566 22332
rect 4566 22276 4570 22332
rect 4506 22272 4570 22276
rect 4586 22332 4650 22336
rect 4586 22276 4590 22332
rect 4590 22276 4646 22332
rect 4646 22276 4650 22332
rect 4586 22272 4650 22276
rect 4666 22332 4730 22336
rect 4666 22276 4670 22332
rect 4670 22276 4726 22332
rect 4726 22276 4730 22332
rect 4666 22272 4730 22276
rect 11374 22332 11438 22336
rect 11374 22276 11378 22332
rect 11378 22276 11434 22332
rect 11434 22276 11438 22332
rect 11374 22272 11438 22276
rect 11454 22332 11518 22336
rect 11454 22276 11458 22332
rect 11458 22276 11514 22332
rect 11514 22276 11518 22332
rect 11454 22272 11518 22276
rect 11534 22332 11598 22336
rect 11534 22276 11538 22332
rect 11538 22276 11594 22332
rect 11594 22276 11598 22332
rect 11534 22272 11598 22276
rect 11614 22332 11678 22336
rect 11614 22276 11618 22332
rect 11618 22276 11674 22332
rect 11674 22276 11678 22332
rect 11614 22272 11678 22276
rect 18322 22332 18386 22336
rect 18322 22276 18326 22332
rect 18326 22276 18382 22332
rect 18382 22276 18386 22332
rect 18322 22272 18386 22276
rect 18402 22332 18466 22336
rect 18402 22276 18406 22332
rect 18406 22276 18462 22332
rect 18462 22276 18466 22332
rect 18402 22272 18466 22276
rect 18482 22332 18546 22336
rect 18482 22276 18486 22332
rect 18486 22276 18542 22332
rect 18542 22276 18546 22332
rect 18482 22272 18546 22276
rect 18562 22332 18626 22336
rect 18562 22276 18566 22332
rect 18566 22276 18622 22332
rect 18622 22276 18626 22332
rect 18562 22272 18626 22276
rect 25270 22332 25334 22336
rect 25270 22276 25274 22332
rect 25274 22276 25330 22332
rect 25330 22276 25334 22332
rect 25270 22272 25334 22276
rect 25350 22332 25414 22336
rect 25350 22276 25354 22332
rect 25354 22276 25410 22332
rect 25410 22276 25414 22332
rect 25350 22272 25414 22276
rect 25430 22332 25494 22336
rect 25430 22276 25434 22332
rect 25434 22276 25490 22332
rect 25490 22276 25494 22332
rect 25430 22272 25494 22276
rect 25510 22332 25574 22336
rect 25510 22276 25514 22332
rect 25514 22276 25570 22332
rect 25570 22276 25574 22332
rect 25510 22272 25574 22276
rect 7900 21788 7964 21792
rect 7900 21732 7904 21788
rect 7904 21732 7960 21788
rect 7960 21732 7964 21788
rect 7900 21728 7964 21732
rect 7980 21788 8044 21792
rect 7980 21732 7984 21788
rect 7984 21732 8040 21788
rect 8040 21732 8044 21788
rect 7980 21728 8044 21732
rect 8060 21788 8124 21792
rect 8060 21732 8064 21788
rect 8064 21732 8120 21788
rect 8120 21732 8124 21788
rect 8060 21728 8124 21732
rect 8140 21788 8204 21792
rect 8140 21732 8144 21788
rect 8144 21732 8200 21788
rect 8200 21732 8204 21788
rect 8140 21728 8204 21732
rect 14848 21788 14912 21792
rect 14848 21732 14852 21788
rect 14852 21732 14908 21788
rect 14908 21732 14912 21788
rect 14848 21728 14912 21732
rect 14928 21788 14992 21792
rect 14928 21732 14932 21788
rect 14932 21732 14988 21788
rect 14988 21732 14992 21788
rect 14928 21728 14992 21732
rect 15008 21788 15072 21792
rect 15008 21732 15012 21788
rect 15012 21732 15068 21788
rect 15068 21732 15072 21788
rect 15008 21728 15072 21732
rect 15088 21788 15152 21792
rect 15088 21732 15092 21788
rect 15092 21732 15148 21788
rect 15148 21732 15152 21788
rect 15088 21728 15152 21732
rect 21796 21788 21860 21792
rect 21796 21732 21800 21788
rect 21800 21732 21856 21788
rect 21856 21732 21860 21788
rect 21796 21728 21860 21732
rect 21876 21788 21940 21792
rect 21876 21732 21880 21788
rect 21880 21732 21936 21788
rect 21936 21732 21940 21788
rect 21876 21728 21940 21732
rect 21956 21788 22020 21792
rect 21956 21732 21960 21788
rect 21960 21732 22016 21788
rect 22016 21732 22020 21788
rect 21956 21728 22020 21732
rect 22036 21788 22100 21792
rect 22036 21732 22040 21788
rect 22040 21732 22096 21788
rect 22096 21732 22100 21788
rect 22036 21728 22100 21732
rect 4426 21244 4490 21248
rect 4426 21188 4430 21244
rect 4430 21188 4486 21244
rect 4486 21188 4490 21244
rect 4426 21184 4490 21188
rect 4506 21244 4570 21248
rect 4506 21188 4510 21244
rect 4510 21188 4566 21244
rect 4566 21188 4570 21244
rect 4506 21184 4570 21188
rect 4586 21244 4650 21248
rect 4586 21188 4590 21244
rect 4590 21188 4646 21244
rect 4646 21188 4650 21244
rect 4586 21184 4650 21188
rect 4666 21244 4730 21248
rect 4666 21188 4670 21244
rect 4670 21188 4726 21244
rect 4726 21188 4730 21244
rect 4666 21184 4730 21188
rect 11374 21244 11438 21248
rect 11374 21188 11378 21244
rect 11378 21188 11434 21244
rect 11434 21188 11438 21244
rect 11374 21184 11438 21188
rect 11454 21244 11518 21248
rect 11454 21188 11458 21244
rect 11458 21188 11514 21244
rect 11514 21188 11518 21244
rect 11454 21184 11518 21188
rect 11534 21244 11598 21248
rect 11534 21188 11538 21244
rect 11538 21188 11594 21244
rect 11594 21188 11598 21244
rect 11534 21184 11598 21188
rect 11614 21244 11678 21248
rect 11614 21188 11618 21244
rect 11618 21188 11674 21244
rect 11674 21188 11678 21244
rect 11614 21184 11678 21188
rect 18322 21244 18386 21248
rect 18322 21188 18326 21244
rect 18326 21188 18382 21244
rect 18382 21188 18386 21244
rect 18322 21184 18386 21188
rect 18402 21244 18466 21248
rect 18402 21188 18406 21244
rect 18406 21188 18462 21244
rect 18462 21188 18466 21244
rect 18402 21184 18466 21188
rect 18482 21244 18546 21248
rect 18482 21188 18486 21244
rect 18486 21188 18542 21244
rect 18542 21188 18546 21244
rect 18482 21184 18546 21188
rect 18562 21244 18626 21248
rect 18562 21188 18566 21244
rect 18566 21188 18622 21244
rect 18622 21188 18626 21244
rect 18562 21184 18626 21188
rect 25270 21244 25334 21248
rect 25270 21188 25274 21244
rect 25274 21188 25330 21244
rect 25330 21188 25334 21244
rect 25270 21184 25334 21188
rect 25350 21244 25414 21248
rect 25350 21188 25354 21244
rect 25354 21188 25410 21244
rect 25410 21188 25414 21244
rect 25350 21184 25414 21188
rect 25430 21244 25494 21248
rect 25430 21188 25434 21244
rect 25434 21188 25490 21244
rect 25490 21188 25494 21244
rect 25430 21184 25494 21188
rect 25510 21244 25574 21248
rect 25510 21188 25514 21244
rect 25514 21188 25570 21244
rect 25570 21188 25574 21244
rect 25510 21184 25574 21188
rect 7900 20700 7964 20704
rect 7900 20644 7904 20700
rect 7904 20644 7960 20700
rect 7960 20644 7964 20700
rect 7900 20640 7964 20644
rect 7980 20700 8044 20704
rect 7980 20644 7984 20700
rect 7984 20644 8040 20700
rect 8040 20644 8044 20700
rect 7980 20640 8044 20644
rect 8060 20700 8124 20704
rect 8060 20644 8064 20700
rect 8064 20644 8120 20700
rect 8120 20644 8124 20700
rect 8060 20640 8124 20644
rect 8140 20700 8204 20704
rect 8140 20644 8144 20700
rect 8144 20644 8200 20700
rect 8200 20644 8204 20700
rect 8140 20640 8204 20644
rect 14848 20700 14912 20704
rect 14848 20644 14852 20700
rect 14852 20644 14908 20700
rect 14908 20644 14912 20700
rect 14848 20640 14912 20644
rect 14928 20700 14992 20704
rect 14928 20644 14932 20700
rect 14932 20644 14988 20700
rect 14988 20644 14992 20700
rect 14928 20640 14992 20644
rect 15008 20700 15072 20704
rect 15008 20644 15012 20700
rect 15012 20644 15068 20700
rect 15068 20644 15072 20700
rect 15008 20640 15072 20644
rect 15088 20700 15152 20704
rect 15088 20644 15092 20700
rect 15092 20644 15148 20700
rect 15148 20644 15152 20700
rect 15088 20640 15152 20644
rect 21796 20700 21860 20704
rect 21796 20644 21800 20700
rect 21800 20644 21856 20700
rect 21856 20644 21860 20700
rect 21796 20640 21860 20644
rect 21876 20700 21940 20704
rect 21876 20644 21880 20700
rect 21880 20644 21936 20700
rect 21936 20644 21940 20700
rect 21876 20640 21940 20644
rect 21956 20700 22020 20704
rect 21956 20644 21960 20700
rect 21960 20644 22016 20700
rect 22016 20644 22020 20700
rect 21956 20640 22020 20644
rect 22036 20700 22100 20704
rect 22036 20644 22040 20700
rect 22040 20644 22096 20700
rect 22096 20644 22100 20700
rect 22036 20640 22100 20644
rect 4426 20156 4490 20160
rect 4426 20100 4430 20156
rect 4430 20100 4486 20156
rect 4486 20100 4490 20156
rect 4426 20096 4490 20100
rect 4506 20156 4570 20160
rect 4506 20100 4510 20156
rect 4510 20100 4566 20156
rect 4566 20100 4570 20156
rect 4506 20096 4570 20100
rect 4586 20156 4650 20160
rect 4586 20100 4590 20156
rect 4590 20100 4646 20156
rect 4646 20100 4650 20156
rect 4586 20096 4650 20100
rect 4666 20156 4730 20160
rect 4666 20100 4670 20156
rect 4670 20100 4726 20156
rect 4726 20100 4730 20156
rect 4666 20096 4730 20100
rect 11374 20156 11438 20160
rect 11374 20100 11378 20156
rect 11378 20100 11434 20156
rect 11434 20100 11438 20156
rect 11374 20096 11438 20100
rect 11454 20156 11518 20160
rect 11454 20100 11458 20156
rect 11458 20100 11514 20156
rect 11514 20100 11518 20156
rect 11454 20096 11518 20100
rect 11534 20156 11598 20160
rect 11534 20100 11538 20156
rect 11538 20100 11594 20156
rect 11594 20100 11598 20156
rect 11534 20096 11598 20100
rect 11614 20156 11678 20160
rect 11614 20100 11618 20156
rect 11618 20100 11674 20156
rect 11674 20100 11678 20156
rect 11614 20096 11678 20100
rect 18322 20156 18386 20160
rect 18322 20100 18326 20156
rect 18326 20100 18382 20156
rect 18382 20100 18386 20156
rect 18322 20096 18386 20100
rect 18402 20156 18466 20160
rect 18402 20100 18406 20156
rect 18406 20100 18462 20156
rect 18462 20100 18466 20156
rect 18402 20096 18466 20100
rect 18482 20156 18546 20160
rect 18482 20100 18486 20156
rect 18486 20100 18542 20156
rect 18542 20100 18546 20156
rect 18482 20096 18546 20100
rect 18562 20156 18626 20160
rect 18562 20100 18566 20156
rect 18566 20100 18622 20156
rect 18622 20100 18626 20156
rect 18562 20096 18626 20100
rect 25270 20156 25334 20160
rect 25270 20100 25274 20156
rect 25274 20100 25330 20156
rect 25330 20100 25334 20156
rect 25270 20096 25334 20100
rect 25350 20156 25414 20160
rect 25350 20100 25354 20156
rect 25354 20100 25410 20156
rect 25410 20100 25414 20156
rect 25350 20096 25414 20100
rect 25430 20156 25494 20160
rect 25430 20100 25434 20156
rect 25434 20100 25490 20156
rect 25490 20100 25494 20156
rect 25430 20096 25494 20100
rect 25510 20156 25574 20160
rect 25510 20100 25514 20156
rect 25514 20100 25570 20156
rect 25570 20100 25574 20156
rect 25510 20096 25574 20100
rect 7900 19612 7964 19616
rect 7900 19556 7904 19612
rect 7904 19556 7960 19612
rect 7960 19556 7964 19612
rect 7900 19552 7964 19556
rect 7980 19612 8044 19616
rect 7980 19556 7984 19612
rect 7984 19556 8040 19612
rect 8040 19556 8044 19612
rect 7980 19552 8044 19556
rect 8060 19612 8124 19616
rect 8060 19556 8064 19612
rect 8064 19556 8120 19612
rect 8120 19556 8124 19612
rect 8060 19552 8124 19556
rect 8140 19612 8204 19616
rect 8140 19556 8144 19612
rect 8144 19556 8200 19612
rect 8200 19556 8204 19612
rect 8140 19552 8204 19556
rect 14848 19612 14912 19616
rect 14848 19556 14852 19612
rect 14852 19556 14908 19612
rect 14908 19556 14912 19612
rect 14848 19552 14912 19556
rect 14928 19612 14992 19616
rect 14928 19556 14932 19612
rect 14932 19556 14988 19612
rect 14988 19556 14992 19612
rect 14928 19552 14992 19556
rect 15008 19612 15072 19616
rect 15008 19556 15012 19612
rect 15012 19556 15068 19612
rect 15068 19556 15072 19612
rect 15008 19552 15072 19556
rect 15088 19612 15152 19616
rect 15088 19556 15092 19612
rect 15092 19556 15148 19612
rect 15148 19556 15152 19612
rect 15088 19552 15152 19556
rect 21796 19612 21860 19616
rect 21796 19556 21800 19612
rect 21800 19556 21856 19612
rect 21856 19556 21860 19612
rect 21796 19552 21860 19556
rect 21876 19612 21940 19616
rect 21876 19556 21880 19612
rect 21880 19556 21936 19612
rect 21936 19556 21940 19612
rect 21876 19552 21940 19556
rect 21956 19612 22020 19616
rect 21956 19556 21960 19612
rect 21960 19556 22016 19612
rect 22016 19556 22020 19612
rect 21956 19552 22020 19556
rect 22036 19612 22100 19616
rect 22036 19556 22040 19612
rect 22040 19556 22096 19612
rect 22096 19556 22100 19612
rect 22036 19552 22100 19556
rect 4426 19068 4490 19072
rect 4426 19012 4430 19068
rect 4430 19012 4486 19068
rect 4486 19012 4490 19068
rect 4426 19008 4490 19012
rect 4506 19068 4570 19072
rect 4506 19012 4510 19068
rect 4510 19012 4566 19068
rect 4566 19012 4570 19068
rect 4506 19008 4570 19012
rect 4586 19068 4650 19072
rect 4586 19012 4590 19068
rect 4590 19012 4646 19068
rect 4646 19012 4650 19068
rect 4586 19008 4650 19012
rect 4666 19068 4730 19072
rect 4666 19012 4670 19068
rect 4670 19012 4726 19068
rect 4726 19012 4730 19068
rect 4666 19008 4730 19012
rect 11374 19068 11438 19072
rect 11374 19012 11378 19068
rect 11378 19012 11434 19068
rect 11434 19012 11438 19068
rect 11374 19008 11438 19012
rect 11454 19068 11518 19072
rect 11454 19012 11458 19068
rect 11458 19012 11514 19068
rect 11514 19012 11518 19068
rect 11454 19008 11518 19012
rect 11534 19068 11598 19072
rect 11534 19012 11538 19068
rect 11538 19012 11594 19068
rect 11594 19012 11598 19068
rect 11534 19008 11598 19012
rect 11614 19068 11678 19072
rect 11614 19012 11618 19068
rect 11618 19012 11674 19068
rect 11674 19012 11678 19068
rect 11614 19008 11678 19012
rect 18322 19068 18386 19072
rect 18322 19012 18326 19068
rect 18326 19012 18382 19068
rect 18382 19012 18386 19068
rect 18322 19008 18386 19012
rect 18402 19068 18466 19072
rect 18402 19012 18406 19068
rect 18406 19012 18462 19068
rect 18462 19012 18466 19068
rect 18402 19008 18466 19012
rect 18482 19068 18546 19072
rect 18482 19012 18486 19068
rect 18486 19012 18542 19068
rect 18542 19012 18546 19068
rect 18482 19008 18546 19012
rect 18562 19068 18626 19072
rect 18562 19012 18566 19068
rect 18566 19012 18622 19068
rect 18622 19012 18626 19068
rect 18562 19008 18626 19012
rect 25270 19068 25334 19072
rect 25270 19012 25274 19068
rect 25274 19012 25330 19068
rect 25330 19012 25334 19068
rect 25270 19008 25334 19012
rect 25350 19068 25414 19072
rect 25350 19012 25354 19068
rect 25354 19012 25410 19068
rect 25410 19012 25414 19068
rect 25350 19008 25414 19012
rect 25430 19068 25494 19072
rect 25430 19012 25434 19068
rect 25434 19012 25490 19068
rect 25490 19012 25494 19068
rect 25430 19008 25494 19012
rect 25510 19068 25574 19072
rect 25510 19012 25514 19068
rect 25514 19012 25570 19068
rect 25570 19012 25574 19068
rect 25510 19008 25574 19012
rect 7900 18524 7964 18528
rect 7900 18468 7904 18524
rect 7904 18468 7960 18524
rect 7960 18468 7964 18524
rect 7900 18464 7964 18468
rect 7980 18524 8044 18528
rect 7980 18468 7984 18524
rect 7984 18468 8040 18524
rect 8040 18468 8044 18524
rect 7980 18464 8044 18468
rect 8060 18524 8124 18528
rect 8060 18468 8064 18524
rect 8064 18468 8120 18524
rect 8120 18468 8124 18524
rect 8060 18464 8124 18468
rect 8140 18524 8204 18528
rect 8140 18468 8144 18524
rect 8144 18468 8200 18524
rect 8200 18468 8204 18524
rect 8140 18464 8204 18468
rect 14848 18524 14912 18528
rect 14848 18468 14852 18524
rect 14852 18468 14908 18524
rect 14908 18468 14912 18524
rect 14848 18464 14912 18468
rect 14928 18524 14992 18528
rect 14928 18468 14932 18524
rect 14932 18468 14988 18524
rect 14988 18468 14992 18524
rect 14928 18464 14992 18468
rect 15008 18524 15072 18528
rect 15008 18468 15012 18524
rect 15012 18468 15068 18524
rect 15068 18468 15072 18524
rect 15008 18464 15072 18468
rect 15088 18524 15152 18528
rect 15088 18468 15092 18524
rect 15092 18468 15148 18524
rect 15148 18468 15152 18524
rect 15088 18464 15152 18468
rect 21796 18524 21860 18528
rect 21796 18468 21800 18524
rect 21800 18468 21856 18524
rect 21856 18468 21860 18524
rect 21796 18464 21860 18468
rect 21876 18524 21940 18528
rect 21876 18468 21880 18524
rect 21880 18468 21936 18524
rect 21936 18468 21940 18524
rect 21876 18464 21940 18468
rect 21956 18524 22020 18528
rect 21956 18468 21960 18524
rect 21960 18468 22016 18524
rect 22016 18468 22020 18524
rect 21956 18464 22020 18468
rect 22036 18524 22100 18528
rect 22036 18468 22040 18524
rect 22040 18468 22096 18524
rect 22096 18468 22100 18524
rect 22036 18464 22100 18468
rect 4426 17980 4490 17984
rect 4426 17924 4430 17980
rect 4430 17924 4486 17980
rect 4486 17924 4490 17980
rect 4426 17920 4490 17924
rect 4506 17980 4570 17984
rect 4506 17924 4510 17980
rect 4510 17924 4566 17980
rect 4566 17924 4570 17980
rect 4506 17920 4570 17924
rect 4586 17980 4650 17984
rect 4586 17924 4590 17980
rect 4590 17924 4646 17980
rect 4646 17924 4650 17980
rect 4586 17920 4650 17924
rect 4666 17980 4730 17984
rect 4666 17924 4670 17980
rect 4670 17924 4726 17980
rect 4726 17924 4730 17980
rect 4666 17920 4730 17924
rect 11374 17980 11438 17984
rect 11374 17924 11378 17980
rect 11378 17924 11434 17980
rect 11434 17924 11438 17980
rect 11374 17920 11438 17924
rect 11454 17980 11518 17984
rect 11454 17924 11458 17980
rect 11458 17924 11514 17980
rect 11514 17924 11518 17980
rect 11454 17920 11518 17924
rect 11534 17980 11598 17984
rect 11534 17924 11538 17980
rect 11538 17924 11594 17980
rect 11594 17924 11598 17980
rect 11534 17920 11598 17924
rect 11614 17980 11678 17984
rect 11614 17924 11618 17980
rect 11618 17924 11674 17980
rect 11674 17924 11678 17980
rect 11614 17920 11678 17924
rect 18322 17980 18386 17984
rect 18322 17924 18326 17980
rect 18326 17924 18382 17980
rect 18382 17924 18386 17980
rect 18322 17920 18386 17924
rect 18402 17980 18466 17984
rect 18402 17924 18406 17980
rect 18406 17924 18462 17980
rect 18462 17924 18466 17980
rect 18402 17920 18466 17924
rect 18482 17980 18546 17984
rect 18482 17924 18486 17980
rect 18486 17924 18542 17980
rect 18542 17924 18546 17980
rect 18482 17920 18546 17924
rect 18562 17980 18626 17984
rect 18562 17924 18566 17980
rect 18566 17924 18622 17980
rect 18622 17924 18626 17980
rect 18562 17920 18626 17924
rect 25270 17980 25334 17984
rect 25270 17924 25274 17980
rect 25274 17924 25330 17980
rect 25330 17924 25334 17980
rect 25270 17920 25334 17924
rect 25350 17980 25414 17984
rect 25350 17924 25354 17980
rect 25354 17924 25410 17980
rect 25410 17924 25414 17980
rect 25350 17920 25414 17924
rect 25430 17980 25494 17984
rect 25430 17924 25434 17980
rect 25434 17924 25490 17980
rect 25490 17924 25494 17980
rect 25430 17920 25494 17924
rect 25510 17980 25574 17984
rect 25510 17924 25514 17980
rect 25514 17924 25570 17980
rect 25570 17924 25574 17980
rect 25510 17920 25574 17924
rect 7900 17436 7964 17440
rect 7900 17380 7904 17436
rect 7904 17380 7960 17436
rect 7960 17380 7964 17436
rect 7900 17376 7964 17380
rect 7980 17436 8044 17440
rect 7980 17380 7984 17436
rect 7984 17380 8040 17436
rect 8040 17380 8044 17436
rect 7980 17376 8044 17380
rect 8060 17436 8124 17440
rect 8060 17380 8064 17436
rect 8064 17380 8120 17436
rect 8120 17380 8124 17436
rect 8060 17376 8124 17380
rect 8140 17436 8204 17440
rect 8140 17380 8144 17436
rect 8144 17380 8200 17436
rect 8200 17380 8204 17436
rect 8140 17376 8204 17380
rect 14848 17436 14912 17440
rect 14848 17380 14852 17436
rect 14852 17380 14908 17436
rect 14908 17380 14912 17436
rect 14848 17376 14912 17380
rect 14928 17436 14992 17440
rect 14928 17380 14932 17436
rect 14932 17380 14988 17436
rect 14988 17380 14992 17436
rect 14928 17376 14992 17380
rect 15008 17436 15072 17440
rect 15008 17380 15012 17436
rect 15012 17380 15068 17436
rect 15068 17380 15072 17436
rect 15008 17376 15072 17380
rect 15088 17436 15152 17440
rect 15088 17380 15092 17436
rect 15092 17380 15148 17436
rect 15148 17380 15152 17436
rect 15088 17376 15152 17380
rect 21796 17436 21860 17440
rect 21796 17380 21800 17436
rect 21800 17380 21856 17436
rect 21856 17380 21860 17436
rect 21796 17376 21860 17380
rect 21876 17436 21940 17440
rect 21876 17380 21880 17436
rect 21880 17380 21936 17436
rect 21936 17380 21940 17436
rect 21876 17376 21940 17380
rect 21956 17436 22020 17440
rect 21956 17380 21960 17436
rect 21960 17380 22016 17436
rect 22016 17380 22020 17436
rect 21956 17376 22020 17380
rect 22036 17436 22100 17440
rect 22036 17380 22040 17436
rect 22040 17380 22096 17436
rect 22096 17380 22100 17436
rect 22036 17376 22100 17380
rect 4426 16892 4490 16896
rect 4426 16836 4430 16892
rect 4430 16836 4486 16892
rect 4486 16836 4490 16892
rect 4426 16832 4490 16836
rect 4506 16892 4570 16896
rect 4506 16836 4510 16892
rect 4510 16836 4566 16892
rect 4566 16836 4570 16892
rect 4506 16832 4570 16836
rect 4586 16892 4650 16896
rect 4586 16836 4590 16892
rect 4590 16836 4646 16892
rect 4646 16836 4650 16892
rect 4586 16832 4650 16836
rect 4666 16892 4730 16896
rect 4666 16836 4670 16892
rect 4670 16836 4726 16892
rect 4726 16836 4730 16892
rect 4666 16832 4730 16836
rect 11374 16892 11438 16896
rect 11374 16836 11378 16892
rect 11378 16836 11434 16892
rect 11434 16836 11438 16892
rect 11374 16832 11438 16836
rect 11454 16892 11518 16896
rect 11454 16836 11458 16892
rect 11458 16836 11514 16892
rect 11514 16836 11518 16892
rect 11454 16832 11518 16836
rect 11534 16892 11598 16896
rect 11534 16836 11538 16892
rect 11538 16836 11594 16892
rect 11594 16836 11598 16892
rect 11534 16832 11598 16836
rect 11614 16892 11678 16896
rect 11614 16836 11618 16892
rect 11618 16836 11674 16892
rect 11674 16836 11678 16892
rect 11614 16832 11678 16836
rect 18322 16892 18386 16896
rect 18322 16836 18326 16892
rect 18326 16836 18382 16892
rect 18382 16836 18386 16892
rect 18322 16832 18386 16836
rect 18402 16892 18466 16896
rect 18402 16836 18406 16892
rect 18406 16836 18462 16892
rect 18462 16836 18466 16892
rect 18402 16832 18466 16836
rect 18482 16892 18546 16896
rect 18482 16836 18486 16892
rect 18486 16836 18542 16892
rect 18542 16836 18546 16892
rect 18482 16832 18546 16836
rect 18562 16892 18626 16896
rect 18562 16836 18566 16892
rect 18566 16836 18622 16892
rect 18622 16836 18626 16892
rect 18562 16832 18626 16836
rect 25270 16892 25334 16896
rect 25270 16836 25274 16892
rect 25274 16836 25330 16892
rect 25330 16836 25334 16892
rect 25270 16832 25334 16836
rect 25350 16892 25414 16896
rect 25350 16836 25354 16892
rect 25354 16836 25410 16892
rect 25410 16836 25414 16892
rect 25350 16832 25414 16836
rect 25430 16892 25494 16896
rect 25430 16836 25434 16892
rect 25434 16836 25490 16892
rect 25490 16836 25494 16892
rect 25430 16832 25494 16836
rect 25510 16892 25574 16896
rect 25510 16836 25514 16892
rect 25514 16836 25570 16892
rect 25570 16836 25574 16892
rect 25510 16832 25574 16836
rect 7900 16348 7964 16352
rect 7900 16292 7904 16348
rect 7904 16292 7960 16348
rect 7960 16292 7964 16348
rect 7900 16288 7964 16292
rect 7980 16348 8044 16352
rect 7980 16292 7984 16348
rect 7984 16292 8040 16348
rect 8040 16292 8044 16348
rect 7980 16288 8044 16292
rect 8060 16348 8124 16352
rect 8060 16292 8064 16348
rect 8064 16292 8120 16348
rect 8120 16292 8124 16348
rect 8060 16288 8124 16292
rect 8140 16348 8204 16352
rect 8140 16292 8144 16348
rect 8144 16292 8200 16348
rect 8200 16292 8204 16348
rect 8140 16288 8204 16292
rect 14848 16348 14912 16352
rect 14848 16292 14852 16348
rect 14852 16292 14908 16348
rect 14908 16292 14912 16348
rect 14848 16288 14912 16292
rect 14928 16348 14992 16352
rect 14928 16292 14932 16348
rect 14932 16292 14988 16348
rect 14988 16292 14992 16348
rect 14928 16288 14992 16292
rect 15008 16348 15072 16352
rect 15008 16292 15012 16348
rect 15012 16292 15068 16348
rect 15068 16292 15072 16348
rect 15008 16288 15072 16292
rect 15088 16348 15152 16352
rect 15088 16292 15092 16348
rect 15092 16292 15148 16348
rect 15148 16292 15152 16348
rect 15088 16288 15152 16292
rect 21796 16348 21860 16352
rect 21796 16292 21800 16348
rect 21800 16292 21856 16348
rect 21856 16292 21860 16348
rect 21796 16288 21860 16292
rect 21876 16348 21940 16352
rect 21876 16292 21880 16348
rect 21880 16292 21936 16348
rect 21936 16292 21940 16348
rect 21876 16288 21940 16292
rect 21956 16348 22020 16352
rect 21956 16292 21960 16348
rect 21960 16292 22016 16348
rect 22016 16292 22020 16348
rect 21956 16288 22020 16292
rect 22036 16348 22100 16352
rect 22036 16292 22040 16348
rect 22040 16292 22096 16348
rect 22096 16292 22100 16348
rect 22036 16288 22100 16292
rect 4426 15804 4490 15808
rect 4426 15748 4430 15804
rect 4430 15748 4486 15804
rect 4486 15748 4490 15804
rect 4426 15744 4490 15748
rect 4506 15804 4570 15808
rect 4506 15748 4510 15804
rect 4510 15748 4566 15804
rect 4566 15748 4570 15804
rect 4506 15744 4570 15748
rect 4586 15804 4650 15808
rect 4586 15748 4590 15804
rect 4590 15748 4646 15804
rect 4646 15748 4650 15804
rect 4586 15744 4650 15748
rect 4666 15804 4730 15808
rect 4666 15748 4670 15804
rect 4670 15748 4726 15804
rect 4726 15748 4730 15804
rect 4666 15744 4730 15748
rect 11374 15804 11438 15808
rect 11374 15748 11378 15804
rect 11378 15748 11434 15804
rect 11434 15748 11438 15804
rect 11374 15744 11438 15748
rect 11454 15804 11518 15808
rect 11454 15748 11458 15804
rect 11458 15748 11514 15804
rect 11514 15748 11518 15804
rect 11454 15744 11518 15748
rect 11534 15804 11598 15808
rect 11534 15748 11538 15804
rect 11538 15748 11594 15804
rect 11594 15748 11598 15804
rect 11534 15744 11598 15748
rect 11614 15804 11678 15808
rect 11614 15748 11618 15804
rect 11618 15748 11674 15804
rect 11674 15748 11678 15804
rect 11614 15744 11678 15748
rect 18322 15804 18386 15808
rect 18322 15748 18326 15804
rect 18326 15748 18382 15804
rect 18382 15748 18386 15804
rect 18322 15744 18386 15748
rect 18402 15804 18466 15808
rect 18402 15748 18406 15804
rect 18406 15748 18462 15804
rect 18462 15748 18466 15804
rect 18402 15744 18466 15748
rect 18482 15804 18546 15808
rect 18482 15748 18486 15804
rect 18486 15748 18542 15804
rect 18542 15748 18546 15804
rect 18482 15744 18546 15748
rect 18562 15804 18626 15808
rect 18562 15748 18566 15804
rect 18566 15748 18622 15804
rect 18622 15748 18626 15804
rect 18562 15744 18626 15748
rect 25270 15804 25334 15808
rect 25270 15748 25274 15804
rect 25274 15748 25330 15804
rect 25330 15748 25334 15804
rect 25270 15744 25334 15748
rect 25350 15804 25414 15808
rect 25350 15748 25354 15804
rect 25354 15748 25410 15804
rect 25410 15748 25414 15804
rect 25350 15744 25414 15748
rect 25430 15804 25494 15808
rect 25430 15748 25434 15804
rect 25434 15748 25490 15804
rect 25490 15748 25494 15804
rect 25430 15744 25494 15748
rect 25510 15804 25574 15808
rect 25510 15748 25514 15804
rect 25514 15748 25570 15804
rect 25570 15748 25574 15804
rect 25510 15744 25574 15748
rect 7900 15260 7964 15264
rect 7900 15204 7904 15260
rect 7904 15204 7960 15260
rect 7960 15204 7964 15260
rect 7900 15200 7964 15204
rect 7980 15260 8044 15264
rect 7980 15204 7984 15260
rect 7984 15204 8040 15260
rect 8040 15204 8044 15260
rect 7980 15200 8044 15204
rect 8060 15260 8124 15264
rect 8060 15204 8064 15260
rect 8064 15204 8120 15260
rect 8120 15204 8124 15260
rect 8060 15200 8124 15204
rect 8140 15260 8204 15264
rect 8140 15204 8144 15260
rect 8144 15204 8200 15260
rect 8200 15204 8204 15260
rect 8140 15200 8204 15204
rect 14848 15260 14912 15264
rect 14848 15204 14852 15260
rect 14852 15204 14908 15260
rect 14908 15204 14912 15260
rect 14848 15200 14912 15204
rect 14928 15260 14992 15264
rect 14928 15204 14932 15260
rect 14932 15204 14988 15260
rect 14988 15204 14992 15260
rect 14928 15200 14992 15204
rect 15008 15260 15072 15264
rect 15008 15204 15012 15260
rect 15012 15204 15068 15260
rect 15068 15204 15072 15260
rect 15008 15200 15072 15204
rect 15088 15260 15152 15264
rect 15088 15204 15092 15260
rect 15092 15204 15148 15260
rect 15148 15204 15152 15260
rect 15088 15200 15152 15204
rect 21796 15260 21860 15264
rect 21796 15204 21800 15260
rect 21800 15204 21856 15260
rect 21856 15204 21860 15260
rect 21796 15200 21860 15204
rect 21876 15260 21940 15264
rect 21876 15204 21880 15260
rect 21880 15204 21936 15260
rect 21936 15204 21940 15260
rect 21876 15200 21940 15204
rect 21956 15260 22020 15264
rect 21956 15204 21960 15260
rect 21960 15204 22016 15260
rect 22016 15204 22020 15260
rect 21956 15200 22020 15204
rect 22036 15260 22100 15264
rect 22036 15204 22040 15260
rect 22040 15204 22096 15260
rect 22096 15204 22100 15260
rect 22036 15200 22100 15204
rect 4426 14716 4490 14720
rect 4426 14660 4430 14716
rect 4430 14660 4486 14716
rect 4486 14660 4490 14716
rect 4426 14656 4490 14660
rect 4506 14716 4570 14720
rect 4506 14660 4510 14716
rect 4510 14660 4566 14716
rect 4566 14660 4570 14716
rect 4506 14656 4570 14660
rect 4586 14716 4650 14720
rect 4586 14660 4590 14716
rect 4590 14660 4646 14716
rect 4646 14660 4650 14716
rect 4586 14656 4650 14660
rect 4666 14716 4730 14720
rect 4666 14660 4670 14716
rect 4670 14660 4726 14716
rect 4726 14660 4730 14716
rect 4666 14656 4730 14660
rect 11374 14716 11438 14720
rect 11374 14660 11378 14716
rect 11378 14660 11434 14716
rect 11434 14660 11438 14716
rect 11374 14656 11438 14660
rect 11454 14716 11518 14720
rect 11454 14660 11458 14716
rect 11458 14660 11514 14716
rect 11514 14660 11518 14716
rect 11454 14656 11518 14660
rect 11534 14716 11598 14720
rect 11534 14660 11538 14716
rect 11538 14660 11594 14716
rect 11594 14660 11598 14716
rect 11534 14656 11598 14660
rect 11614 14716 11678 14720
rect 11614 14660 11618 14716
rect 11618 14660 11674 14716
rect 11674 14660 11678 14716
rect 11614 14656 11678 14660
rect 18322 14716 18386 14720
rect 18322 14660 18326 14716
rect 18326 14660 18382 14716
rect 18382 14660 18386 14716
rect 18322 14656 18386 14660
rect 18402 14716 18466 14720
rect 18402 14660 18406 14716
rect 18406 14660 18462 14716
rect 18462 14660 18466 14716
rect 18402 14656 18466 14660
rect 18482 14716 18546 14720
rect 18482 14660 18486 14716
rect 18486 14660 18542 14716
rect 18542 14660 18546 14716
rect 18482 14656 18546 14660
rect 18562 14716 18626 14720
rect 18562 14660 18566 14716
rect 18566 14660 18622 14716
rect 18622 14660 18626 14716
rect 18562 14656 18626 14660
rect 25270 14716 25334 14720
rect 25270 14660 25274 14716
rect 25274 14660 25330 14716
rect 25330 14660 25334 14716
rect 25270 14656 25334 14660
rect 25350 14716 25414 14720
rect 25350 14660 25354 14716
rect 25354 14660 25410 14716
rect 25410 14660 25414 14716
rect 25350 14656 25414 14660
rect 25430 14716 25494 14720
rect 25430 14660 25434 14716
rect 25434 14660 25490 14716
rect 25490 14660 25494 14716
rect 25430 14656 25494 14660
rect 25510 14716 25574 14720
rect 25510 14660 25514 14716
rect 25514 14660 25570 14716
rect 25570 14660 25574 14716
rect 25510 14656 25574 14660
rect 7900 14172 7964 14176
rect 7900 14116 7904 14172
rect 7904 14116 7960 14172
rect 7960 14116 7964 14172
rect 7900 14112 7964 14116
rect 7980 14172 8044 14176
rect 7980 14116 7984 14172
rect 7984 14116 8040 14172
rect 8040 14116 8044 14172
rect 7980 14112 8044 14116
rect 8060 14172 8124 14176
rect 8060 14116 8064 14172
rect 8064 14116 8120 14172
rect 8120 14116 8124 14172
rect 8060 14112 8124 14116
rect 8140 14172 8204 14176
rect 8140 14116 8144 14172
rect 8144 14116 8200 14172
rect 8200 14116 8204 14172
rect 8140 14112 8204 14116
rect 14848 14172 14912 14176
rect 14848 14116 14852 14172
rect 14852 14116 14908 14172
rect 14908 14116 14912 14172
rect 14848 14112 14912 14116
rect 14928 14172 14992 14176
rect 14928 14116 14932 14172
rect 14932 14116 14988 14172
rect 14988 14116 14992 14172
rect 14928 14112 14992 14116
rect 15008 14172 15072 14176
rect 15008 14116 15012 14172
rect 15012 14116 15068 14172
rect 15068 14116 15072 14172
rect 15008 14112 15072 14116
rect 15088 14172 15152 14176
rect 15088 14116 15092 14172
rect 15092 14116 15148 14172
rect 15148 14116 15152 14172
rect 15088 14112 15152 14116
rect 21796 14172 21860 14176
rect 21796 14116 21800 14172
rect 21800 14116 21856 14172
rect 21856 14116 21860 14172
rect 21796 14112 21860 14116
rect 21876 14172 21940 14176
rect 21876 14116 21880 14172
rect 21880 14116 21936 14172
rect 21936 14116 21940 14172
rect 21876 14112 21940 14116
rect 21956 14172 22020 14176
rect 21956 14116 21960 14172
rect 21960 14116 22016 14172
rect 22016 14116 22020 14172
rect 21956 14112 22020 14116
rect 22036 14172 22100 14176
rect 22036 14116 22040 14172
rect 22040 14116 22096 14172
rect 22096 14116 22100 14172
rect 22036 14112 22100 14116
rect 4426 13628 4490 13632
rect 4426 13572 4430 13628
rect 4430 13572 4486 13628
rect 4486 13572 4490 13628
rect 4426 13568 4490 13572
rect 4506 13628 4570 13632
rect 4506 13572 4510 13628
rect 4510 13572 4566 13628
rect 4566 13572 4570 13628
rect 4506 13568 4570 13572
rect 4586 13628 4650 13632
rect 4586 13572 4590 13628
rect 4590 13572 4646 13628
rect 4646 13572 4650 13628
rect 4586 13568 4650 13572
rect 4666 13628 4730 13632
rect 4666 13572 4670 13628
rect 4670 13572 4726 13628
rect 4726 13572 4730 13628
rect 4666 13568 4730 13572
rect 11374 13628 11438 13632
rect 11374 13572 11378 13628
rect 11378 13572 11434 13628
rect 11434 13572 11438 13628
rect 11374 13568 11438 13572
rect 11454 13628 11518 13632
rect 11454 13572 11458 13628
rect 11458 13572 11514 13628
rect 11514 13572 11518 13628
rect 11454 13568 11518 13572
rect 11534 13628 11598 13632
rect 11534 13572 11538 13628
rect 11538 13572 11594 13628
rect 11594 13572 11598 13628
rect 11534 13568 11598 13572
rect 11614 13628 11678 13632
rect 11614 13572 11618 13628
rect 11618 13572 11674 13628
rect 11674 13572 11678 13628
rect 11614 13568 11678 13572
rect 18322 13628 18386 13632
rect 18322 13572 18326 13628
rect 18326 13572 18382 13628
rect 18382 13572 18386 13628
rect 18322 13568 18386 13572
rect 18402 13628 18466 13632
rect 18402 13572 18406 13628
rect 18406 13572 18462 13628
rect 18462 13572 18466 13628
rect 18402 13568 18466 13572
rect 18482 13628 18546 13632
rect 18482 13572 18486 13628
rect 18486 13572 18542 13628
rect 18542 13572 18546 13628
rect 18482 13568 18546 13572
rect 18562 13628 18626 13632
rect 18562 13572 18566 13628
rect 18566 13572 18622 13628
rect 18622 13572 18626 13628
rect 18562 13568 18626 13572
rect 25270 13628 25334 13632
rect 25270 13572 25274 13628
rect 25274 13572 25330 13628
rect 25330 13572 25334 13628
rect 25270 13568 25334 13572
rect 25350 13628 25414 13632
rect 25350 13572 25354 13628
rect 25354 13572 25410 13628
rect 25410 13572 25414 13628
rect 25350 13568 25414 13572
rect 25430 13628 25494 13632
rect 25430 13572 25434 13628
rect 25434 13572 25490 13628
rect 25490 13572 25494 13628
rect 25430 13568 25494 13572
rect 25510 13628 25574 13632
rect 25510 13572 25514 13628
rect 25514 13572 25570 13628
rect 25570 13572 25574 13628
rect 25510 13568 25574 13572
rect 7900 13084 7964 13088
rect 7900 13028 7904 13084
rect 7904 13028 7960 13084
rect 7960 13028 7964 13084
rect 7900 13024 7964 13028
rect 7980 13084 8044 13088
rect 7980 13028 7984 13084
rect 7984 13028 8040 13084
rect 8040 13028 8044 13084
rect 7980 13024 8044 13028
rect 8060 13084 8124 13088
rect 8060 13028 8064 13084
rect 8064 13028 8120 13084
rect 8120 13028 8124 13084
rect 8060 13024 8124 13028
rect 8140 13084 8204 13088
rect 8140 13028 8144 13084
rect 8144 13028 8200 13084
rect 8200 13028 8204 13084
rect 8140 13024 8204 13028
rect 14848 13084 14912 13088
rect 14848 13028 14852 13084
rect 14852 13028 14908 13084
rect 14908 13028 14912 13084
rect 14848 13024 14912 13028
rect 14928 13084 14992 13088
rect 14928 13028 14932 13084
rect 14932 13028 14988 13084
rect 14988 13028 14992 13084
rect 14928 13024 14992 13028
rect 15008 13084 15072 13088
rect 15008 13028 15012 13084
rect 15012 13028 15068 13084
rect 15068 13028 15072 13084
rect 15008 13024 15072 13028
rect 15088 13084 15152 13088
rect 15088 13028 15092 13084
rect 15092 13028 15148 13084
rect 15148 13028 15152 13084
rect 15088 13024 15152 13028
rect 21796 13084 21860 13088
rect 21796 13028 21800 13084
rect 21800 13028 21856 13084
rect 21856 13028 21860 13084
rect 21796 13024 21860 13028
rect 21876 13084 21940 13088
rect 21876 13028 21880 13084
rect 21880 13028 21936 13084
rect 21936 13028 21940 13084
rect 21876 13024 21940 13028
rect 21956 13084 22020 13088
rect 21956 13028 21960 13084
rect 21960 13028 22016 13084
rect 22016 13028 22020 13084
rect 21956 13024 22020 13028
rect 22036 13084 22100 13088
rect 22036 13028 22040 13084
rect 22040 13028 22096 13084
rect 22096 13028 22100 13084
rect 22036 13024 22100 13028
rect 4426 12540 4490 12544
rect 4426 12484 4430 12540
rect 4430 12484 4486 12540
rect 4486 12484 4490 12540
rect 4426 12480 4490 12484
rect 4506 12540 4570 12544
rect 4506 12484 4510 12540
rect 4510 12484 4566 12540
rect 4566 12484 4570 12540
rect 4506 12480 4570 12484
rect 4586 12540 4650 12544
rect 4586 12484 4590 12540
rect 4590 12484 4646 12540
rect 4646 12484 4650 12540
rect 4586 12480 4650 12484
rect 4666 12540 4730 12544
rect 4666 12484 4670 12540
rect 4670 12484 4726 12540
rect 4726 12484 4730 12540
rect 4666 12480 4730 12484
rect 11374 12540 11438 12544
rect 11374 12484 11378 12540
rect 11378 12484 11434 12540
rect 11434 12484 11438 12540
rect 11374 12480 11438 12484
rect 11454 12540 11518 12544
rect 11454 12484 11458 12540
rect 11458 12484 11514 12540
rect 11514 12484 11518 12540
rect 11454 12480 11518 12484
rect 11534 12540 11598 12544
rect 11534 12484 11538 12540
rect 11538 12484 11594 12540
rect 11594 12484 11598 12540
rect 11534 12480 11598 12484
rect 11614 12540 11678 12544
rect 11614 12484 11618 12540
rect 11618 12484 11674 12540
rect 11674 12484 11678 12540
rect 11614 12480 11678 12484
rect 18322 12540 18386 12544
rect 18322 12484 18326 12540
rect 18326 12484 18382 12540
rect 18382 12484 18386 12540
rect 18322 12480 18386 12484
rect 18402 12540 18466 12544
rect 18402 12484 18406 12540
rect 18406 12484 18462 12540
rect 18462 12484 18466 12540
rect 18402 12480 18466 12484
rect 18482 12540 18546 12544
rect 18482 12484 18486 12540
rect 18486 12484 18542 12540
rect 18542 12484 18546 12540
rect 18482 12480 18546 12484
rect 18562 12540 18626 12544
rect 18562 12484 18566 12540
rect 18566 12484 18622 12540
rect 18622 12484 18626 12540
rect 18562 12480 18626 12484
rect 25270 12540 25334 12544
rect 25270 12484 25274 12540
rect 25274 12484 25330 12540
rect 25330 12484 25334 12540
rect 25270 12480 25334 12484
rect 25350 12540 25414 12544
rect 25350 12484 25354 12540
rect 25354 12484 25410 12540
rect 25410 12484 25414 12540
rect 25350 12480 25414 12484
rect 25430 12540 25494 12544
rect 25430 12484 25434 12540
rect 25434 12484 25490 12540
rect 25490 12484 25494 12540
rect 25430 12480 25494 12484
rect 25510 12540 25574 12544
rect 25510 12484 25514 12540
rect 25514 12484 25570 12540
rect 25570 12484 25574 12540
rect 25510 12480 25574 12484
rect 7900 11996 7964 12000
rect 7900 11940 7904 11996
rect 7904 11940 7960 11996
rect 7960 11940 7964 11996
rect 7900 11936 7964 11940
rect 7980 11996 8044 12000
rect 7980 11940 7984 11996
rect 7984 11940 8040 11996
rect 8040 11940 8044 11996
rect 7980 11936 8044 11940
rect 8060 11996 8124 12000
rect 8060 11940 8064 11996
rect 8064 11940 8120 11996
rect 8120 11940 8124 11996
rect 8060 11936 8124 11940
rect 8140 11996 8204 12000
rect 8140 11940 8144 11996
rect 8144 11940 8200 11996
rect 8200 11940 8204 11996
rect 8140 11936 8204 11940
rect 14848 11996 14912 12000
rect 14848 11940 14852 11996
rect 14852 11940 14908 11996
rect 14908 11940 14912 11996
rect 14848 11936 14912 11940
rect 14928 11996 14992 12000
rect 14928 11940 14932 11996
rect 14932 11940 14988 11996
rect 14988 11940 14992 11996
rect 14928 11936 14992 11940
rect 15008 11996 15072 12000
rect 15008 11940 15012 11996
rect 15012 11940 15068 11996
rect 15068 11940 15072 11996
rect 15008 11936 15072 11940
rect 15088 11996 15152 12000
rect 15088 11940 15092 11996
rect 15092 11940 15148 11996
rect 15148 11940 15152 11996
rect 15088 11936 15152 11940
rect 21796 11996 21860 12000
rect 21796 11940 21800 11996
rect 21800 11940 21856 11996
rect 21856 11940 21860 11996
rect 21796 11936 21860 11940
rect 21876 11996 21940 12000
rect 21876 11940 21880 11996
rect 21880 11940 21936 11996
rect 21936 11940 21940 11996
rect 21876 11936 21940 11940
rect 21956 11996 22020 12000
rect 21956 11940 21960 11996
rect 21960 11940 22016 11996
rect 22016 11940 22020 11996
rect 21956 11936 22020 11940
rect 22036 11996 22100 12000
rect 22036 11940 22040 11996
rect 22040 11940 22096 11996
rect 22096 11940 22100 11996
rect 22036 11936 22100 11940
rect 4426 11452 4490 11456
rect 4426 11396 4430 11452
rect 4430 11396 4486 11452
rect 4486 11396 4490 11452
rect 4426 11392 4490 11396
rect 4506 11452 4570 11456
rect 4506 11396 4510 11452
rect 4510 11396 4566 11452
rect 4566 11396 4570 11452
rect 4506 11392 4570 11396
rect 4586 11452 4650 11456
rect 4586 11396 4590 11452
rect 4590 11396 4646 11452
rect 4646 11396 4650 11452
rect 4586 11392 4650 11396
rect 4666 11452 4730 11456
rect 4666 11396 4670 11452
rect 4670 11396 4726 11452
rect 4726 11396 4730 11452
rect 4666 11392 4730 11396
rect 11374 11452 11438 11456
rect 11374 11396 11378 11452
rect 11378 11396 11434 11452
rect 11434 11396 11438 11452
rect 11374 11392 11438 11396
rect 11454 11452 11518 11456
rect 11454 11396 11458 11452
rect 11458 11396 11514 11452
rect 11514 11396 11518 11452
rect 11454 11392 11518 11396
rect 11534 11452 11598 11456
rect 11534 11396 11538 11452
rect 11538 11396 11594 11452
rect 11594 11396 11598 11452
rect 11534 11392 11598 11396
rect 11614 11452 11678 11456
rect 11614 11396 11618 11452
rect 11618 11396 11674 11452
rect 11674 11396 11678 11452
rect 11614 11392 11678 11396
rect 18322 11452 18386 11456
rect 18322 11396 18326 11452
rect 18326 11396 18382 11452
rect 18382 11396 18386 11452
rect 18322 11392 18386 11396
rect 18402 11452 18466 11456
rect 18402 11396 18406 11452
rect 18406 11396 18462 11452
rect 18462 11396 18466 11452
rect 18402 11392 18466 11396
rect 18482 11452 18546 11456
rect 18482 11396 18486 11452
rect 18486 11396 18542 11452
rect 18542 11396 18546 11452
rect 18482 11392 18546 11396
rect 18562 11452 18626 11456
rect 18562 11396 18566 11452
rect 18566 11396 18622 11452
rect 18622 11396 18626 11452
rect 18562 11392 18626 11396
rect 25270 11452 25334 11456
rect 25270 11396 25274 11452
rect 25274 11396 25330 11452
rect 25330 11396 25334 11452
rect 25270 11392 25334 11396
rect 25350 11452 25414 11456
rect 25350 11396 25354 11452
rect 25354 11396 25410 11452
rect 25410 11396 25414 11452
rect 25350 11392 25414 11396
rect 25430 11452 25494 11456
rect 25430 11396 25434 11452
rect 25434 11396 25490 11452
rect 25490 11396 25494 11452
rect 25430 11392 25494 11396
rect 25510 11452 25574 11456
rect 25510 11396 25514 11452
rect 25514 11396 25570 11452
rect 25570 11396 25574 11452
rect 25510 11392 25574 11396
rect 7900 10908 7964 10912
rect 7900 10852 7904 10908
rect 7904 10852 7960 10908
rect 7960 10852 7964 10908
rect 7900 10848 7964 10852
rect 7980 10908 8044 10912
rect 7980 10852 7984 10908
rect 7984 10852 8040 10908
rect 8040 10852 8044 10908
rect 7980 10848 8044 10852
rect 8060 10908 8124 10912
rect 8060 10852 8064 10908
rect 8064 10852 8120 10908
rect 8120 10852 8124 10908
rect 8060 10848 8124 10852
rect 8140 10908 8204 10912
rect 8140 10852 8144 10908
rect 8144 10852 8200 10908
rect 8200 10852 8204 10908
rect 8140 10848 8204 10852
rect 14848 10908 14912 10912
rect 14848 10852 14852 10908
rect 14852 10852 14908 10908
rect 14908 10852 14912 10908
rect 14848 10848 14912 10852
rect 14928 10908 14992 10912
rect 14928 10852 14932 10908
rect 14932 10852 14988 10908
rect 14988 10852 14992 10908
rect 14928 10848 14992 10852
rect 15008 10908 15072 10912
rect 15008 10852 15012 10908
rect 15012 10852 15068 10908
rect 15068 10852 15072 10908
rect 15008 10848 15072 10852
rect 15088 10908 15152 10912
rect 15088 10852 15092 10908
rect 15092 10852 15148 10908
rect 15148 10852 15152 10908
rect 15088 10848 15152 10852
rect 21796 10908 21860 10912
rect 21796 10852 21800 10908
rect 21800 10852 21856 10908
rect 21856 10852 21860 10908
rect 21796 10848 21860 10852
rect 21876 10908 21940 10912
rect 21876 10852 21880 10908
rect 21880 10852 21936 10908
rect 21936 10852 21940 10908
rect 21876 10848 21940 10852
rect 21956 10908 22020 10912
rect 21956 10852 21960 10908
rect 21960 10852 22016 10908
rect 22016 10852 22020 10908
rect 21956 10848 22020 10852
rect 22036 10908 22100 10912
rect 22036 10852 22040 10908
rect 22040 10852 22096 10908
rect 22096 10852 22100 10908
rect 22036 10848 22100 10852
rect 4426 10364 4490 10368
rect 4426 10308 4430 10364
rect 4430 10308 4486 10364
rect 4486 10308 4490 10364
rect 4426 10304 4490 10308
rect 4506 10364 4570 10368
rect 4506 10308 4510 10364
rect 4510 10308 4566 10364
rect 4566 10308 4570 10364
rect 4506 10304 4570 10308
rect 4586 10364 4650 10368
rect 4586 10308 4590 10364
rect 4590 10308 4646 10364
rect 4646 10308 4650 10364
rect 4586 10304 4650 10308
rect 4666 10364 4730 10368
rect 4666 10308 4670 10364
rect 4670 10308 4726 10364
rect 4726 10308 4730 10364
rect 4666 10304 4730 10308
rect 11374 10364 11438 10368
rect 11374 10308 11378 10364
rect 11378 10308 11434 10364
rect 11434 10308 11438 10364
rect 11374 10304 11438 10308
rect 11454 10364 11518 10368
rect 11454 10308 11458 10364
rect 11458 10308 11514 10364
rect 11514 10308 11518 10364
rect 11454 10304 11518 10308
rect 11534 10364 11598 10368
rect 11534 10308 11538 10364
rect 11538 10308 11594 10364
rect 11594 10308 11598 10364
rect 11534 10304 11598 10308
rect 11614 10364 11678 10368
rect 11614 10308 11618 10364
rect 11618 10308 11674 10364
rect 11674 10308 11678 10364
rect 11614 10304 11678 10308
rect 18322 10364 18386 10368
rect 18322 10308 18326 10364
rect 18326 10308 18382 10364
rect 18382 10308 18386 10364
rect 18322 10304 18386 10308
rect 18402 10364 18466 10368
rect 18402 10308 18406 10364
rect 18406 10308 18462 10364
rect 18462 10308 18466 10364
rect 18402 10304 18466 10308
rect 18482 10364 18546 10368
rect 18482 10308 18486 10364
rect 18486 10308 18542 10364
rect 18542 10308 18546 10364
rect 18482 10304 18546 10308
rect 18562 10364 18626 10368
rect 18562 10308 18566 10364
rect 18566 10308 18622 10364
rect 18622 10308 18626 10364
rect 18562 10304 18626 10308
rect 25270 10364 25334 10368
rect 25270 10308 25274 10364
rect 25274 10308 25330 10364
rect 25330 10308 25334 10364
rect 25270 10304 25334 10308
rect 25350 10364 25414 10368
rect 25350 10308 25354 10364
rect 25354 10308 25410 10364
rect 25410 10308 25414 10364
rect 25350 10304 25414 10308
rect 25430 10364 25494 10368
rect 25430 10308 25434 10364
rect 25434 10308 25490 10364
rect 25490 10308 25494 10364
rect 25430 10304 25494 10308
rect 25510 10364 25574 10368
rect 25510 10308 25514 10364
rect 25514 10308 25570 10364
rect 25570 10308 25574 10364
rect 25510 10304 25574 10308
rect 7900 9820 7964 9824
rect 7900 9764 7904 9820
rect 7904 9764 7960 9820
rect 7960 9764 7964 9820
rect 7900 9760 7964 9764
rect 7980 9820 8044 9824
rect 7980 9764 7984 9820
rect 7984 9764 8040 9820
rect 8040 9764 8044 9820
rect 7980 9760 8044 9764
rect 8060 9820 8124 9824
rect 8060 9764 8064 9820
rect 8064 9764 8120 9820
rect 8120 9764 8124 9820
rect 8060 9760 8124 9764
rect 8140 9820 8204 9824
rect 8140 9764 8144 9820
rect 8144 9764 8200 9820
rect 8200 9764 8204 9820
rect 8140 9760 8204 9764
rect 14848 9820 14912 9824
rect 14848 9764 14852 9820
rect 14852 9764 14908 9820
rect 14908 9764 14912 9820
rect 14848 9760 14912 9764
rect 14928 9820 14992 9824
rect 14928 9764 14932 9820
rect 14932 9764 14988 9820
rect 14988 9764 14992 9820
rect 14928 9760 14992 9764
rect 15008 9820 15072 9824
rect 15008 9764 15012 9820
rect 15012 9764 15068 9820
rect 15068 9764 15072 9820
rect 15008 9760 15072 9764
rect 15088 9820 15152 9824
rect 15088 9764 15092 9820
rect 15092 9764 15148 9820
rect 15148 9764 15152 9820
rect 15088 9760 15152 9764
rect 21796 9820 21860 9824
rect 21796 9764 21800 9820
rect 21800 9764 21856 9820
rect 21856 9764 21860 9820
rect 21796 9760 21860 9764
rect 21876 9820 21940 9824
rect 21876 9764 21880 9820
rect 21880 9764 21936 9820
rect 21936 9764 21940 9820
rect 21876 9760 21940 9764
rect 21956 9820 22020 9824
rect 21956 9764 21960 9820
rect 21960 9764 22016 9820
rect 22016 9764 22020 9820
rect 21956 9760 22020 9764
rect 22036 9820 22100 9824
rect 22036 9764 22040 9820
rect 22040 9764 22096 9820
rect 22096 9764 22100 9820
rect 22036 9760 22100 9764
rect 4426 9276 4490 9280
rect 4426 9220 4430 9276
rect 4430 9220 4486 9276
rect 4486 9220 4490 9276
rect 4426 9216 4490 9220
rect 4506 9276 4570 9280
rect 4506 9220 4510 9276
rect 4510 9220 4566 9276
rect 4566 9220 4570 9276
rect 4506 9216 4570 9220
rect 4586 9276 4650 9280
rect 4586 9220 4590 9276
rect 4590 9220 4646 9276
rect 4646 9220 4650 9276
rect 4586 9216 4650 9220
rect 4666 9276 4730 9280
rect 4666 9220 4670 9276
rect 4670 9220 4726 9276
rect 4726 9220 4730 9276
rect 4666 9216 4730 9220
rect 11374 9276 11438 9280
rect 11374 9220 11378 9276
rect 11378 9220 11434 9276
rect 11434 9220 11438 9276
rect 11374 9216 11438 9220
rect 11454 9276 11518 9280
rect 11454 9220 11458 9276
rect 11458 9220 11514 9276
rect 11514 9220 11518 9276
rect 11454 9216 11518 9220
rect 11534 9276 11598 9280
rect 11534 9220 11538 9276
rect 11538 9220 11594 9276
rect 11594 9220 11598 9276
rect 11534 9216 11598 9220
rect 11614 9276 11678 9280
rect 11614 9220 11618 9276
rect 11618 9220 11674 9276
rect 11674 9220 11678 9276
rect 11614 9216 11678 9220
rect 18322 9276 18386 9280
rect 18322 9220 18326 9276
rect 18326 9220 18382 9276
rect 18382 9220 18386 9276
rect 18322 9216 18386 9220
rect 18402 9276 18466 9280
rect 18402 9220 18406 9276
rect 18406 9220 18462 9276
rect 18462 9220 18466 9276
rect 18402 9216 18466 9220
rect 18482 9276 18546 9280
rect 18482 9220 18486 9276
rect 18486 9220 18542 9276
rect 18542 9220 18546 9276
rect 18482 9216 18546 9220
rect 18562 9276 18626 9280
rect 18562 9220 18566 9276
rect 18566 9220 18622 9276
rect 18622 9220 18626 9276
rect 18562 9216 18626 9220
rect 25270 9276 25334 9280
rect 25270 9220 25274 9276
rect 25274 9220 25330 9276
rect 25330 9220 25334 9276
rect 25270 9216 25334 9220
rect 25350 9276 25414 9280
rect 25350 9220 25354 9276
rect 25354 9220 25410 9276
rect 25410 9220 25414 9276
rect 25350 9216 25414 9220
rect 25430 9276 25494 9280
rect 25430 9220 25434 9276
rect 25434 9220 25490 9276
rect 25490 9220 25494 9276
rect 25430 9216 25494 9220
rect 25510 9276 25574 9280
rect 25510 9220 25514 9276
rect 25514 9220 25570 9276
rect 25570 9220 25574 9276
rect 25510 9216 25574 9220
rect 7900 8732 7964 8736
rect 7900 8676 7904 8732
rect 7904 8676 7960 8732
rect 7960 8676 7964 8732
rect 7900 8672 7964 8676
rect 7980 8732 8044 8736
rect 7980 8676 7984 8732
rect 7984 8676 8040 8732
rect 8040 8676 8044 8732
rect 7980 8672 8044 8676
rect 8060 8732 8124 8736
rect 8060 8676 8064 8732
rect 8064 8676 8120 8732
rect 8120 8676 8124 8732
rect 8060 8672 8124 8676
rect 8140 8732 8204 8736
rect 8140 8676 8144 8732
rect 8144 8676 8200 8732
rect 8200 8676 8204 8732
rect 8140 8672 8204 8676
rect 14848 8732 14912 8736
rect 14848 8676 14852 8732
rect 14852 8676 14908 8732
rect 14908 8676 14912 8732
rect 14848 8672 14912 8676
rect 14928 8732 14992 8736
rect 14928 8676 14932 8732
rect 14932 8676 14988 8732
rect 14988 8676 14992 8732
rect 14928 8672 14992 8676
rect 15008 8732 15072 8736
rect 15008 8676 15012 8732
rect 15012 8676 15068 8732
rect 15068 8676 15072 8732
rect 15008 8672 15072 8676
rect 15088 8732 15152 8736
rect 15088 8676 15092 8732
rect 15092 8676 15148 8732
rect 15148 8676 15152 8732
rect 15088 8672 15152 8676
rect 21796 8732 21860 8736
rect 21796 8676 21800 8732
rect 21800 8676 21856 8732
rect 21856 8676 21860 8732
rect 21796 8672 21860 8676
rect 21876 8732 21940 8736
rect 21876 8676 21880 8732
rect 21880 8676 21936 8732
rect 21936 8676 21940 8732
rect 21876 8672 21940 8676
rect 21956 8732 22020 8736
rect 21956 8676 21960 8732
rect 21960 8676 22016 8732
rect 22016 8676 22020 8732
rect 21956 8672 22020 8676
rect 22036 8732 22100 8736
rect 22036 8676 22040 8732
rect 22040 8676 22096 8732
rect 22096 8676 22100 8732
rect 22036 8672 22100 8676
rect 4426 8188 4490 8192
rect 4426 8132 4430 8188
rect 4430 8132 4486 8188
rect 4486 8132 4490 8188
rect 4426 8128 4490 8132
rect 4506 8188 4570 8192
rect 4506 8132 4510 8188
rect 4510 8132 4566 8188
rect 4566 8132 4570 8188
rect 4506 8128 4570 8132
rect 4586 8188 4650 8192
rect 4586 8132 4590 8188
rect 4590 8132 4646 8188
rect 4646 8132 4650 8188
rect 4586 8128 4650 8132
rect 4666 8188 4730 8192
rect 4666 8132 4670 8188
rect 4670 8132 4726 8188
rect 4726 8132 4730 8188
rect 4666 8128 4730 8132
rect 11374 8188 11438 8192
rect 11374 8132 11378 8188
rect 11378 8132 11434 8188
rect 11434 8132 11438 8188
rect 11374 8128 11438 8132
rect 11454 8188 11518 8192
rect 11454 8132 11458 8188
rect 11458 8132 11514 8188
rect 11514 8132 11518 8188
rect 11454 8128 11518 8132
rect 11534 8188 11598 8192
rect 11534 8132 11538 8188
rect 11538 8132 11594 8188
rect 11594 8132 11598 8188
rect 11534 8128 11598 8132
rect 11614 8188 11678 8192
rect 11614 8132 11618 8188
rect 11618 8132 11674 8188
rect 11674 8132 11678 8188
rect 11614 8128 11678 8132
rect 18322 8188 18386 8192
rect 18322 8132 18326 8188
rect 18326 8132 18382 8188
rect 18382 8132 18386 8188
rect 18322 8128 18386 8132
rect 18402 8188 18466 8192
rect 18402 8132 18406 8188
rect 18406 8132 18462 8188
rect 18462 8132 18466 8188
rect 18402 8128 18466 8132
rect 18482 8188 18546 8192
rect 18482 8132 18486 8188
rect 18486 8132 18542 8188
rect 18542 8132 18546 8188
rect 18482 8128 18546 8132
rect 18562 8188 18626 8192
rect 18562 8132 18566 8188
rect 18566 8132 18622 8188
rect 18622 8132 18626 8188
rect 18562 8128 18626 8132
rect 25270 8188 25334 8192
rect 25270 8132 25274 8188
rect 25274 8132 25330 8188
rect 25330 8132 25334 8188
rect 25270 8128 25334 8132
rect 25350 8188 25414 8192
rect 25350 8132 25354 8188
rect 25354 8132 25410 8188
rect 25410 8132 25414 8188
rect 25350 8128 25414 8132
rect 25430 8188 25494 8192
rect 25430 8132 25434 8188
rect 25434 8132 25490 8188
rect 25490 8132 25494 8188
rect 25430 8128 25494 8132
rect 25510 8188 25574 8192
rect 25510 8132 25514 8188
rect 25514 8132 25570 8188
rect 25570 8132 25574 8188
rect 25510 8128 25574 8132
rect 7900 7644 7964 7648
rect 7900 7588 7904 7644
rect 7904 7588 7960 7644
rect 7960 7588 7964 7644
rect 7900 7584 7964 7588
rect 7980 7644 8044 7648
rect 7980 7588 7984 7644
rect 7984 7588 8040 7644
rect 8040 7588 8044 7644
rect 7980 7584 8044 7588
rect 8060 7644 8124 7648
rect 8060 7588 8064 7644
rect 8064 7588 8120 7644
rect 8120 7588 8124 7644
rect 8060 7584 8124 7588
rect 8140 7644 8204 7648
rect 8140 7588 8144 7644
rect 8144 7588 8200 7644
rect 8200 7588 8204 7644
rect 8140 7584 8204 7588
rect 14848 7644 14912 7648
rect 14848 7588 14852 7644
rect 14852 7588 14908 7644
rect 14908 7588 14912 7644
rect 14848 7584 14912 7588
rect 14928 7644 14992 7648
rect 14928 7588 14932 7644
rect 14932 7588 14988 7644
rect 14988 7588 14992 7644
rect 14928 7584 14992 7588
rect 15008 7644 15072 7648
rect 15008 7588 15012 7644
rect 15012 7588 15068 7644
rect 15068 7588 15072 7644
rect 15008 7584 15072 7588
rect 15088 7644 15152 7648
rect 15088 7588 15092 7644
rect 15092 7588 15148 7644
rect 15148 7588 15152 7644
rect 15088 7584 15152 7588
rect 21796 7644 21860 7648
rect 21796 7588 21800 7644
rect 21800 7588 21856 7644
rect 21856 7588 21860 7644
rect 21796 7584 21860 7588
rect 21876 7644 21940 7648
rect 21876 7588 21880 7644
rect 21880 7588 21936 7644
rect 21936 7588 21940 7644
rect 21876 7584 21940 7588
rect 21956 7644 22020 7648
rect 21956 7588 21960 7644
rect 21960 7588 22016 7644
rect 22016 7588 22020 7644
rect 21956 7584 22020 7588
rect 22036 7644 22100 7648
rect 22036 7588 22040 7644
rect 22040 7588 22096 7644
rect 22096 7588 22100 7644
rect 22036 7584 22100 7588
rect 4426 7100 4490 7104
rect 4426 7044 4430 7100
rect 4430 7044 4486 7100
rect 4486 7044 4490 7100
rect 4426 7040 4490 7044
rect 4506 7100 4570 7104
rect 4506 7044 4510 7100
rect 4510 7044 4566 7100
rect 4566 7044 4570 7100
rect 4506 7040 4570 7044
rect 4586 7100 4650 7104
rect 4586 7044 4590 7100
rect 4590 7044 4646 7100
rect 4646 7044 4650 7100
rect 4586 7040 4650 7044
rect 4666 7100 4730 7104
rect 4666 7044 4670 7100
rect 4670 7044 4726 7100
rect 4726 7044 4730 7100
rect 4666 7040 4730 7044
rect 11374 7100 11438 7104
rect 11374 7044 11378 7100
rect 11378 7044 11434 7100
rect 11434 7044 11438 7100
rect 11374 7040 11438 7044
rect 11454 7100 11518 7104
rect 11454 7044 11458 7100
rect 11458 7044 11514 7100
rect 11514 7044 11518 7100
rect 11454 7040 11518 7044
rect 11534 7100 11598 7104
rect 11534 7044 11538 7100
rect 11538 7044 11594 7100
rect 11594 7044 11598 7100
rect 11534 7040 11598 7044
rect 11614 7100 11678 7104
rect 11614 7044 11618 7100
rect 11618 7044 11674 7100
rect 11674 7044 11678 7100
rect 11614 7040 11678 7044
rect 18322 7100 18386 7104
rect 18322 7044 18326 7100
rect 18326 7044 18382 7100
rect 18382 7044 18386 7100
rect 18322 7040 18386 7044
rect 18402 7100 18466 7104
rect 18402 7044 18406 7100
rect 18406 7044 18462 7100
rect 18462 7044 18466 7100
rect 18402 7040 18466 7044
rect 18482 7100 18546 7104
rect 18482 7044 18486 7100
rect 18486 7044 18542 7100
rect 18542 7044 18546 7100
rect 18482 7040 18546 7044
rect 18562 7100 18626 7104
rect 18562 7044 18566 7100
rect 18566 7044 18622 7100
rect 18622 7044 18626 7100
rect 18562 7040 18626 7044
rect 25270 7100 25334 7104
rect 25270 7044 25274 7100
rect 25274 7044 25330 7100
rect 25330 7044 25334 7100
rect 25270 7040 25334 7044
rect 25350 7100 25414 7104
rect 25350 7044 25354 7100
rect 25354 7044 25410 7100
rect 25410 7044 25414 7100
rect 25350 7040 25414 7044
rect 25430 7100 25494 7104
rect 25430 7044 25434 7100
rect 25434 7044 25490 7100
rect 25490 7044 25494 7100
rect 25430 7040 25494 7044
rect 25510 7100 25574 7104
rect 25510 7044 25514 7100
rect 25514 7044 25570 7100
rect 25570 7044 25574 7100
rect 25510 7040 25574 7044
rect 7900 6556 7964 6560
rect 7900 6500 7904 6556
rect 7904 6500 7960 6556
rect 7960 6500 7964 6556
rect 7900 6496 7964 6500
rect 7980 6556 8044 6560
rect 7980 6500 7984 6556
rect 7984 6500 8040 6556
rect 8040 6500 8044 6556
rect 7980 6496 8044 6500
rect 8060 6556 8124 6560
rect 8060 6500 8064 6556
rect 8064 6500 8120 6556
rect 8120 6500 8124 6556
rect 8060 6496 8124 6500
rect 8140 6556 8204 6560
rect 8140 6500 8144 6556
rect 8144 6500 8200 6556
rect 8200 6500 8204 6556
rect 8140 6496 8204 6500
rect 14848 6556 14912 6560
rect 14848 6500 14852 6556
rect 14852 6500 14908 6556
rect 14908 6500 14912 6556
rect 14848 6496 14912 6500
rect 14928 6556 14992 6560
rect 14928 6500 14932 6556
rect 14932 6500 14988 6556
rect 14988 6500 14992 6556
rect 14928 6496 14992 6500
rect 15008 6556 15072 6560
rect 15008 6500 15012 6556
rect 15012 6500 15068 6556
rect 15068 6500 15072 6556
rect 15008 6496 15072 6500
rect 15088 6556 15152 6560
rect 15088 6500 15092 6556
rect 15092 6500 15148 6556
rect 15148 6500 15152 6556
rect 15088 6496 15152 6500
rect 21796 6556 21860 6560
rect 21796 6500 21800 6556
rect 21800 6500 21856 6556
rect 21856 6500 21860 6556
rect 21796 6496 21860 6500
rect 21876 6556 21940 6560
rect 21876 6500 21880 6556
rect 21880 6500 21936 6556
rect 21936 6500 21940 6556
rect 21876 6496 21940 6500
rect 21956 6556 22020 6560
rect 21956 6500 21960 6556
rect 21960 6500 22016 6556
rect 22016 6500 22020 6556
rect 21956 6496 22020 6500
rect 22036 6556 22100 6560
rect 22036 6500 22040 6556
rect 22040 6500 22096 6556
rect 22096 6500 22100 6556
rect 22036 6496 22100 6500
rect 4426 6012 4490 6016
rect 4426 5956 4430 6012
rect 4430 5956 4486 6012
rect 4486 5956 4490 6012
rect 4426 5952 4490 5956
rect 4506 6012 4570 6016
rect 4506 5956 4510 6012
rect 4510 5956 4566 6012
rect 4566 5956 4570 6012
rect 4506 5952 4570 5956
rect 4586 6012 4650 6016
rect 4586 5956 4590 6012
rect 4590 5956 4646 6012
rect 4646 5956 4650 6012
rect 4586 5952 4650 5956
rect 4666 6012 4730 6016
rect 4666 5956 4670 6012
rect 4670 5956 4726 6012
rect 4726 5956 4730 6012
rect 4666 5952 4730 5956
rect 11374 6012 11438 6016
rect 11374 5956 11378 6012
rect 11378 5956 11434 6012
rect 11434 5956 11438 6012
rect 11374 5952 11438 5956
rect 11454 6012 11518 6016
rect 11454 5956 11458 6012
rect 11458 5956 11514 6012
rect 11514 5956 11518 6012
rect 11454 5952 11518 5956
rect 11534 6012 11598 6016
rect 11534 5956 11538 6012
rect 11538 5956 11594 6012
rect 11594 5956 11598 6012
rect 11534 5952 11598 5956
rect 11614 6012 11678 6016
rect 11614 5956 11618 6012
rect 11618 5956 11674 6012
rect 11674 5956 11678 6012
rect 11614 5952 11678 5956
rect 18322 6012 18386 6016
rect 18322 5956 18326 6012
rect 18326 5956 18382 6012
rect 18382 5956 18386 6012
rect 18322 5952 18386 5956
rect 18402 6012 18466 6016
rect 18402 5956 18406 6012
rect 18406 5956 18462 6012
rect 18462 5956 18466 6012
rect 18402 5952 18466 5956
rect 18482 6012 18546 6016
rect 18482 5956 18486 6012
rect 18486 5956 18542 6012
rect 18542 5956 18546 6012
rect 18482 5952 18546 5956
rect 18562 6012 18626 6016
rect 18562 5956 18566 6012
rect 18566 5956 18622 6012
rect 18622 5956 18626 6012
rect 18562 5952 18626 5956
rect 25270 6012 25334 6016
rect 25270 5956 25274 6012
rect 25274 5956 25330 6012
rect 25330 5956 25334 6012
rect 25270 5952 25334 5956
rect 25350 6012 25414 6016
rect 25350 5956 25354 6012
rect 25354 5956 25410 6012
rect 25410 5956 25414 6012
rect 25350 5952 25414 5956
rect 25430 6012 25494 6016
rect 25430 5956 25434 6012
rect 25434 5956 25490 6012
rect 25490 5956 25494 6012
rect 25430 5952 25494 5956
rect 25510 6012 25574 6016
rect 25510 5956 25514 6012
rect 25514 5956 25570 6012
rect 25570 5956 25574 6012
rect 25510 5952 25574 5956
rect 7900 5468 7964 5472
rect 7900 5412 7904 5468
rect 7904 5412 7960 5468
rect 7960 5412 7964 5468
rect 7900 5408 7964 5412
rect 7980 5468 8044 5472
rect 7980 5412 7984 5468
rect 7984 5412 8040 5468
rect 8040 5412 8044 5468
rect 7980 5408 8044 5412
rect 8060 5468 8124 5472
rect 8060 5412 8064 5468
rect 8064 5412 8120 5468
rect 8120 5412 8124 5468
rect 8060 5408 8124 5412
rect 8140 5468 8204 5472
rect 8140 5412 8144 5468
rect 8144 5412 8200 5468
rect 8200 5412 8204 5468
rect 8140 5408 8204 5412
rect 14848 5468 14912 5472
rect 14848 5412 14852 5468
rect 14852 5412 14908 5468
rect 14908 5412 14912 5468
rect 14848 5408 14912 5412
rect 14928 5468 14992 5472
rect 14928 5412 14932 5468
rect 14932 5412 14988 5468
rect 14988 5412 14992 5468
rect 14928 5408 14992 5412
rect 15008 5468 15072 5472
rect 15008 5412 15012 5468
rect 15012 5412 15068 5468
rect 15068 5412 15072 5468
rect 15008 5408 15072 5412
rect 15088 5468 15152 5472
rect 15088 5412 15092 5468
rect 15092 5412 15148 5468
rect 15148 5412 15152 5468
rect 15088 5408 15152 5412
rect 21796 5468 21860 5472
rect 21796 5412 21800 5468
rect 21800 5412 21856 5468
rect 21856 5412 21860 5468
rect 21796 5408 21860 5412
rect 21876 5468 21940 5472
rect 21876 5412 21880 5468
rect 21880 5412 21936 5468
rect 21936 5412 21940 5468
rect 21876 5408 21940 5412
rect 21956 5468 22020 5472
rect 21956 5412 21960 5468
rect 21960 5412 22016 5468
rect 22016 5412 22020 5468
rect 21956 5408 22020 5412
rect 22036 5468 22100 5472
rect 22036 5412 22040 5468
rect 22040 5412 22096 5468
rect 22096 5412 22100 5468
rect 22036 5408 22100 5412
rect 4426 4924 4490 4928
rect 4426 4868 4430 4924
rect 4430 4868 4486 4924
rect 4486 4868 4490 4924
rect 4426 4864 4490 4868
rect 4506 4924 4570 4928
rect 4506 4868 4510 4924
rect 4510 4868 4566 4924
rect 4566 4868 4570 4924
rect 4506 4864 4570 4868
rect 4586 4924 4650 4928
rect 4586 4868 4590 4924
rect 4590 4868 4646 4924
rect 4646 4868 4650 4924
rect 4586 4864 4650 4868
rect 4666 4924 4730 4928
rect 4666 4868 4670 4924
rect 4670 4868 4726 4924
rect 4726 4868 4730 4924
rect 4666 4864 4730 4868
rect 11374 4924 11438 4928
rect 11374 4868 11378 4924
rect 11378 4868 11434 4924
rect 11434 4868 11438 4924
rect 11374 4864 11438 4868
rect 11454 4924 11518 4928
rect 11454 4868 11458 4924
rect 11458 4868 11514 4924
rect 11514 4868 11518 4924
rect 11454 4864 11518 4868
rect 11534 4924 11598 4928
rect 11534 4868 11538 4924
rect 11538 4868 11594 4924
rect 11594 4868 11598 4924
rect 11534 4864 11598 4868
rect 11614 4924 11678 4928
rect 11614 4868 11618 4924
rect 11618 4868 11674 4924
rect 11674 4868 11678 4924
rect 11614 4864 11678 4868
rect 18322 4924 18386 4928
rect 18322 4868 18326 4924
rect 18326 4868 18382 4924
rect 18382 4868 18386 4924
rect 18322 4864 18386 4868
rect 18402 4924 18466 4928
rect 18402 4868 18406 4924
rect 18406 4868 18462 4924
rect 18462 4868 18466 4924
rect 18402 4864 18466 4868
rect 18482 4924 18546 4928
rect 18482 4868 18486 4924
rect 18486 4868 18542 4924
rect 18542 4868 18546 4924
rect 18482 4864 18546 4868
rect 18562 4924 18626 4928
rect 18562 4868 18566 4924
rect 18566 4868 18622 4924
rect 18622 4868 18626 4924
rect 18562 4864 18626 4868
rect 25270 4924 25334 4928
rect 25270 4868 25274 4924
rect 25274 4868 25330 4924
rect 25330 4868 25334 4924
rect 25270 4864 25334 4868
rect 25350 4924 25414 4928
rect 25350 4868 25354 4924
rect 25354 4868 25410 4924
rect 25410 4868 25414 4924
rect 25350 4864 25414 4868
rect 25430 4924 25494 4928
rect 25430 4868 25434 4924
rect 25434 4868 25490 4924
rect 25490 4868 25494 4924
rect 25430 4864 25494 4868
rect 25510 4924 25574 4928
rect 25510 4868 25514 4924
rect 25514 4868 25570 4924
rect 25570 4868 25574 4924
rect 25510 4864 25574 4868
rect 7900 4380 7964 4384
rect 7900 4324 7904 4380
rect 7904 4324 7960 4380
rect 7960 4324 7964 4380
rect 7900 4320 7964 4324
rect 7980 4380 8044 4384
rect 7980 4324 7984 4380
rect 7984 4324 8040 4380
rect 8040 4324 8044 4380
rect 7980 4320 8044 4324
rect 8060 4380 8124 4384
rect 8060 4324 8064 4380
rect 8064 4324 8120 4380
rect 8120 4324 8124 4380
rect 8060 4320 8124 4324
rect 8140 4380 8204 4384
rect 8140 4324 8144 4380
rect 8144 4324 8200 4380
rect 8200 4324 8204 4380
rect 8140 4320 8204 4324
rect 14848 4380 14912 4384
rect 14848 4324 14852 4380
rect 14852 4324 14908 4380
rect 14908 4324 14912 4380
rect 14848 4320 14912 4324
rect 14928 4380 14992 4384
rect 14928 4324 14932 4380
rect 14932 4324 14988 4380
rect 14988 4324 14992 4380
rect 14928 4320 14992 4324
rect 15008 4380 15072 4384
rect 15008 4324 15012 4380
rect 15012 4324 15068 4380
rect 15068 4324 15072 4380
rect 15008 4320 15072 4324
rect 15088 4380 15152 4384
rect 15088 4324 15092 4380
rect 15092 4324 15148 4380
rect 15148 4324 15152 4380
rect 15088 4320 15152 4324
rect 21796 4380 21860 4384
rect 21796 4324 21800 4380
rect 21800 4324 21856 4380
rect 21856 4324 21860 4380
rect 21796 4320 21860 4324
rect 21876 4380 21940 4384
rect 21876 4324 21880 4380
rect 21880 4324 21936 4380
rect 21936 4324 21940 4380
rect 21876 4320 21940 4324
rect 21956 4380 22020 4384
rect 21956 4324 21960 4380
rect 21960 4324 22016 4380
rect 22016 4324 22020 4380
rect 21956 4320 22020 4324
rect 22036 4380 22100 4384
rect 22036 4324 22040 4380
rect 22040 4324 22096 4380
rect 22096 4324 22100 4380
rect 22036 4320 22100 4324
rect 4426 3836 4490 3840
rect 4426 3780 4430 3836
rect 4430 3780 4486 3836
rect 4486 3780 4490 3836
rect 4426 3776 4490 3780
rect 4506 3836 4570 3840
rect 4506 3780 4510 3836
rect 4510 3780 4566 3836
rect 4566 3780 4570 3836
rect 4506 3776 4570 3780
rect 4586 3836 4650 3840
rect 4586 3780 4590 3836
rect 4590 3780 4646 3836
rect 4646 3780 4650 3836
rect 4586 3776 4650 3780
rect 4666 3836 4730 3840
rect 4666 3780 4670 3836
rect 4670 3780 4726 3836
rect 4726 3780 4730 3836
rect 4666 3776 4730 3780
rect 11374 3836 11438 3840
rect 11374 3780 11378 3836
rect 11378 3780 11434 3836
rect 11434 3780 11438 3836
rect 11374 3776 11438 3780
rect 11454 3836 11518 3840
rect 11454 3780 11458 3836
rect 11458 3780 11514 3836
rect 11514 3780 11518 3836
rect 11454 3776 11518 3780
rect 11534 3836 11598 3840
rect 11534 3780 11538 3836
rect 11538 3780 11594 3836
rect 11594 3780 11598 3836
rect 11534 3776 11598 3780
rect 11614 3836 11678 3840
rect 11614 3780 11618 3836
rect 11618 3780 11674 3836
rect 11674 3780 11678 3836
rect 11614 3776 11678 3780
rect 18322 3836 18386 3840
rect 18322 3780 18326 3836
rect 18326 3780 18382 3836
rect 18382 3780 18386 3836
rect 18322 3776 18386 3780
rect 18402 3836 18466 3840
rect 18402 3780 18406 3836
rect 18406 3780 18462 3836
rect 18462 3780 18466 3836
rect 18402 3776 18466 3780
rect 18482 3836 18546 3840
rect 18482 3780 18486 3836
rect 18486 3780 18542 3836
rect 18542 3780 18546 3836
rect 18482 3776 18546 3780
rect 18562 3836 18626 3840
rect 18562 3780 18566 3836
rect 18566 3780 18622 3836
rect 18622 3780 18626 3836
rect 18562 3776 18626 3780
rect 25270 3836 25334 3840
rect 25270 3780 25274 3836
rect 25274 3780 25330 3836
rect 25330 3780 25334 3836
rect 25270 3776 25334 3780
rect 25350 3836 25414 3840
rect 25350 3780 25354 3836
rect 25354 3780 25410 3836
rect 25410 3780 25414 3836
rect 25350 3776 25414 3780
rect 25430 3836 25494 3840
rect 25430 3780 25434 3836
rect 25434 3780 25490 3836
rect 25490 3780 25494 3836
rect 25430 3776 25494 3780
rect 25510 3836 25574 3840
rect 25510 3780 25514 3836
rect 25514 3780 25570 3836
rect 25570 3780 25574 3836
rect 25510 3776 25574 3780
rect 7900 3292 7964 3296
rect 7900 3236 7904 3292
rect 7904 3236 7960 3292
rect 7960 3236 7964 3292
rect 7900 3232 7964 3236
rect 7980 3292 8044 3296
rect 7980 3236 7984 3292
rect 7984 3236 8040 3292
rect 8040 3236 8044 3292
rect 7980 3232 8044 3236
rect 8060 3292 8124 3296
rect 8060 3236 8064 3292
rect 8064 3236 8120 3292
rect 8120 3236 8124 3292
rect 8060 3232 8124 3236
rect 8140 3292 8204 3296
rect 8140 3236 8144 3292
rect 8144 3236 8200 3292
rect 8200 3236 8204 3292
rect 8140 3232 8204 3236
rect 14848 3292 14912 3296
rect 14848 3236 14852 3292
rect 14852 3236 14908 3292
rect 14908 3236 14912 3292
rect 14848 3232 14912 3236
rect 14928 3292 14992 3296
rect 14928 3236 14932 3292
rect 14932 3236 14988 3292
rect 14988 3236 14992 3292
rect 14928 3232 14992 3236
rect 15008 3292 15072 3296
rect 15008 3236 15012 3292
rect 15012 3236 15068 3292
rect 15068 3236 15072 3292
rect 15008 3232 15072 3236
rect 15088 3292 15152 3296
rect 15088 3236 15092 3292
rect 15092 3236 15148 3292
rect 15148 3236 15152 3292
rect 15088 3232 15152 3236
rect 21796 3292 21860 3296
rect 21796 3236 21800 3292
rect 21800 3236 21856 3292
rect 21856 3236 21860 3292
rect 21796 3232 21860 3236
rect 21876 3292 21940 3296
rect 21876 3236 21880 3292
rect 21880 3236 21936 3292
rect 21936 3236 21940 3292
rect 21876 3232 21940 3236
rect 21956 3292 22020 3296
rect 21956 3236 21960 3292
rect 21960 3236 22016 3292
rect 22016 3236 22020 3292
rect 21956 3232 22020 3236
rect 22036 3292 22100 3296
rect 22036 3236 22040 3292
rect 22040 3236 22096 3292
rect 22096 3236 22100 3292
rect 22036 3232 22100 3236
rect 4426 2748 4490 2752
rect 4426 2692 4430 2748
rect 4430 2692 4486 2748
rect 4486 2692 4490 2748
rect 4426 2688 4490 2692
rect 4506 2748 4570 2752
rect 4506 2692 4510 2748
rect 4510 2692 4566 2748
rect 4566 2692 4570 2748
rect 4506 2688 4570 2692
rect 4586 2748 4650 2752
rect 4586 2692 4590 2748
rect 4590 2692 4646 2748
rect 4646 2692 4650 2748
rect 4586 2688 4650 2692
rect 4666 2748 4730 2752
rect 4666 2692 4670 2748
rect 4670 2692 4726 2748
rect 4726 2692 4730 2748
rect 4666 2688 4730 2692
rect 11374 2748 11438 2752
rect 11374 2692 11378 2748
rect 11378 2692 11434 2748
rect 11434 2692 11438 2748
rect 11374 2688 11438 2692
rect 11454 2748 11518 2752
rect 11454 2692 11458 2748
rect 11458 2692 11514 2748
rect 11514 2692 11518 2748
rect 11454 2688 11518 2692
rect 11534 2748 11598 2752
rect 11534 2692 11538 2748
rect 11538 2692 11594 2748
rect 11594 2692 11598 2748
rect 11534 2688 11598 2692
rect 11614 2748 11678 2752
rect 11614 2692 11618 2748
rect 11618 2692 11674 2748
rect 11674 2692 11678 2748
rect 11614 2688 11678 2692
rect 18322 2748 18386 2752
rect 18322 2692 18326 2748
rect 18326 2692 18382 2748
rect 18382 2692 18386 2748
rect 18322 2688 18386 2692
rect 18402 2748 18466 2752
rect 18402 2692 18406 2748
rect 18406 2692 18462 2748
rect 18462 2692 18466 2748
rect 18402 2688 18466 2692
rect 18482 2748 18546 2752
rect 18482 2692 18486 2748
rect 18486 2692 18542 2748
rect 18542 2692 18546 2748
rect 18482 2688 18546 2692
rect 18562 2748 18626 2752
rect 18562 2692 18566 2748
rect 18566 2692 18622 2748
rect 18622 2692 18626 2748
rect 18562 2688 18626 2692
rect 25270 2748 25334 2752
rect 25270 2692 25274 2748
rect 25274 2692 25330 2748
rect 25330 2692 25334 2748
rect 25270 2688 25334 2692
rect 25350 2748 25414 2752
rect 25350 2692 25354 2748
rect 25354 2692 25410 2748
rect 25410 2692 25414 2748
rect 25350 2688 25414 2692
rect 25430 2748 25494 2752
rect 25430 2692 25434 2748
rect 25434 2692 25490 2748
rect 25490 2692 25494 2748
rect 25430 2688 25494 2692
rect 25510 2748 25574 2752
rect 25510 2692 25514 2748
rect 25514 2692 25570 2748
rect 25570 2692 25574 2748
rect 25510 2688 25574 2692
rect 7900 2204 7964 2208
rect 7900 2148 7904 2204
rect 7904 2148 7960 2204
rect 7960 2148 7964 2204
rect 7900 2144 7964 2148
rect 7980 2204 8044 2208
rect 7980 2148 7984 2204
rect 7984 2148 8040 2204
rect 8040 2148 8044 2204
rect 7980 2144 8044 2148
rect 8060 2204 8124 2208
rect 8060 2148 8064 2204
rect 8064 2148 8120 2204
rect 8120 2148 8124 2204
rect 8060 2144 8124 2148
rect 8140 2204 8204 2208
rect 8140 2148 8144 2204
rect 8144 2148 8200 2204
rect 8200 2148 8204 2204
rect 8140 2144 8204 2148
rect 14848 2204 14912 2208
rect 14848 2148 14852 2204
rect 14852 2148 14908 2204
rect 14908 2148 14912 2204
rect 14848 2144 14912 2148
rect 14928 2204 14992 2208
rect 14928 2148 14932 2204
rect 14932 2148 14988 2204
rect 14988 2148 14992 2204
rect 14928 2144 14992 2148
rect 15008 2204 15072 2208
rect 15008 2148 15012 2204
rect 15012 2148 15068 2204
rect 15068 2148 15072 2204
rect 15008 2144 15072 2148
rect 15088 2204 15152 2208
rect 15088 2148 15092 2204
rect 15092 2148 15148 2204
rect 15148 2148 15152 2204
rect 15088 2144 15152 2148
rect 21796 2204 21860 2208
rect 21796 2148 21800 2204
rect 21800 2148 21856 2204
rect 21856 2148 21860 2204
rect 21796 2144 21860 2148
rect 21876 2204 21940 2208
rect 21876 2148 21880 2204
rect 21880 2148 21936 2204
rect 21936 2148 21940 2204
rect 21876 2144 21940 2148
rect 21956 2204 22020 2208
rect 21956 2148 21960 2204
rect 21960 2148 22016 2204
rect 22016 2148 22020 2204
rect 21956 2144 22020 2148
rect 22036 2204 22100 2208
rect 22036 2148 22040 2204
rect 22040 2148 22096 2204
rect 22096 2148 22100 2204
rect 22036 2144 22100 2148
<< metal4 >>
rect 4418 27776 4738 27792
rect 4418 27712 4426 27776
rect 4490 27712 4506 27776
rect 4570 27712 4586 27776
rect 4650 27712 4666 27776
rect 4730 27712 4738 27776
rect 4418 26688 4738 27712
rect 4418 26624 4426 26688
rect 4490 26624 4506 26688
rect 4570 26624 4586 26688
rect 4650 26624 4666 26688
rect 4730 26624 4738 26688
rect 4418 25600 4738 26624
rect 4418 25536 4426 25600
rect 4490 25536 4506 25600
rect 4570 25536 4586 25600
rect 4650 25536 4666 25600
rect 4730 25536 4738 25600
rect 4418 24512 4738 25536
rect 4418 24448 4426 24512
rect 4490 24448 4506 24512
rect 4570 24448 4586 24512
rect 4650 24448 4666 24512
rect 4730 24448 4738 24512
rect 4418 23424 4738 24448
rect 4418 23360 4426 23424
rect 4490 23360 4506 23424
rect 4570 23360 4586 23424
rect 4650 23360 4666 23424
rect 4730 23360 4738 23424
rect 4418 22336 4738 23360
rect 4418 22272 4426 22336
rect 4490 22272 4506 22336
rect 4570 22272 4586 22336
rect 4650 22272 4666 22336
rect 4730 22272 4738 22336
rect 4418 21248 4738 22272
rect 4418 21184 4426 21248
rect 4490 21184 4506 21248
rect 4570 21184 4586 21248
rect 4650 21184 4666 21248
rect 4730 21184 4738 21248
rect 4418 20160 4738 21184
rect 4418 20096 4426 20160
rect 4490 20096 4506 20160
rect 4570 20096 4586 20160
rect 4650 20096 4666 20160
rect 4730 20096 4738 20160
rect 4418 19072 4738 20096
rect 4418 19008 4426 19072
rect 4490 19008 4506 19072
rect 4570 19008 4586 19072
rect 4650 19008 4666 19072
rect 4730 19008 4738 19072
rect 4418 17984 4738 19008
rect 4418 17920 4426 17984
rect 4490 17920 4506 17984
rect 4570 17920 4586 17984
rect 4650 17920 4666 17984
rect 4730 17920 4738 17984
rect 4418 16896 4738 17920
rect 4418 16832 4426 16896
rect 4490 16832 4506 16896
rect 4570 16832 4586 16896
rect 4650 16832 4666 16896
rect 4730 16832 4738 16896
rect 4418 15808 4738 16832
rect 4418 15744 4426 15808
rect 4490 15744 4506 15808
rect 4570 15744 4586 15808
rect 4650 15744 4666 15808
rect 4730 15744 4738 15808
rect 4418 14720 4738 15744
rect 4418 14656 4426 14720
rect 4490 14656 4506 14720
rect 4570 14656 4586 14720
rect 4650 14656 4666 14720
rect 4730 14656 4738 14720
rect 4418 13632 4738 14656
rect 4418 13568 4426 13632
rect 4490 13568 4506 13632
rect 4570 13568 4586 13632
rect 4650 13568 4666 13632
rect 4730 13568 4738 13632
rect 4418 12544 4738 13568
rect 4418 12480 4426 12544
rect 4490 12480 4506 12544
rect 4570 12480 4586 12544
rect 4650 12480 4666 12544
rect 4730 12480 4738 12544
rect 4418 11456 4738 12480
rect 4418 11392 4426 11456
rect 4490 11392 4506 11456
rect 4570 11392 4586 11456
rect 4650 11392 4666 11456
rect 4730 11392 4738 11456
rect 4418 10368 4738 11392
rect 4418 10304 4426 10368
rect 4490 10304 4506 10368
rect 4570 10304 4586 10368
rect 4650 10304 4666 10368
rect 4730 10304 4738 10368
rect 4418 9280 4738 10304
rect 4418 9216 4426 9280
rect 4490 9216 4506 9280
rect 4570 9216 4586 9280
rect 4650 9216 4666 9280
rect 4730 9216 4738 9280
rect 4418 8192 4738 9216
rect 4418 8128 4426 8192
rect 4490 8128 4506 8192
rect 4570 8128 4586 8192
rect 4650 8128 4666 8192
rect 4730 8128 4738 8192
rect 4418 7104 4738 8128
rect 4418 7040 4426 7104
rect 4490 7040 4506 7104
rect 4570 7040 4586 7104
rect 4650 7040 4666 7104
rect 4730 7040 4738 7104
rect 4418 6016 4738 7040
rect 4418 5952 4426 6016
rect 4490 5952 4506 6016
rect 4570 5952 4586 6016
rect 4650 5952 4666 6016
rect 4730 5952 4738 6016
rect 4418 4928 4738 5952
rect 4418 4864 4426 4928
rect 4490 4864 4506 4928
rect 4570 4864 4586 4928
rect 4650 4864 4666 4928
rect 4730 4864 4738 4928
rect 4418 3840 4738 4864
rect 4418 3776 4426 3840
rect 4490 3776 4506 3840
rect 4570 3776 4586 3840
rect 4650 3776 4666 3840
rect 4730 3776 4738 3840
rect 4418 2752 4738 3776
rect 4418 2688 4426 2752
rect 4490 2688 4506 2752
rect 4570 2688 4586 2752
rect 4650 2688 4666 2752
rect 4730 2688 4738 2752
rect 4418 2128 4738 2688
rect 7892 27232 8212 27792
rect 7892 27168 7900 27232
rect 7964 27168 7980 27232
rect 8044 27168 8060 27232
rect 8124 27168 8140 27232
rect 8204 27168 8212 27232
rect 7892 26144 8212 27168
rect 7892 26080 7900 26144
rect 7964 26080 7980 26144
rect 8044 26080 8060 26144
rect 8124 26080 8140 26144
rect 8204 26080 8212 26144
rect 7892 25056 8212 26080
rect 7892 24992 7900 25056
rect 7964 24992 7980 25056
rect 8044 24992 8060 25056
rect 8124 24992 8140 25056
rect 8204 24992 8212 25056
rect 7892 23968 8212 24992
rect 7892 23904 7900 23968
rect 7964 23904 7980 23968
rect 8044 23904 8060 23968
rect 8124 23904 8140 23968
rect 8204 23904 8212 23968
rect 7892 22880 8212 23904
rect 7892 22816 7900 22880
rect 7964 22816 7980 22880
rect 8044 22816 8060 22880
rect 8124 22816 8140 22880
rect 8204 22816 8212 22880
rect 7892 21792 8212 22816
rect 7892 21728 7900 21792
rect 7964 21728 7980 21792
rect 8044 21728 8060 21792
rect 8124 21728 8140 21792
rect 8204 21728 8212 21792
rect 7892 20704 8212 21728
rect 7892 20640 7900 20704
rect 7964 20640 7980 20704
rect 8044 20640 8060 20704
rect 8124 20640 8140 20704
rect 8204 20640 8212 20704
rect 7892 19616 8212 20640
rect 7892 19552 7900 19616
rect 7964 19552 7980 19616
rect 8044 19552 8060 19616
rect 8124 19552 8140 19616
rect 8204 19552 8212 19616
rect 7892 18528 8212 19552
rect 7892 18464 7900 18528
rect 7964 18464 7980 18528
rect 8044 18464 8060 18528
rect 8124 18464 8140 18528
rect 8204 18464 8212 18528
rect 7892 17440 8212 18464
rect 7892 17376 7900 17440
rect 7964 17376 7980 17440
rect 8044 17376 8060 17440
rect 8124 17376 8140 17440
rect 8204 17376 8212 17440
rect 7892 16352 8212 17376
rect 7892 16288 7900 16352
rect 7964 16288 7980 16352
rect 8044 16288 8060 16352
rect 8124 16288 8140 16352
rect 8204 16288 8212 16352
rect 7892 15264 8212 16288
rect 7892 15200 7900 15264
rect 7964 15200 7980 15264
rect 8044 15200 8060 15264
rect 8124 15200 8140 15264
rect 8204 15200 8212 15264
rect 7892 14176 8212 15200
rect 7892 14112 7900 14176
rect 7964 14112 7980 14176
rect 8044 14112 8060 14176
rect 8124 14112 8140 14176
rect 8204 14112 8212 14176
rect 7892 13088 8212 14112
rect 7892 13024 7900 13088
rect 7964 13024 7980 13088
rect 8044 13024 8060 13088
rect 8124 13024 8140 13088
rect 8204 13024 8212 13088
rect 7892 12000 8212 13024
rect 7892 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8212 12000
rect 7892 10912 8212 11936
rect 7892 10848 7900 10912
rect 7964 10848 7980 10912
rect 8044 10848 8060 10912
rect 8124 10848 8140 10912
rect 8204 10848 8212 10912
rect 7892 9824 8212 10848
rect 7892 9760 7900 9824
rect 7964 9760 7980 9824
rect 8044 9760 8060 9824
rect 8124 9760 8140 9824
rect 8204 9760 8212 9824
rect 7892 8736 8212 9760
rect 7892 8672 7900 8736
rect 7964 8672 7980 8736
rect 8044 8672 8060 8736
rect 8124 8672 8140 8736
rect 8204 8672 8212 8736
rect 7892 7648 8212 8672
rect 7892 7584 7900 7648
rect 7964 7584 7980 7648
rect 8044 7584 8060 7648
rect 8124 7584 8140 7648
rect 8204 7584 8212 7648
rect 7892 6560 8212 7584
rect 7892 6496 7900 6560
rect 7964 6496 7980 6560
rect 8044 6496 8060 6560
rect 8124 6496 8140 6560
rect 8204 6496 8212 6560
rect 7892 5472 8212 6496
rect 7892 5408 7900 5472
rect 7964 5408 7980 5472
rect 8044 5408 8060 5472
rect 8124 5408 8140 5472
rect 8204 5408 8212 5472
rect 7892 4384 8212 5408
rect 7892 4320 7900 4384
rect 7964 4320 7980 4384
rect 8044 4320 8060 4384
rect 8124 4320 8140 4384
rect 8204 4320 8212 4384
rect 7892 3296 8212 4320
rect 7892 3232 7900 3296
rect 7964 3232 7980 3296
rect 8044 3232 8060 3296
rect 8124 3232 8140 3296
rect 8204 3232 8212 3296
rect 7892 2208 8212 3232
rect 7892 2144 7900 2208
rect 7964 2144 7980 2208
rect 8044 2144 8060 2208
rect 8124 2144 8140 2208
rect 8204 2144 8212 2208
rect 7892 2128 8212 2144
rect 11366 27776 11686 27792
rect 11366 27712 11374 27776
rect 11438 27712 11454 27776
rect 11518 27712 11534 27776
rect 11598 27712 11614 27776
rect 11678 27712 11686 27776
rect 11366 26688 11686 27712
rect 11366 26624 11374 26688
rect 11438 26624 11454 26688
rect 11518 26624 11534 26688
rect 11598 26624 11614 26688
rect 11678 26624 11686 26688
rect 11366 25600 11686 26624
rect 11366 25536 11374 25600
rect 11438 25536 11454 25600
rect 11518 25536 11534 25600
rect 11598 25536 11614 25600
rect 11678 25536 11686 25600
rect 11366 24512 11686 25536
rect 11366 24448 11374 24512
rect 11438 24448 11454 24512
rect 11518 24448 11534 24512
rect 11598 24448 11614 24512
rect 11678 24448 11686 24512
rect 11366 23424 11686 24448
rect 11366 23360 11374 23424
rect 11438 23360 11454 23424
rect 11518 23360 11534 23424
rect 11598 23360 11614 23424
rect 11678 23360 11686 23424
rect 11366 22336 11686 23360
rect 11366 22272 11374 22336
rect 11438 22272 11454 22336
rect 11518 22272 11534 22336
rect 11598 22272 11614 22336
rect 11678 22272 11686 22336
rect 11366 21248 11686 22272
rect 11366 21184 11374 21248
rect 11438 21184 11454 21248
rect 11518 21184 11534 21248
rect 11598 21184 11614 21248
rect 11678 21184 11686 21248
rect 11366 20160 11686 21184
rect 11366 20096 11374 20160
rect 11438 20096 11454 20160
rect 11518 20096 11534 20160
rect 11598 20096 11614 20160
rect 11678 20096 11686 20160
rect 11366 19072 11686 20096
rect 11366 19008 11374 19072
rect 11438 19008 11454 19072
rect 11518 19008 11534 19072
rect 11598 19008 11614 19072
rect 11678 19008 11686 19072
rect 11366 17984 11686 19008
rect 11366 17920 11374 17984
rect 11438 17920 11454 17984
rect 11518 17920 11534 17984
rect 11598 17920 11614 17984
rect 11678 17920 11686 17984
rect 11366 16896 11686 17920
rect 11366 16832 11374 16896
rect 11438 16832 11454 16896
rect 11518 16832 11534 16896
rect 11598 16832 11614 16896
rect 11678 16832 11686 16896
rect 11366 15808 11686 16832
rect 11366 15744 11374 15808
rect 11438 15744 11454 15808
rect 11518 15744 11534 15808
rect 11598 15744 11614 15808
rect 11678 15744 11686 15808
rect 11366 14720 11686 15744
rect 11366 14656 11374 14720
rect 11438 14656 11454 14720
rect 11518 14656 11534 14720
rect 11598 14656 11614 14720
rect 11678 14656 11686 14720
rect 11366 13632 11686 14656
rect 11366 13568 11374 13632
rect 11438 13568 11454 13632
rect 11518 13568 11534 13632
rect 11598 13568 11614 13632
rect 11678 13568 11686 13632
rect 11366 12544 11686 13568
rect 11366 12480 11374 12544
rect 11438 12480 11454 12544
rect 11518 12480 11534 12544
rect 11598 12480 11614 12544
rect 11678 12480 11686 12544
rect 11366 11456 11686 12480
rect 11366 11392 11374 11456
rect 11438 11392 11454 11456
rect 11518 11392 11534 11456
rect 11598 11392 11614 11456
rect 11678 11392 11686 11456
rect 11366 10368 11686 11392
rect 11366 10304 11374 10368
rect 11438 10304 11454 10368
rect 11518 10304 11534 10368
rect 11598 10304 11614 10368
rect 11678 10304 11686 10368
rect 11366 9280 11686 10304
rect 11366 9216 11374 9280
rect 11438 9216 11454 9280
rect 11518 9216 11534 9280
rect 11598 9216 11614 9280
rect 11678 9216 11686 9280
rect 11366 8192 11686 9216
rect 11366 8128 11374 8192
rect 11438 8128 11454 8192
rect 11518 8128 11534 8192
rect 11598 8128 11614 8192
rect 11678 8128 11686 8192
rect 11366 7104 11686 8128
rect 11366 7040 11374 7104
rect 11438 7040 11454 7104
rect 11518 7040 11534 7104
rect 11598 7040 11614 7104
rect 11678 7040 11686 7104
rect 11366 6016 11686 7040
rect 11366 5952 11374 6016
rect 11438 5952 11454 6016
rect 11518 5952 11534 6016
rect 11598 5952 11614 6016
rect 11678 5952 11686 6016
rect 11366 4928 11686 5952
rect 11366 4864 11374 4928
rect 11438 4864 11454 4928
rect 11518 4864 11534 4928
rect 11598 4864 11614 4928
rect 11678 4864 11686 4928
rect 11366 3840 11686 4864
rect 11366 3776 11374 3840
rect 11438 3776 11454 3840
rect 11518 3776 11534 3840
rect 11598 3776 11614 3840
rect 11678 3776 11686 3840
rect 11366 2752 11686 3776
rect 11366 2688 11374 2752
rect 11438 2688 11454 2752
rect 11518 2688 11534 2752
rect 11598 2688 11614 2752
rect 11678 2688 11686 2752
rect 11366 2128 11686 2688
rect 14840 27232 15160 27792
rect 14840 27168 14848 27232
rect 14912 27168 14928 27232
rect 14992 27168 15008 27232
rect 15072 27168 15088 27232
rect 15152 27168 15160 27232
rect 14840 26144 15160 27168
rect 14840 26080 14848 26144
rect 14912 26080 14928 26144
rect 14992 26080 15008 26144
rect 15072 26080 15088 26144
rect 15152 26080 15160 26144
rect 14840 25056 15160 26080
rect 14840 24992 14848 25056
rect 14912 24992 14928 25056
rect 14992 24992 15008 25056
rect 15072 24992 15088 25056
rect 15152 24992 15160 25056
rect 14840 23968 15160 24992
rect 14840 23904 14848 23968
rect 14912 23904 14928 23968
rect 14992 23904 15008 23968
rect 15072 23904 15088 23968
rect 15152 23904 15160 23968
rect 14840 22880 15160 23904
rect 14840 22816 14848 22880
rect 14912 22816 14928 22880
rect 14992 22816 15008 22880
rect 15072 22816 15088 22880
rect 15152 22816 15160 22880
rect 14840 21792 15160 22816
rect 14840 21728 14848 21792
rect 14912 21728 14928 21792
rect 14992 21728 15008 21792
rect 15072 21728 15088 21792
rect 15152 21728 15160 21792
rect 14840 20704 15160 21728
rect 14840 20640 14848 20704
rect 14912 20640 14928 20704
rect 14992 20640 15008 20704
rect 15072 20640 15088 20704
rect 15152 20640 15160 20704
rect 14840 19616 15160 20640
rect 14840 19552 14848 19616
rect 14912 19552 14928 19616
rect 14992 19552 15008 19616
rect 15072 19552 15088 19616
rect 15152 19552 15160 19616
rect 14840 18528 15160 19552
rect 14840 18464 14848 18528
rect 14912 18464 14928 18528
rect 14992 18464 15008 18528
rect 15072 18464 15088 18528
rect 15152 18464 15160 18528
rect 14840 17440 15160 18464
rect 14840 17376 14848 17440
rect 14912 17376 14928 17440
rect 14992 17376 15008 17440
rect 15072 17376 15088 17440
rect 15152 17376 15160 17440
rect 14840 16352 15160 17376
rect 14840 16288 14848 16352
rect 14912 16288 14928 16352
rect 14992 16288 15008 16352
rect 15072 16288 15088 16352
rect 15152 16288 15160 16352
rect 14840 15264 15160 16288
rect 14840 15200 14848 15264
rect 14912 15200 14928 15264
rect 14992 15200 15008 15264
rect 15072 15200 15088 15264
rect 15152 15200 15160 15264
rect 14840 14176 15160 15200
rect 14840 14112 14848 14176
rect 14912 14112 14928 14176
rect 14992 14112 15008 14176
rect 15072 14112 15088 14176
rect 15152 14112 15160 14176
rect 14840 13088 15160 14112
rect 14840 13024 14848 13088
rect 14912 13024 14928 13088
rect 14992 13024 15008 13088
rect 15072 13024 15088 13088
rect 15152 13024 15160 13088
rect 14840 12000 15160 13024
rect 14840 11936 14848 12000
rect 14912 11936 14928 12000
rect 14992 11936 15008 12000
rect 15072 11936 15088 12000
rect 15152 11936 15160 12000
rect 14840 10912 15160 11936
rect 14840 10848 14848 10912
rect 14912 10848 14928 10912
rect 14992 10848 15008 10912
rect 15072 10848 15088 10912
rect 15152 10848 15160 10912
rect 14840 9824 15160 10848
rect 14840 9760 14848 9824
rect 14912 9760 14928 9824
rect 14992 9760 15008 9824
rect 15072 9760 15088 9824
rect 15152 9760 15160 9824
rect 14840 8736 15160 9760
rect 14840 8672 14848 8736
rect 14912 8672 14928 8736
rect 14992 8672 15008 8736
rect 15072 8672 15088 8736
rect 15152 8672 15160 8736
rect 14840 7648 15160 8672
rect 14840 7584 14848 7648
rect 14912 7584 14928 7648
rect 14992 7584 15008 7648
rect 15072 7584 15088 7648
rect 15152 7584 15160 7648
rect 14840 6560 15160 7584
rect 14840 6496 14848 6560
rect 14912 6496 14928 6560
rect 14992 6496 15008 6560
rect 15072 6496 15088 6560
rect 15152 6496 15160 6560
rect 14840 5472 15160 6496
rect 14840 5408 14848 5472
rect 14912 5408 14928 5472
rect 14992 5408 15008 5472
rect 15072 5408 15088 5472
rect 15152 5408 15160 5472
rect 14840 4384 15160 5408
rect 14840 4320 14848 4384
rect 14912 4320 14928 4384
rect 14992 4320 15008 4384
rect 15072 4320 15088 4384
rect 15152 4320 15160 4384
rect 14840 3296 15160 4320
rect 14840 3232 14848 3296
rect 14912 3232 14928 3296
rect 14992 3232 15008 3296
rect 15072 3232 15088 3296
rect 15152 3232 15160 3296
rect 14840 2208 15160 3232
rect 14840 2144 14848 2208
rect 14912 2144 14928 2208
rect 14992 2144 15008 2208
rect 15072 2144 15088 2208
rect 15152 2144 15160 2208
rect 14840 2128 15160 2144
rect 18314 27776 18634 27792
rect 18314 27712 18322 27776
rect 18386 27712 18402 27776
rect 18466 27712 18482 27776
rect 18546 27712 18562 27776
rect 18626 27712 18634 27776
rect 18314 26688 18634 27712
rect 18314 26624 18322 26688
rect 18386 26624 18402 26688
rect 18466 26624 18482 26688
rect 18546 26624 18562 26688
rect 18626 26624 18634 26688
rect 18314 25600 18634 26624
rect 18314 25536 18322 25600
rect 18386 25536 18402 25600
rect 18466 25536 18482 25600
rect 18546 25536 18562 25600
rect 18626 25536 18634 25600
rect 18314 24512 18634 25536
rect 18314 24448 18322 24512
rect 18386 24448 18402 24512
rect 18466 24448 18482 24512
rect 18546 24448 18562 24512
rect 18626 24448 18634 24512
rect 18314 23424 18634 24448
rect 18314 23360 18322 23424
rect 18386 23360 18402 23424
rect 18466 23360 18482 23424
rect 18546 23360 18562 23424
rect 18626 23360 18634 23424
rect 18314 22336 18634 23360
rect 18314 22272 18322 22336
rect 18386 22272 18402 22336
rect 18466 22272 18482 22336
rect 18546 22272 18562 22336
rect 18626 22272 18634 22336
rect 18314 21248 18634 22272
rect 18314 21184 18322 21248
rect 18386 21184 18402 21248
rect 18466 21184 18482 21248
rect 18546 21184 18562 21248
rect 18626 21184 18634 21248
rect 18314 20160 18634 21184
rect 18314 20096 18322 20160
rect 18386 20096 18402 20160
rect 18466 20096 18482 20160
rect 18546 20096 18562 20160
rect 18626 20096 18634 20160
rect 18314 19072 18634 20096
rect 18314 19008 18322 19072
rect 18386 19008 18402 19072
rect 18466 19008 18482 19072
rect 18546 19008 18562 19072
rect 18626 19008 18634 19072
rect 18314 17984 18634 19008
rect 18314 17920 18322 17984
rect 18386 17920 18402 17984
rect 18466 17920 18482 17984
rect 18546 17920 18562 17984
rect 18626 17920 18634 17984
rect 18314 16896 18634 17920
rect 18314 16832 18322 16896
rect 18386 16832 18402 16896
rect 18466 16832 18482 16896
rect 18546 16832 18562 16896
rect 18626 16832 18634 16896
rect 18314 15808 18634 16832
rect 18314 15744 18322 15808
rect 18386 15744 18402 15808
rect 18466 15744 18482 15808
rect 18546 15744 18562 15808
rect 18626 15744 18634 15808
rect 18314 14720 18634 15744
rect 18314 14656 18322 14720
rect 18386 14656 18402 14720
rect 18466 14656 18482 14720
rect 18546 14656 18562 14720
rect 18626 14656 18634 14720
rect 18314 13632 18634 14656
rect 18314 13568 18322 13632
rect 18386 13568 18402 13632
rect 18466 13568 18482 13632
rect 18546 13568 18562 13632
rect 18626 13568 18634 13632
rect 18314 12544 18634 13568
rect 18314 12480 18322 12544
rect 18386 12480 18402 12544
rect 18466 12480 18482 12544
rect 18546 12480 18562 12544
rect 18626 12480 18634 12544
rect 18314 11456 18634 12480
rect 18314 11392 18322 11456
rect 18386 11392 18402 11456
rect 18466 11392 18482 11456
rect 18546 11392 18562 11456
rect 18626 11392 18634 11456
rect 18314 10368 18634 11392
rect 18314 10304 18322 10368
rect 18386 10304 18402 10368
rect 18466 10304 18482 10368
rect 18546 10304 18562 10368
rect 18626 10304 18634 10368
rect 18314 9280 18634 10304
rect 18314 9216 18322 9280
rect 18386 9216 18402 9280
rect 18466 9216 18482 9280
rect 18546 9216 18562 9280
rect 18626 9216 18634 9280
rect 18314 8192 18634 9216
rect 18314 8128 18322 8192
rect 18386 8128 18402 8192
rect 18466 8128 18482 8192
rect 18546 8128 18562 8192
rect 18626 8128 18634 8192
rect 18314 7104 18634 8128
rect 18314 7040 18322 7104
rect 18386 7040 18402 7104
rect 18466 7040 18482 7104
rect 18546 7040 18562 7104
rect 18626 7040 18634 7104
rect 18314 6016 18634 7040
rect 18314 5952 18322 6016
rect 18386 5952 18402 6016
rect 18466 5952 18482 6016
rect 18546 5952 18562 6016
rect 18626 5952 18634 6016
rect 18314 4928 18634 5952
rect 18314 4864 18322 4928
rect 18386 4864 18402 4928
rect 18466 4864 18482 4928
rect 18546 4864 18562 4928
rect 18626 4864 18634 4928
rect 18314 3840 18634 4864
rect 18314 3776 18322 3840
rect 18386 3776 18402 3840
rect 18466 3776 18482 3840
rect 18546 3776 18562 3840
rect 18626 3776 18634 3840
rect 18314 2752 18634 3776
rect 18314 2688 18322 2752
rect 18386 2688 18402 2752
rect 18466 2688 18482 2752
rect 18546 2688 18562 2752
rect 18626 2688 18634 2752
rect 18314 2128 18634 2688
rect 21788 27232 22108 27792
rect 21788 27168 21796 27232
rect 21860 27168 21876 27232
rect 21940 27168 21956 27232
rect 22020 27168 22036 27232
rect 22100 27168 22108 27232
rect 21788 26144 22108 27168
rect 21788 26080 21796 26144
rect 21860 26080 21876 26144
rect 21940 26080 21956 26144
rect 22020 26080 22036 26144
rect 22100 26080 22108 26144
rect 21788 25056 22108 26080
rect 21788 24992 21796 25056
rect 21860 24992 21876 25056
rect 21940 24992 21956 25056
rect 22020 24992 22036 25056
rect 22100 24992 22108 25056
rect 21788 23968 22108 24992
rect 21788 23904 21796 23968
rect 21860 23904 21876 23968
rect 21940 23904 21956 23968
rect 22020 23904 22036 23968
rect 22100 23904 22108 23968
rect 21788 22880 22108 23904
rect 21788 22816 21796 22880
rect 21860 22816 21876 22880
rect 21940 22816 21956 22880
rect 22020 22816 22036 22880
rect 22100 22816 22108 22880
rect 21788 21792 22108 22816
rect 21788 21728 21796 21792
rect 21860 21728 21876 21792
rect 21940 21728 21956 21792
rect 22020 21728 22036 21792
rect 22100 21728 22108 21792
rect 21788 20704 22108 21728
rect 21788 20640 21796 20704
rect 21860 20640 21876 20704
rect 21940 20640 21956 20704
rect 22020 20640 22036 20704
rect 22100 20640 22108 20704
rect 21788 19616 22108 20640
rect 21788 19552 21796 19616
rect 21860 19552 21876 19616
rect 21940 19552 21956 19616
rect 22020 19552 22036 19616
rect 22100 19552 22108 19616
rect 21788 18528 22108 19552
rect 21788 18464 21796 18528
rect 21860 18464 21876 18528
rect 21940 18464 21956 18528
rect 22020 18464 22036 18528
rect 22100 18464 22108 18528
rect 21788 17440 22108 18464
rect 21788 17376 21796 17440
rect 21860 17376 21876 17440
rect 21940 17376 21956 17440
rect 22020 17376 22036 17440
rect 22100 17376 22108 17440
rect 21788 16352 22108 17376
rect 21788 16288 21796 16352
rect 21860 16288 21876 16352
rect 21940 16288 21956 16352
rect 22020 16288 22036 16352
rect 22100 16288 22108 16352
rect 21788 15264 22108 16288
rect 21788 15200 21796 15264
rect 21860 15200 21876 15264
rect 21940 15200 21956 15264
rect 22020 15200 22036 15264
rect 22100 15200 22108 15264
rect 21788 14176 22108 15200
rect 21788 14112 21796 14176
rect 21860 14112 21876 14176
rect 21940 14112 21956 14176
rect 22020 14112 22036 14176
rect 22100 14112 22108 14176
rect 21788 13088 22108 14112
rect 21788 13024 21796 13088
rect 21860 13024 21876 13088
rect 21940 13024 21956 13088
rect 22020 13024 22036 13088
rect 22100 13024 22108 13088
rect 21788 12000 22108 13024
rect 21788 11936 21796 12000
rect 21860 11936 21876 12000
rect 21940 11936 21956 12000
rect 22020 11936 22036 12000
rect 22100 11936 22108 12000
rect 21788 10912 22108 11936
rect 21788 10848 21796 10912
rect 21860 10848 21876 10912
rect 21940 10848 21956 10912
rect 22020 10848 22036 10912
rect 22100 10848 22108 10912
rect 21788 9824 22108 10848
rect 21788 9760 21796 9824
rect 21860 9760 21876 9824
rect 21940 9760 21956 9824
rect 22020 9760 22036 9824
rect 22100 9760 22108 9824
rect 21788 8736 22108 9760
rect 21788 8672 21796 8736
rect 21860 8672 21876 8736
rect 21940 8672 21956 8736
rect 22020 8672 22036 8736
rect 22100 8672 22108 8736
rect 21788 7648 22108 8672
rect 21788 7584 21796 7648
rect 21860 7584 21876 7648
rect 21940 7584 21956 7648
rect 22020 7584 22036 7648
rect 22100 7584 22108 7648
rect 21788 6560 22108 7584
rect 21788 6496 21796 6560
rect 21860 6496 21876 6560
rect 21940 6496 21956 6560
rect 22020 6496 22036 6560
rect 22100 6496 22108 6560
rect 21788 5472 22108 6496
rect 21788 5408 21796 5472
rect 21860 5408 21876 5472
rect 21940 5408 21956 5472
rect 22020 5408 22036 5472
rect 22100 5408 22108 5472
rect 21788 4384 22108 5408
rect 21788 4320 21796 4384
rect 21860 4320 21876 4384
rect 21940 4320 21956 4384
rect 22020 4320 22036 4384
rect 22100 4320 22108 4384
rect 21788 3296 22108 4320
rect 21788 3232 21796 3296
rect 21860 3232 21876 3296
rect 21940 3232 21956 3296
rect 22020 3232 22036 3296
rect 22100 3232 22108 3296
rect 21788 2208 22108 3232
rect 21788 2144 21796 2208
rect 21860 2144 21876 2208
rect 21940 2144 21956 2208
rect 22020 2144 22036 2208
rect 22100 2144 22108 2208
rect 21788 2128 22108 2144
rect 25262 27776 25582 27792
rect 25262 27712 25270 27776
rect 25334 27712 25350 27776
rect 25414 27712 25430 27776
rect 25494 27712 25510 27776
rect 25574 27712 25582 27776
rect 25262 26688 25582 27712
rect 25262 26624 25270 26688
rect 25334 26624 25350 26688
rect 25414 26624 25430 26688
rect 25494 26624 25510 26688
rect 25574 26624 25582 26688
rect 25262 25600 25582 26624
rect 25262 25536 25270 25600
rect 25334 25536 25350 25600
rect 25414 25536 25430 25600
rect 25494 25536 25510 25600
rect 25574 25536 25582 25600
rect 25262 24512 25582 25536
rect 25262 24448 25270 24512
rect 25334 24448 25350 24512
rect 25414 24448 25430 24512
rect 25494 24448 25510 24512
rect 25574 24448 25582 24512
rect 25262 23424 25582 24448
rect 25262 23360 25270 23424
rect 25334 23360 25350 23424
rect 25414 23360 25430 23424
rect 25494 23360 25510 23424
rect 25574 23360 25582 23424
rect 25262 22336 25582 23360
rect 25262 22272 25270 22336
rect 25334 22272 25350 22336
rect 25414 22272 25430 22336
rect 25494 22272 25510 22336
rect 25574 22272 25582 22336
rect 25262 21248 25582 22272
rect 25262 21184 25270 21248
rect 25334 21184 25350 21248
rect 25414 21184 25430 21248
rect 25494 21184 25510 21248
rect 25574 21184 25582 21248
rect 25262 20160 25582 21184
rect 25262 20096 25270 20160
rect 25334 20096 25350 20160
rect 25414 20096 25430 20160
rect 25494 20096 25510 20160
rect 25574 20096 25582 20160
rect 25262 19072 25582 20096
rect 25262 19008 25270 19072
rect 25334 19008 25350 19072
rect 25414 19008 25430 19072
rect 25494 19008 25510 19072
rect 25574 19008 25582 19072
rect 25262 17984 25582 19008
rect 25262 17920 25270 17984
rect 25334 17920 25350 17984
rect 25414 17920 25430 17984
rect 25494 17920 25510 17984
rect 25574 17920 25582 17984
rect 25262 16896 25582 17920
rect 25262 16832 25270 16896
rect 25334 16832 25350 16896
rect 25414 16832 25430 16896
rect 25494 16832 25510 16896
rect 25574 16832 25582 16896
rect 25262 15808 25582 16832
rect 25262 15744 25270 15808
rect 25334 15744 25350 15808
rect 25414 15744 25430 15808
rect 25494 15744 25510 15808
rect 25574 15744 25582 15808
rect 25262 14720 25582 15744
rect 25262 14656 25270 14720
rect 25334 14656 25350 14720
rect 25414 14656 25430 14720
rect 25494 14656 25510 14720
rect 25574 14656 25582 14720
rect 25262 13632 25582 14656
rect 25262 13568 25270 13632
rect 25334 13568 25350 13632
rect 25414 13568 25430 13632
rect 25494 13568 25510 13632
rect 25574 13568 25582 13632
rect 25262 12544 25582 13568
rect 25262 12480 25270 12544
rect 25334 12480 25350 12544
rect 25414 12480 25430 12544
rect 25494 12480 25510 12544
rect 25574 12480 25582 12544
rect 25262 11456 25582 12480
rect 25262 11392 25270 11456
rect 25334 11392 25350 11456
rect 25414 11392 25430 11456
rect 25494 11392 25510 11456
rect 25574 11392 25582 11456
rect 25262 10368 25582 11392
rect 25262 10304 25270 10368
rect 25334 10304 25350 10368
rect 25414 10304 25430 10368
rect 25494 10304 25510 10368
rect 25574 10304 25582 10368
rect 25262 9280 25582 10304
rect 25262 9216 25270 9280
rect 25334 9216 25350 9280
rect 25414 9216 25430 9280
rect 25494 9216 25510 9280
rect 25574 9216 25582 9280
rect 25262 8192 25582 9216
rect 25262 8128 25270 8192
rect 25334 8128 25350 8192
rect 25414 8128 25430 8192
rect 25494 8128 25510 8192
rect 25574 8128 25582 8192
rect 25262 7104 25582 8128
rect 25262 7040 25270 7104
rect 25334 7040 25350 7104
rect 25414 7040 25430 7104
rect 25494 7040 25510 7104
rect 25574 7040 25582 7104
rect 25262 6016 25582 7040
rect 25262 5952 25270 6016
rect 25334 5952 25350 6016
rect 25414 5952 25430 6016
rect 25494 5952 25510 6016
rect 25574 5952 25582 6016
rect 25262 4928 25582 5952
rect 25262 4864 25270 4928
rect 25334 4864 25350 4928
rect 25414 4864 25430 4928
rect 25494 4864 25510 4928
rect 25574 4864 25582 4928
rect 25262 3840 25582 4864
rect 25262 3776 25270 3840
rect 25334 3776 25350 3840
rect 25414 3776 25430 3840
rect 25494 3776 25510 3840
rect 25574 3776 25582 3840
rect 25262 2752 25582 3776
rect 25262 2688 25270 2752
rect 25334 2688 25350 2752
rect 25414 2688 25430 2752
rect 25494 2688 25510 2752
rect 25574 2688 25582 2752
rect 25262 2128 25582 2688
use sky130_ef_sc_hd__decap_12  FILLER_0_3 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70
timestamp 1649977179
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1649977179
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1649977179
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1649977179
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1649977179
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1649977179
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_153
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1649977179
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1649977179
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1649977179
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_295
timestamp 1649977179
transform 1 0 28244 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1649977179
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1649977179
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1649977179
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_289
timestamp 1649977179
transform 1 0 27692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_295
timestamp 1649977179
transform 1 0 28244 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1649977179
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1649977179
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1649977179
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1649977179
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1649977179
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1649977179
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1649977179
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1649977179
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1649977179
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1649977179
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1649977179
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1649977179
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_57
timestamp 1649977179
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_69
timestamp 1649977179
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1649977179
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_113
timestamp 1649977179
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_125
timestamp 1649977179
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1649977179
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_169
timestamp 1649977179
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_181
timestamp 1649977179
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1649977179
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_225
timestamp 1649977179
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1649977179
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1649977179
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_281
timestamp 1649977179
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_293
timestamp 1649977179
transform 1 0 28060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0_ ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  okk_3 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output2 ~/rioschip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7544 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 hehe_rstn
port 0 nsew signal tristate
flabel metal3 s 29200 16328 30000 16448 0 FreeSans 480 0 0 0 la_data_in[0]
port 1 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 2 nsew signal input
flabel metal3 s 29200 21768 30000 21888 0 FreeSans 480 0 0 0 la_data_in[101]
port 3 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 4 nsew signal input
flabel metal2 s 29642 29200 29698 30000 0 FreeSans 224 90 0 0 la_data_in[103]
port 5 nsew signal input
flabel metal3 s 29200 6808 30000 6928 0 FreeSans 480 0 0 0 la_data_in[104]
port 6 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 la_data_in[105]
port 7 nsew signal input
flabel metal2 s 12898 29200 12954 30000 0 FreeSans 224 90 0 0 la_data_in[106]
port 8 nsew signal input
flabel metal2 s 15474 29200 15530 30000 0 FreeSans 224 90 0 0 la_data_in[107]
port 9 nsew signal input
flabel metal2 s 26422 29200 26478 30000 0 FreeSans 224 90 0 0 la_data_in[108]
port 10 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 11 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 la_data_in[10]
port 12 nsew signal input
flabel metal2 s 28998 29200 29054 30000 0 FreeSans 224 90 0 0 la_data_in[110]
port 13 nsew signal input
flabel metal2 s 2594 29200 2650 30000 0 FreeSans 224 90 0 0 la_data_in[111]
port 14 nsew signal input
flabel metal2 s 24490 29200 24546 30000 0 FreeSans 224 90 0 0 la_data_in[112]
port 15 nsew signal input
flabel metal2 s 12254 29200 12310 30000 0 FreeSans 224 90 0 0 la_data_in[113]
port 16 nsew signal input
flabel metal3 s 29200 10208 30000 10328 0 FreeSans 480 0 0 0 la_data_in[114]
port 17 nsew signal input
flabel metal3 s 29200 14288 30000 14408 0 FreeSans 480 0 0 0 la_data_in[115]
port 18 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 19 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 la_data_in[117]
port 20 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 21 nsew signal input
flabel metal2 s 7746 29200 7802 30000 0 FreeSans 224 90 0 0 la_data_in[119]
port 22 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 23 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 24 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 25 nsew signal input
flabel metal3 s 29200 17008 30000 17128 0 FreeSans 480 0 0 0 la_data_in[122]
port 26 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 27 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 28 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 la_data_in[125]
port 29 nsew signal input
flabel metal3 s 29200 21088 30000 21208 0 FreeSans 480 0 0 0 la_data_in[126]
port 30 nsew signal input
flabel metal2 s 8390 29200 8446 30000 0 FreeSans 224 90 0 0 la_data_in[127]
port 31 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 32 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 la_data_in[13]
port 33 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 la_data_in[14]
port 34 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 la_data_in[15]
port 35 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 la_data_in[16]
port 36 nsew signal input
flabel metal2 s 28354 29200 28410 30000 0 FreeSans 224 90 0 0 la_data_in[17]
port 37 nsew signal input
flabel metal2 s 25134 29200 25190 30000 0 FreeSans 224 90 0 0 la_data_in[18]
port 38 nsew signal input
flabel metal2 s 6458 29200 6514 30000 0 FreeSans 224 90 0 0 la_data_in[19]
port 39 nsew signal input
flabel metal3 s 29200 9528 30000 9648 0 FreeSans 480 0 0 0 la_data_in[1]
port 40 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 41 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 la_data_in[21]
port 42 nsew signal input
flabel metal2 s 4526 29200 4582 30000 0 FreeSans 224 90 0 0 la_data_in[22]
port 43 nsew signal input
flabel metal2 s 16118 29200 16174 30000 0 FreeSans 224 90 0 0 la_data_in[23]
port 44 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 45 nsew signal input
flabel metal2 s 20626 29200 20682 30000 0 FreeSans 224 90 0 0 la_data_in[25]
port 46 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 la_data_in[26]
port 47 nsew signal input
flabel metal2 s 19982 29200 20038 30000 0 FreeSans 224 90 0 0 la_data_in[27]
port 48 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 la_data_in[28]
port 49 nsew signal input
flabel metal3 s 29200 27888 30000 28008 0 FreeSans 480 0 0 0 la_data_in[29]
port 50 nsew signal input
flabel metal3 s 29200 23128 30000 23248 0 FreeSans 480 0 0 0 la_data_in[2]
port 51 nsew signal input
flabel metal3 s 29200 19048 30000 19168 0 FreeSans 480 0 0 0 la_data_in[30]
port 52 nsew signal input
flabel metal3 s 29200 2048 30000 2168 0 FreeSans 480 0 0 0 la_data_in[31]
port 53 nsew signal input
flabel metal2 s 10322 29200 10378 30000 0 FreeSans 224 90 0 0 la_data_in[32]
port 54 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 55 nsew signal input
flabel metal3 s 29200 28568 30000 28688 0 FreeSans 480 0 0 0 la_data_in[34]
port 56 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 57 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 la_data_in[36]
port 58 nsew signal input
flabel metal2 s 18050 29200 18106 30000 0 FreeSans 224 90 0 0 la_data_in[37]
port 59 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 la_data_in[38]
port 60 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 la_data_in[39]
port 61 nsew signal input
flabel metal2 s 1950 29200 2006 30000 0 FreeSans 224 90 0 0 la_data_in[3]
port 62 nsew signal input
flabel metal3 s 29200 25168 30000 25288 0 FreeSans 480 0 0 0 la_data_in[40]
port 63 nsew signal input
flabel metal2 s 3882 29200 3938 30000 0 FreeSans 224 90 0 0 la_data_in[41]
port 64 nsew signal input
flabel metal2 s 10966 29200 11022 30000 0 FreeSans 224 90 0 0 la_data_in[42]
port 65 nsew signal input
flabel metal2 s 13542 29200 13598 30000 0 FreeSans 224 90 0 0 la_data_in[43]
port 66 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 la_data_in[44]
port 67 nsew signal input
flabel metal3 s 29200 11568 30000 11688 0 FreeSans 480 0 0 0 la_data_in[45]
port 68 nsew signal input
flabel metal3 s 29200 7488 30000 7608 0 FreeSans 480 0 0 0 la_data_in[46]
port 69 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 la_data_in[47]
port 70 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 71 nsew signal input
flabel metal3 s 29200 8 30000 128 0 FreeSans 480 0 0 0 la_data_in[49]
port 72 nsew signal input
flabel metal3 s 29200 8848 30000 8968 0 FreeSans 480 0 0 0 la_data_in[4]
port 73 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 la_data_in[50]
port 74 nsew signal input
flabel metal3 s 29200 4768 30000 4888 0 FreeSans 480 0 0 0 la_data_in[51]
port 75 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 la_data_in[52]
port 76 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 77 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 la_data_in[54]
port 78 nsew signal input
flabel metal3 s 29200 26528 30000 26648 0 FreeSans 480 0 0 0 la_data_in[55]
port 79 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 80 nsew signal input
flabel metal3 s 29200 2728 30000 2848 0 FreeSans 480 0 0 0 la_data_in[57]
port 81 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 la_data_in[58]
port 82 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 83 nsew signal input
flabel metal2 s 14830 29200 14886 30000 0 FreeSans 224 90 0 0 la_data_in[5]
port 84 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 85 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 86 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 87 nsew signal input
flabel metal3 s 29200 1368 30000 1488 0 FreeSans 480 0 0 0 la_data_in[63]
port 88 nsew signal input
flabel metal3 s 29200 20408 30000 20528 0 FreeSans 480 0 0 0 la_data_in[64]
port 89 nsew signal input
flabel metal3 s 29200 12248 30000 12368 0 FreeSans 480 0 0 0 la_data_in[65]
port 90 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 91 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 la_data_in[67]
port 92 nsew signal input
flabel metal3 s 29200 6128 30000 6248 0 FreeSans 480 0 0 0 la_data_in[68]
port 93 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 la_data_in[69]
port 94 nsew signal input
flabel metal3 s 29200 15648 30000 15768 0 FreeSans 480 0 0 0 la_data_in[6]
port 95 nsew signal input
flabel metal3 s 29200 23808 30000 23928 0 FreeSans 480 0 0 0 la_data_in[70]
port 96 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 97 nsew signal input
flabel metal3 s 29200 25848 30000 25968 0 FreeSans 480 0 0 0 la_data_in[72]
port 98 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 la_data_in[73]
port 99 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 la_data_in[74]
port 100 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 la_data_in[75]
port 101 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 102 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 103 nsew signal input
flabel metal2 s 18 29200 74 30000 0 FreeSans 224 90 0 0 la_data_in[78]
port 104 nsew signal input
flabel metal2 s 9034 29200 9090 30000 0 FreeSans 224 90 0 0 la_data_in[79]
port 105 nsew signal input
flabel metal2 s 19338 29200 19394 30000 0 FreeSans 224 90 0 0 la_data_in[7]
port 106 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 la_data_in[80]
port 107 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 la_data_in[81]
port 108 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 109 nsew signal input
flabel metal2 s 23846 29200 23902 30000 0 FreeSans 224 90 0 0 la_data_in[83]
port 110 nsew signal input
flabel metal2 s 17406 29200 17462 30000 0 FreeSans 224 90 0 0 la_data_in[84]
port 111 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 112 nsew signal input
flabel metal2 s 27066 29200 27122 30000 0 FreeSans 224 90 0 0 la_data_in[86]
port 113 nsew signal input
flabel metal3 s 29200 4088 30000 4208 0 FreeSans 480 0 0 0 la_data_in[87]
port 114 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 la_data_in[88]
port 115 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 la_data_in[89]
port 116 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 117 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 118 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 119 nsew signal input
flabel metal3 s 29200 18368 30000 18488 0 FreeSans 480 0 0 0 la_data_in[92]
port 120 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 121 nsew signal input
flabel metal2 s 22558 29200 22614 30000 0 FreeSans 224 90 0 0 la_data_in[94]
port 122 nsew signal input
flabel metal2 s 21914 29200 21970 30000 0 FreeSans 224 90 0 0 la_data_in[95]
port 123 nsew signal input
flabel metal2 s 1306 29200 1362 30000 0 FreeSans 224 90 0 0 la_data_in[96]
port 124 nsew signal input
flabel metal2 s 5814 29200 5870 30000 0 FreeSans 224 90 0 0 la_data_in[97]
port 125 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 126 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 la_data_in[99]
port 127 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 la_data_in[9]
port 128 nsew signal input
flabel metal3 s 29200 13608 30000 13728 0 FreeSans 480 0 0 0 meip
port 129 nsew signal tristate
flabel metal4 s 4418 2128 4738 27792 0 FreeSans 1920 90 0 0 vccd1
port 130 nsew power bidirectional
flabel metal4 s 11366 2128 11686 27792 0 FreeSans 1920 90 0 0 vccd1
port 130 nsew power bidirectional
flabel metal4 s 18314 2128 18634 27792 0 FreeSans 1920 90 0 0 vccd1
port 130 nsew power bidirectional
flabel metal4 s 25262 2128 25582 27792 0 FreeSans 1920 90 0 0 vccd1
port 130 nsew power bidirectional
flabel metal4 s 7892 2128 8212 27792 0 FreeSans 1920 90 0 0 vssd1
port 131 nsew ground bidirectional
flabel metal4 s 14840 2128 15160 27792 0 FreeSans 1920 90 0 0 vssd1
port 131 nsew ground bidirectional
flabel metal4 s 21788 2128 22108 27792 0 FreeSans 1920 90 0 0 vssd1
port 131 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
